* File: sky130_osu_sc_18T_ms__mux2_1.pex.spice
* Created: Fri Nov 12 14:05:03 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%GND 1 29 33 54 56
r35 54 56 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r36 31 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r37 29 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r38 29 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r39 29 31 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r40 29 35 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r41 29 35 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r42 1 33 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%VDD 1 9 13 19 23
r30 23 26 0.00227273 $w=2.75e-06 $l=5e-08 $layer=MET1_cond $X=1.375 $Y=6.42
+ $X2=1.375 $Y2=6.47
r31 19 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.38 $Y=6.47
+ $X2=2.38 $Y2=6.47
r32 17 19 76.8925 $w=3.03e-07 $l=2.035e-06 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=2.38 $Y2=6.507
r33 13 16 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r34 11 17 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.345 $Y2=6.507
r35 11 16 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r36 9 19 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r37 1 16 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r38 1 13 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%A_110_115# 1 3 9 11 15 19 24 28 31 34 37
+ 44 49
c69 9 0 3.63536e-20 $X=1.35 $Y=1.79
r70 46 49 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=2.69
+ $X2=0.925 $Y2=2.69
r71 41 44 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.925 $Y2=1.85
r72 37 39 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r73 35 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.855
+ $X2=0.69 $Y2=2.69
r74 35 37 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.69 $Y=2.855 $X2=0.69
+ $Y2=3.455
r75 34 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.525
+ $X2=0.69 $Y2=2.69
r76 33 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.015
+ $X2=0.69 $Y2=1.85
r77 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.69 $Y=2.015
+ $X2=0.69 $Y2=2.525
r78 29 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.685
+ $X2=0.69 $Y2=1.85
r79 29 31 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.69 $Y=1.685
+ $X2=0.69 $Y2=0.825
r80 26 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.69 $X2=0.925 $Y2=2.69
r81 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.69
+ $X2=1.09 $Y2=2.69
r82 22 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.85 $X2=0.925 $Y2=1.85
r83 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.85
+ $X2=1.09 $Y2=1.85
r84 17 19 964 $w=1.5e-07 $l=1.88e-06 $layer=POLY_cond $X=1.855 $Y=2.705
+ $X2=1.855 $Y2=4.585
r85 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.425 $Y=1.715
+ $X2=1.425 $Y2=1.075
r86 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.63
+ $X2=1.855 $Y2=2.705
r87 11 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.78 $Y=2.63
+ $X2=1.09 $Y2=2.63
r88 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=1.79
+ $X2=1.425 $Y2=1.715
r89 9 24 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.35 $Y=1.79 $X2=1.09
+ $Y2=1.79
r90 3 39 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r91 3 37 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r92 1 31 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%S0 3 8 9 11 12 13 15 18 24 26 32
c65 8 0 1.8854e-20 $X=0.475 $Y=4.585
r66 29 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r67 26 29 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.27 $Y=2.305
+ $X2=0.27 $Y2=3.33
r68 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.305
+ $X2=0.55 $Y2=2.305
r69 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.305 $X2=0.27 $Y2=2.305
r70 21 23 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.305
+ $X2=0.475 $Y2=2.305
r71 16 18 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.855 $Y=2.195
+ $X2=1.855 $Y2=1.075
r72 13 15 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.425 $Y=6.16
+ $X2=1.425 $Y2=4.585
r73 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=6.235
+ $X2=1.425 $Y2=6.16
r74 11 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.35 $Y=6.235 $X2=0.55
+ $Y2=6.235
r75 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.27
+ $X2=1.855 $Y2=2.195
r76 9 24 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.78 $Y=2.27
+ $X2=0.55 $Y2=2.27
r77 6 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=6.16
+ $X2=0.55 $Y2=6.235
r78 6 8 807.606 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=6.16
+ $X2=0.475 $Y2=4.585
r79 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=2.305
r80 5 8 1084.5 $w=1.5e-07 $l=2.115e-06 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=4.585
r81 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.14
+ $X2=0.475 $Y2=2.305
r82 1 3 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=0.475 $Y=2.14
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%A0 1 3 11 15 22 24 26 28
c41 28 0 1.8854e-20 $X=1.265 $Y=2.96
r42 25 26 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=3.115
+ $X2=1.237 $Y2=3.285
r43 23 24 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=1.335
+ $X2=1.237 $Y2=1.505
r44 22 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.265 $Y=2.96
+ $X2=1.265 $Y2=2.96
r45 22 25 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.265 $Y=2.96
+ $X2=1.265 $Y2=3.115
r46 22 24 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=1.265 $Y=2.96
+ $X2=1.265 $Y2=1.505
r47 15 17 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.21 $Y=3.455
+ $X2=1.21 $Y2=5.835
r48 15 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.21 $Y=3.455
+ $X2=1.21 $Y2=3.285
r49 11 23 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.21 $Y=0.825
+ $X2=1.21 $Y2=1.335
r50 3 17 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=1.085
+ $Y=3.085 $X2=1.21 $Y2=5.835
r51 3 15 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=1.085
+ $Y=3.085 $X2=1.21 $Y2=3.455
r52 1 11 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%Y 1 3 10 16 24 26 29
c37 29 0 3.63536e-20 $X=1.64 $Y=2.22
r38 24 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=2.105
+ $X2=1.64 $Y2=2.22
r39 23 26 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=1.595
+ $X2=1.64 $Y2=1.48
r40 23 24 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=1.64 $Y=1.595
+ $X2=1.64 $Y2=2.105
r41 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.64 $Y=3.455
+ $X2=1.64 $Y2=5.835
r42 16 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=2.22
+ $X2=1.64 $Y2=2.22
r43 16 19 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.64 $Y=2.22
+ $X2=1.64 $Y2=3.455
r44 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.48
+ $X2=1.64 $Y2=1.48
r45 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.64 $Y=0.825
+ $X2=1.64 $Y2=1.48
r46 3 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=5.835
r47 3 19 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=3.455
r48 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__MUX2_1%A1 1 3 10 20
r17 15 17 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.07 $Y=3.455
+ $X2=2.07 $Y2=5.835
r18 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.59
+ $X2=2.07 $Y2=2.59
r19 13 15 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.07 $Y=2.59
+ $X2=2.07 $Y2=3.455
r20 10 13 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.07 $Y=0.825
+ $X2=2.07 $Y2=2.59
r21 3 17 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=5.835
r22 3 15 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=3.455
r23 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

