* File: sky130_osu_sc_15T_ms__dffs_1.pex.spice
* Created: Fri Nov 12 14:42:48 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%GND 1 2 3 4 5 6 97 99 107 113 115 125
+ 127 137 139 149 151 158 180 182
c197 137 0 1.67294e-19 $X=5.14 $Y=0.865
c198 113 0 3.07193e-19 $X=1.64 $Y=0.865
c199 97 0 1.27355e-19 $X=-0.05 $Y=0
r200 180 182 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=7.815 $Y2=0.152
r201 156 158 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.74
r202 152 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=0.152
+ $X2=6.88 $Y2=0.152
r203 147 172 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.152
r204 147 149 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.74
r205 139 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=0.152
+ $X2=6.88 $Y2=0.152
r206 135 137 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.14 $Y=0.305
+ $X2=5.14 $Y2=0.865
r207 128 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.152
+ $X2=3.39 $Y2=0.152
r208 123 168 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.152
r209 123 125 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.74
r210 115 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.152
+ $X2=3.39 $Y2=0.152
r211 111 113 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.64 $Y=0.305
+ $X2=1.64 $Y2=0.865
r212 109 110 15.8697 $w=3.03e-07 $l=4.2e-07 $layer=LI1_cond $X=1.555 $Y=0.152
+ $X2=1.135 $Y2=0.152
r213 105 107 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r214 97 182 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=0.19
+ $X2=7.815 $Y2=0.19
r215 97 180 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r216 97 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r217 97 151 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r218 97 135 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.14 $Y2=0.305
r219 97 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.055 $Y2=0.152
r220 97 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.225 $Y2=0.152
r221 97 111 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.64 $Y2=0.305
r222 97 109 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.555 $Y2=0.152
r223 97 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.725 $Y2=0.152
r224 97 105 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r225 97 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r226 97 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r227 97 151 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r228 97 152 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.965 $Y2=0.152
r229 97 139 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.795 $Y2=0.152
r230 97 140 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=5.225 $Y2=0.152
r231 97 127 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=5.055 $Y2=0.152
r232 97 128 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.475 $Y2=0.152
r233 97 115 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=3.305 $Y2=0.152
r234 97 116 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=1.725 $Y2=0.152
r235 97 99 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=0.335 $Y=0.152
+ $X2=0.965 $Y2=0.152
r236 6 158 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.74
r237 5 149 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.575 $X2=6.88 $Y2=0.74
r238 4 137 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=5
+ $Y=0.575 $X2=5.14 $Y2=0.865
r239 3 125 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.575 $X2=3.39 $Y2=0.74
r240 2 113 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.575 $X2=1.64 $Y2=0.865
r241 1 107 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%VDD 1 2 3 4 5 6 7 8 81 85 87 93 99 103
+ 111 115 123 127 133 135 141 143 149 165 168 172
r104 168 172 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=5.397
+ $X2=7.815 $Y2=5.397
r105 165 172 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=5.36
+ $X2=7.815 $Y2=5.36
r106 154 168 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=5.36
+ $X2=0.335 $Y2=5.36
r107 147 165 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=5.245
+ $X2=7.9 $Y2=5.397
r108 147 149 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.9 $Y=5.245
+ $X2=7.9 $Y2=4.225
r109 144 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.035 $Y=5.397
+ $X2=6.95 $Y2=5.397
r110 144 146 3.7785 $w=3.03e-07 $l=1e-07 $layer=LI1_cond $X=7.035 $Y=5.397
+ $X2=7.135 $Y2=5.397
r111 143 165 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=5.397
+ $X2=7.9 $Y2=5.397
r112 143 146 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=5.397
+ $X2=7.135 $Y2=5.397
r113 139 163 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.95 $Y=5.245
+ $X2=6.95 $Y2=5.397
r114 139 141 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.95 $Y=5.245
+ $X2=6.95 $Y2=4.565
r115 136 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=5.397
+ $X2=6.09 $Y2=5.397
r116 136 138 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=5.397
+ $X2=6.455 $Y2=5.397
r117 135 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=5.397
+ $X2=6.95 $Y2=5.397
r118 135 138 15.4919 $w=3.03e-07 $l=4.1e-07 $layer=LI1_cond $X=6.865 $Y=5.397
+ $X2=6.455 $Y2=5.397
r119 131 162 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=5.245
+ $X2=6.09 $Y2=5.397
r120 131 133 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.09 $Y=5.245
+ $X2=6.09 $Y2=4.565
r121 128 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=5.397
+ $X2=5.14 $Y2=5.397
r122 128 130 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.225 $Y=5.397
+ $X2=5.775 $Y2=5.397
r123 127 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=5.397
+ $X2=6.09 $Y2=5.397
r124 127 130 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=5.397
+ $X2=5.775 $Y2=5.397
r125 123 126 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=5.14 $Y=3.205
+ $X2=5.14 $Y2=4.565
r126 121 161 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.14 $Y=5.245
+ $X2=5.14 $Y2=5.397
r127 121 126 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.14 $Y=5.245
+ $X2=5.14 $Y2=4.565
r128 118 120 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=5.397
+ $X2=4.415 $Y2=5.397
r129 116 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=5.397
+ $X2=3.39 $Y2=5.397
r130 116 118 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.475 $Y=5.397
+ $X2=3.735 $Y2=5.397
r131 115 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=5.397
+ $X2=5.14 $Y2=5.397
r132 115 120 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=5.055 $Y=5.397
+ $X2=4.415 $Y2=5.397
r133 111 114 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.39 $Y=3.545
+ $X2=3.39 $Y2=4.565
r134 109 159 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.39 $Y=5.245
+ $X2=3.39 $Y2=5.397
r135 109 114 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.39 $Y=5.245
+ $X2=3.39 $Y2=4.565
r136 106 108 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.375 $Y=5.397
+ $X2=3.055 $Y2=5.397
r137 104 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=5.397
+ $X2=1.64 $Y2=5.397
r138 104 106 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=1.725 $Y=5.397
+ $X2=2.375 $Y2=5.397
r139 103 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=5.397
+ $X2=3.39 $Y2=5.397
r140 103 108 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.305 $Y=5.397
+ $X2=3.055 $Y2=5.397
r141 99 102 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.64 $Y=3.545
+ $X2=1.64 $Y2=4.565
r142 97 158 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.64 $Y=5.245
+ $X2=1.64 $Y2=5.397
r143 97 102 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.64 $Y=5.245
+ $X2=1.64 $Y2=4.565
r144 96 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r145 95 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=5.397
+ $X2=1.64 $Y2=5.397
r146 95 96 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=1.555 $Y=5.397
+ $X2=1.205 $Y2=5.397
r147 91 156 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r148 91 93 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r149 88 154 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r150 88 90 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.015 $Y2=5.397
r151 87 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r152 87 90 0.7557 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.015 $Y2=5.397
r153 83 154 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r154 83 85 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r155 81 165 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=5.245 $X2=7.815 $Y2=5.33
r156 81 146 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=5.245 $X2=7.135 $Y2=5.33
r157 81 138 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=5.245 $X2=6.455 $Y2=5.33
r158 81 130 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=5.245 $X2=5.775 $Y2=5.33
r159 81 161 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=5.245 $X2=5.095 $Y2=5.33
r160 81 120 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=5.245 $X2=4.415 $Y2=5.33
r161 81 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=5.245 $X2=3.735 $Y2=5.33
r162 81 108 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=5.245 $X2=3.055 $Y2=5.33
r163 81 106 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=5.245 $X2=2.375 $Y2=5.33
r164 81 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=5.245 $X2=1.695 $Y2=5.33
r165 81 90 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=5.245 $X2=1.015 $Y2=5.33
r166 81 154 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=5.245 $X2=0.335 $Y2=5.33
r167 8 149 300 $w=1.7e-07 $l=1.46833e-06 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=2.825 $X2=7.9 $Y2=4.225
r168 7 141 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=3.565 $X2=6.95 $Y2=4.565
r169 6 133 600 $w=1.7e-07 $l=1.06066e-06 $layer=licon1_PDIFF $count=1 $X=5.965
+ $Y=3.565 $X2=6.09 $Y2=4.565
r170 5 126 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=5
+ $Y=2.825 $X2=5.14 $Y2=4.565
r171 5 123 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=5
+ $Y=2.825 $X2=5.14 $Y2=3.205
r172 4 114 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.25
+ $Y=2.825 $X2=3.39 $Y2=4.565
r173 4 111 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=3.25
+ $Y=2.825 $X2=3.39 $Y2=3.545
r174 3 102 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=2.825 $X2=1.64 $Y2=4.565
r175 3 99 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=2.825 $X2=1.64 $Y2=3.545
r176 2 93 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=3.565 $X2=1.12 $Y2=4.565
r177 1 85 600 $w=1.7e-07 $l=1.06066e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.565
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%SN 3 7 9 11 14 17 21 25 31 36 37 39 44
c131 31 0 7.745e-20 $X=6.86 $Y=1.22
r132 37 39 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.465 $Y=1.22
+ $X2=0.32 $Y2=1.22
r133 36 44 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.715 $Y=1.22
+ $X2=6.86 $Y2=1.22
r134 36 37 6.01801 $w=1.7e-07 $l=6.25e-06 $layer=MET1_cond $X=6.715 $Y=1.22
+ $X2=0.465 $Y2=1.22
r135 31 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.86 $Y=1.22
+ $X2=6.86 $Y2=1.22
r136 31 34 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.86 $Y=1.22
+ $X2=6.86 $Y2=1.37
r137 25 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=1.22
+ $X2=0.32 $Y2=1.22
r138 25 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.22
+ $X2=0.32 $Y2=1.59
r139 23 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.37 $X2=6.86 $Y2=1.37
r140 21 23 19.4984 $w=3.09e-07 $l=1.25e-07 $layer=POLY_cond $X=6.735 $Y=1.37
+ $X2=6.86 $Y2=1.37
r141 20 21 10.9191 $w=3.09e-07 $l=7e-08 $layer=POLY_cond $X=6.665 $Y=1.37
+ $X2=6.735 $Y2=1.37
r142 17 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.59 $X2=0.32 $Y2=1.59
r143 17 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.59
+ $X2=0.367 $Y2=1.755
r144 17 18 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.59
+ $X2=0.367 $Y2=1.425
r145 12 21 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.535
+ $X2=6.735 $Y2=1.37
r146 12 14 1363.96 $w=1.5e-07 $l=2.66e-06 $layer=POLY_cond $X=6.735 $Y=1.535
+ $X2=6.735 $Y2=4.195
r147 9 20 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.665 $Y=1.205
+ $X2=6.665 $Y2=1.37
r148 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.665 $Y=1.205
+ $X2=6.665 $Y2=0.835
r149 7 19 1251.15 $w=1.5e-07 $l=2.44e-06 $layer=POLY_cond $X=0.475 $Y=4.195
+ $X2=0.475 $Y2=1.755
r150 3 18 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.425
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%A_152_89# 1 3 11 15 21 26 27 28 29 30 32
+ 35 39 44
c86 44 0 1.71621e-19 $X=2.507 $Y=1.155
c87 27 0 1.29912e-19 $X=2.33 $Y=1.505
r88 43 44 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.507 $Y=0.985
+ $X2=2.507 $Y2=1.155
r89 39 41 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=2.515 $Y=3.205
+ $X2=2.515 $Y2=4.565
r90 37 39 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=2.515 $Y=3.01
+ $X2=2.515 $Y2=3.205
r91 35 43 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=2.515 $Y=0.865
+ $X2=2.515 $Y2=0.985
r92 32 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.415 $Y=1.42
+ $X2=2.415 $Y2=1.155
r93 29 37 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.345 $Y=2.925
+ $X2=2.515 $Y2=3.01
r94 29 30 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.345 $Y=2.925
+ $X2=1.115 $Y2=2.925
r95 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=1.505
+ $X2=2.415 $Y2=1.42
r96 27 28 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.33 $Y=1.505
+ $X2=1.115 $Y2=1.505
r97 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=2.84
+ $X2=1.115 $Y2=2.925
r98 24 26 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.03 $Y=2.84
+ $X2=1.03 $Y2=2.045
r99 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=1.59
+ $X2=1.115 $Y2=1.505
r100 23 26 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.03 $Y=1.59
+ $X2=1.03 $Y2=2.045
r101 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=2.045 $X2=1.03 $Y2=2.045
r102 19 21 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.905 $Y=2.045
+ $X2=1.03 $Y2=2.045
r103 17 19 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.835 $Y=2.045
+ $X2=0.905 $Y2=2.045
r104 13 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.21
+ $X2=0.905 $Y2=2.045
r105 13 15 1017.84 $w=1.5e-07 $l=1.985e-06 $layer=POLY_cond $X=0.905 $Y=2.21
+ $X2=0.905 $Y2=4.195
r106 9 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=1.88
+ $X2=0.835 $Y2=2.045
r107 9 11 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=0.835 $Y=1.88
+ $X2=0.835 $Y2=0.835
r108 3 41 240 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=2.825 $X2=2.515 $Y2=4.565
r109 3 39 240 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=2.825 $X2=2.515 $Y2=3.205
r110 1 35 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.575 $X2=2.515 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%D 3 7 10 14 19
c41 19 0 1.41836e-19 $X=1.915 $Y=1.96
c42 10 0 1.12321e-19 $X=1.915 $Y=1.96
r43 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.915 $Y=1.96
+ $X2=1.915 $Y2=1.96
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.96 $X2=1.915 $Y2=1.96
r45 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.96
+ $X2=1.915 $Y2=2.125
r46 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.96
+ $X2=1.915 $Y2=1.795
r47 7 12 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=1.855 $Y=3.825
+ $X2=1.855 $Y2=2.125
r48 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.855 $Y=0.945
+ $X2=1.855 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c218 55 0 6.79641e-20 $X=4.11 $Y=2.33
c219 48 0 1.98654e-19 $X=2.755 $Y=1.59
c220 44 0 1.86602e-19 $X=2.67 $Y=2.33
c221 30 0 1.29912e-19 $X=2.755 $Y=1.425
c222 25 0 1.41836e-19 $X=2.275 $Y=2.505
r223 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.65 $Y=2.33
+ $X2=4.505 $Y2=2.33
r224 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.355 $Y=2.33
+ $X2=5.5 $Y2=2.33
r225 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=5.355 $Y=2.33
+ $X2=4.65 $Y2=2.33
r226 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.42 $Y=2.33
+ $X2=2.275 $Y2=2.33
r227 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.36 $Y=2.33
+ $X2=4.505 $Y2=2.33
r228 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=4.36 $Y=2.33
+ $X2=2.42 $Y2=2.33
r229 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.505 $Y=2.33
+ $X2=4.505 $Y2=2.33
r230 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.505 $Y=2.33
+ $X2=4.505 $Y2=2.505
r231 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.275 $Y=2.33
+ $X2=2.275 $Y2=2.33
r232 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.275 $Y=2.33
+ $X2=2.275 $Y2=2.505
r233 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.5 $Y=2.33 $X2=5.5
+ $Y2=2.33
r234 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.5 $Y=2.33
+ $X2=5.5 $Y2=2.505
r235 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.33
+ $X2=4.505 $Y2=2.33
r236 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.42 $Y=2.33
+ $X2=4.11 $Y2=2.33
r237 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=2.245
+ $X2=4.11 $Y2=2.33
r238 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.025 $Y=2.245
+ $X2=4.025 $Y2=1.59
r239 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.755 $Y=2.245
+ $X2=2.755 $Y2=1.59
r240 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.33
+ $X2=2.275 $Y2=2.33
r241 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.67 $Y=2.33
+ $X2=2.755 $Y2=2.245
r242 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.67 $Y=2.33
+ $X2=2.36 $Y2=2.33
r243 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=2.505 $X2=5.5 $Y2=2.505
r244 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=5.382 $Y=1.425
+ $X2=5.382 $Y2=1.575
r245 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=2.505 $X2=4.505 $Y2=2.505
r246 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=2.505
+ $X2=4.505 $Y2=2.67
r247 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.59 $X2=4.025 $Y2=1.59
r248 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.59
+ $X2=4.025 $Y2=1.425
r249 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.59 $X2=2.755 $Y2=1.59
r250 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.59
+ $X2=2.755 $Y2=1.425
r251 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=2.505 $X2=2.275 $Y2=2.505
r252 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=2.505
+ $X2=2.275 $Y2=2.67
r253 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=5.41 $Y=2.34
+ $X2=5.457 $Y2=2.505
r254 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=5.41 $Y=2.34
+ $X2=5.41 $Y2=1.575
r255 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=5.355 $Y=2.67
+ $X2=5.457 $Y2=2.505
r256 18 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=5.355 $Y=2.67
+ $X2=5.355 $Y2=3.825
r257 17 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.355 $Y=0.945
+ $X2=5.355 $Y2=1.425
r258 13 39 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=4.565 $Y=3.825
+ $X2=4.565 $Y2=2.67
r259 10 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.965 $Y=0.945
+ $X2=3.965 $Y2=1.425
r260 7 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.815 $Y=0.945
+ $X2=2.815 $Y2=1.425
r261 3 27 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=2.215 $Y=3.825
+ $X2=2.215 $Y2=2.67
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%A_27_115# 1 3 11 15 17 18 21 22 27 31 33
+ 37 43 46 53 54 55 60
c129 54 0 1.35571e-19 $X=3.11 $Y=1.59
c130 43 0 1.5821e-19 $X=3.345 $Y=2.505
c131 31 0 6.36774e-20 $X=3.605 $Y=3.825
c132 22 0 1.86602e-19 $X=3.25 $Y=2.505
c133 21 0 6.79641e-20 $X=3.53 $Y=2.505
c134 15 0 6.36774e-20 $X=3.175 $Y=3.825
r135 55 57 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.59
+ $X2=0.69 $Y2=1.59
r136 54 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.11 $Y=1.59
+ $X2=3.255 $Y2=1.59
r137 54 55 2.19056 $w=1.7e-07 $l=2.275e-06 $layer=MET1_cond $X=3.11 $Y=1.59
+ $X2=0.835 $Y2=1.59
r138 51 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.255 $Y=1.59
+ $X2=3.255 $Y2=1.59
r139 51 53 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=3.255 $Y=1.55
+ $X2=3.345 $Y2=1.55
r140 46 48 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.26 $Y=0.74
+ $X2=0.26 $Y2=0.88
r141 41 53 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=1.675
+ $X2=3.345 $Y2=1.55
r142 41 43 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.345 $Y=1.675
+ $X2=3.345 $Y2=2.505
r143 37 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.59
+ $X2=0.69 $Y2=1.59
r144 37 39 194.091 $w=1.68e-07 $l=2.975e-06 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.69 $Y2=4.565
r145 35 37 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=0.69 $Y=0.965
+ $X2=0.69 $Y2=1.59
r146 34 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.88
+ $X2=0.26 $Y2=0.88
r147 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=0.88
+ $X2=0.69 $Y2=0.965
r148 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.88
+ $X2=0.345 $Y2=0.88
r149 29 31 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=3.605 $Y=2.64
+ $X2=3.605 $Y2=3.825
r150 25 27 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.605 $Y=1.455
+ $X2=3.605 $Y2=0.945
r151 24 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=2.505 $X2=3.345 $Y2=2.505
r152 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=2.505
+ $X2=3.345 $Y2=2.505
r153 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.53 $Y=2.505
+ $X2=3.605 $Y2=2.64
r154 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=2.505
+ $X2=3.345 $Y2=2.505
r155 20 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.59 $X2=3.345 $Y2=1.59
r156 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=1.59
+ $X2=3.345 $Y2=1.59
r157 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.53 $Y=1.59
+ $X2=3.605 $Y2=1.455
r158 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=1.59
+ $X2=3.345 $Y2=1.59
r159 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=2.64
+ $X2=3.25 $Y2=2.505
r160 13 15 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=3.175 $Y=2.64
+ $X2=3.175 $Y2=3.825
r161 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=1.455
+ $X2=3.25 $Y2=1.59
r162 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.175 $Y=1.455
+ $X2=3.175 $Y2=0.945
r163 3 39 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.565 $X2=0.69 $Y2=4.565
r164 1 46 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%A_428_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c187 35 0 1.98654e-19 $X=2.335 $Y=1.5
c188 18 0 1.12321e-19 $X=2.815 $Y=3.825
r189 66 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=2.925
+ $X2=5.845 $Y2=2.925
r190 62 64 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=1.99
+ $X2=5.845 $Y2=1.99
r191 60 68 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.84
+ $X2=5.845 $Y2=2.925
r192 59 64 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.075
+ $X2=5.845 $Y2=1.99
r193 59 60 47.1364 $w=1.78e-07 $l=7.65e-07 $layer=LI1_cond $X=5.845 $Y=2.075
+ $X2=5.845 $Y2=2.84
r194 55 57 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=5.57 $Y=3.205
+ $X2=5.57 $Y2=4.565
r195 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=3.01
+ $X2=5.57 $Y2=2.925
r196 53 55 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.57 $Y=3.01
+ $X2=5.57 $Y2=3.205
r197 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.905
+ $X2=5.57 $Y2=1.99
r198 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.675
+ $X2=5.57 $Y2=1.59
r199 51 52 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.57 $Y=1.675
+ $X2=5.57 $Y2=1.905
r200 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.505
+ $X2=5.57 $Y2=1.59
r201 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.57 $Y=1.505
+ $X2=5.57 $Y2=0.865
r202 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=1.59
+ $X2=5.57 $Y2=1.59
r203 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.485 $Y=1.59
+ $X2=4.505 $Y2=1.59
r204 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=1.59 $X2=4.505 $Y2=1.59
r205 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.59
+ $X2=4.505 $Y2=1.755
r206 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.59
+ $X2=4.505 $Y2=1.425
r207 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.215 $Y=1.5
+ $X2=2.335 $Y2=1.5
r208 32 41 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.565 $Y=0.945
+ $X2=4.565 $Y2=1.425
r209 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.445 $Y=1.965
+ $X2=4.445 $Y2=1.755
r210 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=2.04
+ $X2=3.965 $Y2=2.04
r211 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.37 $Y=2.04
+ $X2=4.445 $Y2=1.965
r212 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.37 $Y=2.04
+ $X2=4.04 $Y2=2.04
r213 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.965 $Y=2.115
+ $X2=3.965 $Y2=2.04
r214 22 24 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=3.965 $Y=2.115
+ $X2=3.965 $Y2=3.825
r215 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.89 $Y=2.04
+ $X2=2.815 $Y2=2.04
r216 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.89 $Y=2.04
+ $X2=3.965 $Y2=2.04
r217 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.89 $Y=2.04 $X2=2.89
+ $Y2=2.04
r218 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.815 $Y=2.115
+ $X2=2.815 $Y2=2.04
r219 16 18 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=2.815 $Y=2.115
+ $X2=2.815 $Y2=3.825
r220 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.74 $Y=2.04
+ $X2=2.815 $Y2=2.04
r221 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.74 $Y=2.04
+ $X2=2.41 $Y2=2.04
r222 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.335 $Y=1.965
+ $X2=2.41 $Y2=2.04
r223 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.335 $Y=1.575
+ $X2=2.335 $Y2=1.5
r224 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.335 $Y=1.575
+ $X2=2.335 $Y2=1.965
r225 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.215 $Y=1.425
+ $X2=2.215 $Y2=1.5
r226 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.215 $Y=1.425
+ $X2=2.215 $Y2=0.945
r227 3 57 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=5.43
+ $Y=2.825 $X2=5.57 $Y2=4.565
r228 3 55 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=5.43
+ $Y=2.825 $X2=5.57 $Y2=3.205
r229 1 49 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.575 $X2=5.57 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%A_970_89# 1 3 11 15 23 26 28 32 33 35 36
+ 37 38 40 44 47 50 54 58 62 63 64 69
c165 37 0 8.77106e-20 $X=7.66 $Y=2.595
c166 36 0 7.745e-20 $X=7.66 $Y=1.54
c167 32 0 2.20654e-19 $X=7.57 $Y=1.93
r168 64 66 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.13 $Y=1.93
+ $X2=4.985 $Y2=1.93
r169 63 69 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.425 $Y=1.93
+ $X2=7.57 $Y2=1.93
r170 63 64 2.20982 $w=1.7e-07 $l=2.295e-06 $layer=MET1_cond $X=7.425 $Y=1.93
+ $X2=5.13 $Y2=1.93
r171 58 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.09 $Y=0.74
+ $X2=6.09 $Y2=0.91
r172 54 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.57 $Y=1.93
+ $X2=7.57 $Y2=1.93
r173 52 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=1.93
+ $X2=6.52 $Y2=1.93
r174 52 54 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=6.605 $Y=1.93
+ $X2=7.57 $Y2=1.93
r175 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.015
+ $X2=6.52 $Y2=1.93
r176 48 50 166.364 $w=1.68e-07 $l=2.55e-06 $layer=LI1_cond $X=6.52 $Y=2.015
+ $X2=6.52 $Y2=4.565
r177 47 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.845
+ $X2=6.52 $Y2=1.93
r178 46 47 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=6.52 $Y=0.995
+ $X2=6.52 $Y2=1.845
r179 45 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.91
+ $X2=6.09 $Y2=0.91
r180 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.435 $Y=0.91
+ $X2=6.52 $Y2=0.995
r181 44 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.435 $Y=0.91
+ $X2=6.175 $Y2=0.91
r182 40 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.985 $Y=1.93
+ $X2=4.985 $Y2=1.93
r183 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=2.595
+ $X2=7.66 $Y2=2.745
r184 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=1.39 $X2=7.66
+ $Y2=1.54
r185 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.635 $Y=2.095
+ $X2=7.635 $Y2=2.595
r186 33 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.635 $Y=1.765
+ $X2=7.635 $Y2=1.54
r187 32 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=1.93 $X2=7.57 $Y2=1.93
r188 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=1.93
+ $X2=7.572 $Y2=2.095
r189 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=1.93
+ $X2=7.572 $Y2=1.765
r190 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.93 $X2=4.985 $Y2=1.93
r191 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.93
+ $X2=4.985 $Y2=2.095
r192 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.93
+ $X2=4.985 $Y2=1.765
r193 26 38 347.04 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=7.685 $Y=3.825
+ $X2=7.685 $Y2=2.745
r194 23 35 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.685 $Y=0.945
+ $X2=7.685 $Y2=1.39
r195 15 30 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=4.925 $Y=3.825
+ $X2=4.925 $Y2=2.095
r196 11 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4.925 $Y=0.945
+ $X2=4.925 $Y2=1.765
r197 3 50 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=3.565 $X2=6.52 $Y2=4.565
r198 1 58 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.965
+ $Y=0.575 $X2=6.09 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%A_808_115# 1 3 11 15 20 25 26 27 28 29
+ 32 36 41 45 46 51
c128 46 0 1.5821e-19 $X=3.83 $Y=1.59
c129 26 0 1.67294e-19 $X=4.095 $Y=1.17
c130 25 0 1.57671e-19 $X=3.685 $Y=1.59
r131 46 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.83 $Y=1.59
+ $X2=3.685 $Y2=1.59
r132 45 51 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.955 $Y=1.59
+ $X2=6.1 $Y2=1.59
r133 45 46 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=5.955 $Y=1.59
+ $X2=3.83 $Y2=1.59
r134 41 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.1 $Y=1.59 $X2=6.1
+ $Y2=1.59
r135 36 38 34.5733 $w=3.38e-07 $l=1.02e-06 $layer=LI1_cond $X=4.265 $Y=3.545
+ $X2=4.265 $Y2=4.565
r136 34 36 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=4.265 $Y=3.01
+ $X2=4.265 $Y2=3.545
r137 30 32 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=4.265 $Y=1.085
+ $X2=4.265 $Y2=0.865
r138 28 34 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=2.925
+ $X2=4.265 $Y2=3.01
r139 28 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=2.925
+ $X2=3.77 $Y2=2.925
r140 26 30 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=1.17
+ $X2=4.265 $Y2=1.085
r141 26 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=1.17
+ $X2=3.77 $Y2=1.17
r142 25 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=1.59
+ $X2=3.685 $Y2=1.59
r143 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=2.84
+ $X2=3.77 $Y2=2.925
r144 23 25 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.685 $Y=2.84
+ $X2=3.685 $Y2=1.59
r145 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=1.255
+ $X2=3.77 $Y2=1.17
r146 22 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.685 $Y=1.255
+ $X2=3.685 $Y2=1.59
r147 18 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.1
+ $Y=1.59 $X2=6.1 $Y2=1.59
r148 18 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.1 $Y=1.59
+ $X2=6.305 $Y2=1.59
r149 13 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.755
+ $X2=6.305 $Y2=1.59
r150 13 15 1251.15 $w=1.5e-07 $l=2.44e-06 $layer=POLY_cond $X=6.305 $Y=1.755
+ $X2=6.305 $Y2=4.195
r151 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.425
+ $X2=6.305 $Y2=1.59
r152 9 11 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.305 $Y=1.425
+ $X2=6.305 $Y2=0.835
r153 3 38 300 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=4.04
+ $Y=2.825 $X2=4.265 $Y2=4.565
r154 3 36 300 $w=1.7e-07 $l=8.24864e-07 $layer=licon1_PDIFF $count=2 $X=4.04
+ $Y=2.825 $X2=4.265 $Y2=3.545
r155 1 32 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.575 $X2=4.265 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c83 42 0 8.77106e-20 $X=7.475 $Y=2.7
c84 33 0 9.99996e-20 $X=7.97 $Y=2.505
c85 31 0 1.20654e-19 $X=7.97 $Y=1.59
r86 40 42 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=7.47 $Y=2.7
+ $X2=7.475 $Y2=2.7
r87 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.055 $Y=2.42
+ $X2=8.055 $Y2=2.135
r88 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.055 $Y=1.675
+ $X2=8.055 $Y2=2.135
r89 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=2.505
+ $X2=8.055 $Y2=2.42
r90 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=2.505
+ $X2=7.555 $Y2=2.505
r91 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=1.59
+ $X2=8.055 $Y2=1.675
r92 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=1.59
+ $X2=7.555 $Y2=1.59
r93 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.47 $Y=2.7 $X2=7.47
+ $Y2=2.7
r94 27 29 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=7.47 $Y=2.7
+ $X2=7.47 $Y2=4.225
r95 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=2.59
+ $X2=7.555 $Y2=2.505
r96 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.47 $Y=2.59
+ $X2=7.47 $Y2=2.7
r97 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=1.505
+ $X2=7.555 $Y2=1.59
r98 21 23 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=7.47 $Y=1.505
+ $X2=7.47 $Y2=0.74
r99 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=2.135 $X2=8.055 $Y2=2.135
r100 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.135
+ $X2=8.055 $Y2=2.3
r101 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.135
+ $X2=8.055 $Y2=1.97
r102 15 20 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=8.115 $Y=3.825
+ $X2=8.115 $Y2=2.3
r103 11 19 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=8.115 $Y=0.945
+ $X2=8.115 $Y2=1.97
r104 3 29 300 $w=1.7e-07 $l=1.46116e-06 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=2.825 $X2=7.47 $Y2=4.225
r105 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFS_1%Q 1 3 11 15 18 21 25 28
r21 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=3.027
+ $X2=8.445 $Y2=3.027
r22 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.325 $Y=3.07
+ $X2=8.325 $Y2=3.07
r23 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=8.325 $Y=3.027
+ $X2=8.33 $Y2=3.027
r24 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=1.255
+ $X2=8.445 $Y2=1.255
r25 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.445 $Y=2.9
+ $X2=8.445 $Y2=3.027
r26 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=1.34
+ $X2=8.445 $Y2=1.255
r27 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=8.445 $Y=1.34
+ $X2=8.445 $Y2=2.9
r28 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.33 $Y=3.155
+ $X2=8.33 $Y2=3.027
r29 13 15 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=8.33 $Y=3.155
+ $X2=8.33 $Y2=4.225
r30 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=1.17 $X2=8.33
+ $Y2=1.255
r31 9 11 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.33 $Y=1.17 $X2=8.33
+ $Y2=0.74
r32 3 15 300 $w=1.7e-07 $l=1.46833e-06 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=2.825 $X2=8.33 $Y2=4.225
r33 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.575 $X2=8.33 $Y2=0.74
.ends

