* File: sky130_osu_sc_15T_ls__inv_1.spice
* Created: Fri Nov 12 14:57:14 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__inv_1.pex.spice"
.subckt sky130_osu_sc_15T_ls__inv_1  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_Y_M1001_d N_A_M1001_g N_GND_M1001_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PHIGHVT L=0.15 W=2
+ AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=3.068 P=7.98
pX3_noxref noxref_5 A A PROBETYPE=1
pX4_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__inv_1.pxi.spice"
*
.ends
*
*
