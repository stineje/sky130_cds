magic
tech sky130A
magscale 1 2
timestamp 1612373608
<< nwell >>
rect -9 529 374 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 252 115 282 243
<< pmos >>
rect 80 565 110 965
rect 152 565 182 965
rect 250 713 280 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 165 166 243
rect 110 131 121 165
rect 155 131 166 165
rect 110 115 166 131
rect 196 215 252 243
rect 196 131 207 215
rect 241 131 252 215
rect 196 115 252 131
rect 282 214 335 243
rect 282 131 293 214
rect 327 131 335 214
rect 282 115 335 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 565 152 965
rect 182 949 250 965
rect 182 809 193 949
rect 227 809 250 949
rect 182 713 250 809
rect 280 949 333 965
rect 280 809 291 949
rect 325 809 333 949
rect 280 713 333 809
rect 182 565 235 713
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 165
rect 207 131 241 215
rect 293 131 327 214
<< pdiffc >>
rect 35 741 69 949
rect 193 809 227 949
rect 291 809 325 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 152 965 182 991
rect 250 965 280 991
rect 80 533 110 565
rect 56 517 110 533
rect 56 483 66 517
rect 100 483 110 517
rect 56 467 110 483
rect 56 318 86 467
rect 152 419 182 565
rect 136 409 202 419
rect 136 375 152 409
rect 186 375 202 409
rect 136 365 202 375
rect 56 268 110 318
rect 80 243 110 268
rect 166 243 196 365
rect 250 357 280 713
rect 250 341 306 357
rect 252 307 262 341
rect 296 307 306 341
rect 252 271 306 307
rect 252 243 282 271
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
<< polycont >>
rect 66 483 100 517
rect 152 375 186 409
rect 262 307 296 341
<< locali >>
rect 0 1089 374 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 374 1089
rect 35 949 69 965
rect 193 949 227 1049
rect 193 793 227 809
rect 291 949 325 965
rect 35 699 69 741
rect 291 699 325 809
rect 35 665 325 699
rect 66 517 100 597
rect 66 467 100 483
rect 152 523 162 557
rect 152 409 186 523
rect 152 359 186 375
rect 223 341 257 449
rect 291 409 325 665
rect 223 307 262 341
rect 296 307 312 341
rect 35 215 241 249
rect 35 115 69 131
rect 121 165 155 181
rect 121 61 155 131
rect 207 115 241 131
rect 293 214 327 227
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 66 597 100 631
rect 162 523 196 557
rect 223 449 257 483
rect 291 375 325 409
rect 293 227 327 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 374 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 374 1089
rect 0 1049 374 1055
rect 54 631 112 637
rect 54 597 66 631
rect 100 597 134 631
rect 54 591 112 597
rect 150 557 208 563
rect 150 523 162 557
rect 196 523 230 557
rect 150 517 208 523
rect 211 483 269 489
rect 189 449 223 483
rect 257 449 269 483
rect 211 443 269 449
rect 279 409 337 415
rect 279 375 291 409
rect 325 375 337 409
rect 279 369 337 375
rect 293 267 327 369
rect 281 261 339 267
rect 281 227 293 261
rect 327 227 339 261
rect 281 221 339 227
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel viali 83 614 83 614 1 A0
port 1 n
rlabel viali 179 540 179 540 1 A1
port 2 n
rlabel viali 308 392 308 392 1 Y
port 3 n
rlabel viali 240 466 240 466 1 B0
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
