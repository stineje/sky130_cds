* File: sky130_osu_sc_15T_ms__addf_l.pxi.spice
* Created: Fri Nov 12 14:39:38 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%GND N_GND_M1009_d N_GND_M1025_d N_GND_M1022_d
+ N_GND_M1020_s N_GND_M1003_d N_GND_M1009_b N_GND_c_14_p N_GND_c_15_p
+ N_GND_c_3_p N_GND_c_4_p N_GND_c_20_p N_GND_c_54_p N_GND_c_26_p N_GND_c_24_p
+ N_GND_c_137_p N_GND_c_108_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%GND
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%VDD N_VDD_M1017_d N_VDD_M1004_d N_VDD_M1027_d
+ N_VDD_M1016_s N_VDD_M1007_d N_VDD_M1017_b N_VDD_c_181_p N_VDD_c_182_p
+ N_VDD_c_185_p N_VDD_c_186_p N_VDD_c_193_p N_VDD_c_212_p N_VDD_c_196_p
+ N_VDD_c_197_p N_VDD_c_245_p N_VDD_c_233_p N_VDD_c_234_p VDD N_VDD_c_183_p
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%VDD
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%A N_A_M1009_g N_A_M1017_g N_A_c_288_n
+ N_A_M1025_g N_A_c_334_n N_A_M1004_g N_A_c_292_n N_A_c_294_n N_A_c_295_n
+ N_A_c_296_n N_A_c_297_n N_A_M1019_g N_A_c_341_n N_A_M1026_g N_A_M1003_g
+ N_A_M1007_g N_A_c_298_n N_A_c_299_n N_A_c_303_n N_A_c_304_n N_A_c_308_n
+ N_A_c_309_n N_A_c_311_n N_A_c_315_n N_A_c_316_n N_A_c_317_n N_A_c_318_n
+ N_A_c_320_n N_A_c_322_n N_A_c_324_n N_A_c_325_n N_A_c_326_n A N_A_c_328_n
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%A
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%B N_B_M1001_g N_B_M1006_g N_B_M1024_g
+ N_B_M1000_g N_B_M1022_g N_B_M1027_g N_B_M1014_g N_B_M1023_g N_B_c_513_n
+ N_B_c_514_n N_B_c_515_n N_B_c_516_n N_B_c_517_n N_B_c_518_n N_B_c_519_n
+ N_B_c_520_n N_B_c_521_n N_B_c_522_n N_B_c_523_n N_B_c_524_n B N_B_c_525_n
+ N_B_c_526_n N_B_c_527_n N_B_c_528_n PM_SKY130_OSU_SC_15T_MS__ADDF_L%B
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%CI N_CI_M1002_g N_CI_M1008_g N_CI_M1012_g
+ N_CI_M1018_g N_CI_M1005_g N_CI_M1010_g N_CI_c_737_n N_CI_c_738_n N_CI_c_739_n
+ N_CI_c_740_n N_CI_c_741_n N_CI_c_742_n N_CI_c_743_n N_CI_c_744_n N_CI_c_745_n
+ N_CI_c_746_n N_CI_c_747_n CI N_CI_c_749_n PM_SKY130_OSU_SC_15T_MS__ADDF_L%CI
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%CON N_CON_M1002_d N_CON_M1008_d N_CON_c_907_n
+ N_CON_M1013_g N_CON_M1021_g N_CON_M1020_g N_CON_M1016_g N_CON_c_914_n
+ N_CON_c_915_n N_CON_c_916_n N_CON_c_947_n N_CON_c_920_n N_CON_c_921_n
+ N_CON_c_922_n N_CON_c_923_n N_CON_c_952_n N_CON_c_924_n N_CON_c_925_n
+ N_CON_c_927_n N_CON_c_931_n N_CON_c_933_n N_CON_c_936_n CON
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%CON
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_784_115# N_A_784_115#_M1013_d
+ N_A_784_115#_M1021_d N_A_784_115#_M1015_g N_A_784_115#_M1011_g
+ N_A_784_115#_c_1098_n N_A_784_115#_c_1099_n N_A_784_115#_c_1100_n
+ N_A_784_115#_c_1101_n N_A_784_115#_c_1114_n N_A_784_115#_c_1115_n
+ N_A_784_115#_c_1118_n N_A_784_115#_c_1102_n N_A_784_115#_c_1121_n
+ N_A_784_115#_c_1103_n N_A_784_115#_c_1106_n
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_784_115#
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_27_565# N_A_27_565#_M1017_s
+ N_A_27_565#_M1006_d N_A_27_565#_c_1217_n N_A_27_565#_c_1220_n
+ N_A_27_565#_c_1222_n PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_27_565#
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_526_565# N_A_526_565#_M1026_d
+ N_A_526_565#_M1018_d N_A_526_565#_c_1230_n N_A_526_565#_c_1233_n
+ N_A_526_565#_c_1235_n PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_526_565#
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%S N_S_M1015_d N_S_M1011_d N_S_c_1244_n
+ N_S_c_1251_n N_S_c_1249_n N_S_c_1250_n N_S_c_1256_n S
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%S
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%CO N_CO_M1020_d N_CO_M1016_d N_CO_c_1296_n CO
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%CO
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_27_115# N_A_27_115#_M1009_s
+ N_A_27_115#_M1001_d N_A_27_115#_c_1313_n N_A_27_115#_c_1316_n
+ N_A_27_115#_c_1327_n N_A_27_115#_c_1318_n
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_27_115#
x_PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_526_115# N_A_526_115#_M1019_d
+ N_A_526_115#_M1012_d N_A_526_115#_c_1333_n N_A_526_115#_c_1338_n
+ N_A_526_115#_c_1340_n N_A_526_115#_c_1341_n
+ PM_SKY130_OSU_SC_15T_MS__ADDF_L%A_526_115#
cc_1 N_GND_M1009_b N_A_M1017_g 0.0637211f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_2 N_GND_M1009_b N_A_c_288_n 0.0173144f $X=-0.045 $Y=0 $X2=2.125 $Y2=1.425
cc_3 N_GND_c_3_p N_A_c_288_n 0.0063578f $X=2.255 $Y=0.152 $X2=2.125 $Y2=1.425
cc_4 N_GND_c_4_p N_A_c_288_n 0.0042622f $X=2.34 $Y=0.74 $X2=2.125 $Y2=1.425
cc_5 N_GND_c_5_p N_A_c_288_n 0.00478641f $X=6.46 $Y=0.19 $X2=2.125 $Y2=1.425
cc_6 N_GND_M1009_b N_A_c_292_n 0.00927148f $X=-0.045 $Y=0 $X2=2.36 $Y2=1.5
cc_7 N_GND_c_4_p N_A_c_292_n 0.00269245f $X=2.34 $Y=0.74 $X2=2.36 $Y2=1.5
cc_8 N_GND_M1009_b N_A_c_294_n 0.0080793f $X=-0.045 $Y=0 $X2=2.2 $Y2=1.5
cc_9 N_GND_M1009_b N_A_c_295_n 0.00539004f $X=-0.045 $Y=0 $X2=2.36 $Y2=2.625
cc_10 N_GND_M1009_b N_A_c_296_n 0.00610054f $X=-0.045 $Y=0 $X2=2.2 $Y2=2.625
cc_11 N_GND_M1009_b N_A_c_297_n 0.0423913f $X=-0.045 $Y=0 $X2=2.435 $Y2=2.55
cc_12 N_GND_M1009_b N_A_c_298_n 0.0324507f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.59
cc_13 N_GND_M1009_b N_A_c_299_n 0.0266765f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.425
cc_14 N_GND_c_14_p N_A_c_299_n 0.00640094f $X=0.605 $Y=0.152 $X2=0.485 $Y2=1.425
cc_15 N_GND_c_15_p N_A_c_299_n 0.00411218f $X=0.69 $Y=0.74 $X2=0.485 $Y2=1.425
cc_16 N_GND_c_5_p N_A_c_299_n 0.0048006f $X=6.46 $Y=0.19 $X2=0.485 $Y2=1.425
cc_17 N_GND_M1009_b N_A_c_303_n 0.0213093f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.5
cc_18 N_GND_M1009_b N_A_c_304_n 0.0181429f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.425
cc_19 N_GND_c_4_p N_A_c_304_n 0.00404553f $X=2.34 $Y=0.74 $X2=2.495 $Y2=1.425
cc_20 N_GND_c_20_p N_A_c_304_n 0.0063578f $X=3.115 $Y=0.152 $X2=2.495 $Y2=1.425
cc_21 N_GND_c_5_p N_A_c_304_n 0.00478641f $X=6.46 $Y=0.19 $X2=2.495 $Y2=1.425
cc_22 N_GND_M1009_b N_A_c_308_n 0.0092911f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.625
cc_23 N_GND_M1009_b N_A_c_309_n 0.0285814f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.59
cc_24 N_GND_c_24_p N_A_c_309_n 0.00152586f $X=5.31 $Y=0.74 $X2=5.155 $Y2=1.59
cc_25 N_GND_M1009_b N_A_c_311_n 0.0189719f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.425
cc_26 N_GND_c_26_p N_A_c_311_n 0.0063578f $X=5.225 $Y=0.152 $X2=5.155 $Y2=1.425
cc_27 N_GND_c_24_p N_A_c_311_n 0.00496483f $X=5.31 $Y=0.74 $X2=5.155 $Y2=1.425
cc_28 N_GND_c_5_p N_A_c_311_n 0.00478641f $X=6.46 $Y=0.19 $X2=5.155 $Y2=1.425
cc_29 N_GND_M1009_b N_A_c_315_n 0.0401101f $X=-0.045 $Y=0 $X2=5.13 $Y2=2.515
cc_30 N_GND_M1009_b N_A_c_316_n 0.011447f $X=-0.045 $Y=0 $X2=5.13 $Y2=2.665
cc_31 N_GND_M1009_b N_A_c_317_n 0.0100075f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.59
cc_32 N_GND_M1009_b N_A_c_318_n 0.0025848f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.59
cc_33 N_GND_c_4_p N_A_c_318_n 0.00404679f $X=2.34 $Y=0.74 $X2=2.495 $Y2=1.59
cc_34 N_GND_M1009_b N_A_c_320_n 0.00463768f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.59
cc_35 N_GND_c_24_p N_A_c_320_n 0.00405692f $X=5.31 $Y=0.74 $X2=5.155 $Y2=1.59
cc_36 N_GND_M1009_b N_A_c_322_n 0.015289f $X=-0.045 $Y=0 $X2=2.35 $Y2=1.59
cc_37 N_GND_c_4_p N_A_c_322_n 4.76205e-19 $X=2.34 $Y=0.74 $X2=2.35 $Y2=1.59
cc_38 N_GND_M1009_b N_A_c_324_n 0.00354071f $X=-0.045 $Y=0 $X2=0.63 $Y2=1.59
cc_39 N_GND_M1009_b N_A_c_325_n 0.0199945f $X=-0.045 $Y=0 $X2=5.01 $Y2=1.59
cc_40 N_GND_M1009_b N_A_c_326_n 0.00110006f $X=-0.045 $Y=0 $X2=2.64 $Y2=1.59
cc_41 N_GND_c_4_p N_A_c_326_n 2.14981e-19 $X=2.34 $Y=0.74 $X2=2.64 $Y2=1.59
cc_42 N_GND_M1009_b N_A_c_328_n 0.00220872f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.59
cc_43 N_GND_c_24_p N_A_c_328_n 2.21784e-19 $X=5.31 $Y=0.74 $X2=5.155 $Y2=1.59
cc_44 N_GND_M1009_b N_B_M1001_g 0.0614047f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.945
cc_45 N_GND_c_15_p N_B_M1001_g 0.00385579f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.945
cc_46 N_GND_c_3_p N_B_M1001_g 0.0063578f $X=2.255 $Y=0.152 $X2=0.905 $Y2=0.945
cc_47 N_GND_c_5_p N_B_M1001_g 0.00478641f $X=6.46 $Y=0.19 $X2=0.905 $Y2=0.945
cc_48 N_GND_M1009_b N_B_M1024_g 0.0477186f $X=-0.045 $Y=0 $X2=1.765 $Y2=0.945
cc_49 N_GND_c_3_p N_B_M1024_g 0.0063578f $X=2.255 $Y=0.152 $X2=1.765 $Y2=0.945
cc_50 N_GND_c_5_p N_B_M1024_g 0.00478641f $X=6.46 $Y=0.19 $X2=1.765 $Y2=0.945
cc_51 N_GND_M1009_b N_B_M1000_g 0.0177314f $X=-0.045 $Y=0 $X2=1.765 $Y2=3.825
cc_52 N_GND_M1009_b N_B_M1022_g 0.0215112f $X=-0.045 $Y=0 $X2=2.985 $Y2=0.945
cc_53 N_GND_c_20_p N_B_M1022_g 0.0063578f $X=3.115 $Y=0.152 $X2=2.985 $Y2=0.945
cc_54 N_GND_c_54_p N_B_M1022_g 0.00385579f $X=3.2 $Y=0.74 $X2=2.985 $Y2=0.945
cc_55 N_GND_c_5_p N_B_M1022_g 0.00478641f $X=6.46 $Y=0.19 $X2=2.985 $Y2=0.945
cc_56 N_GND_M1009_b N_B_M1027_g 0.0416759f $X=-0.045 $Y=0 $X2=2.985 $Y2=3.825
cc_57 N_GND_M1009_b N_B_M1014_g 0.050864f $X=-0.045 $Y=0 $X2=4.275 $Y2=0.945
cc_58 N_GND_c_26_p N_B_M1014_g 0.00452019f $X=5.225 $Y=0.152 $X2=4.275 $Y2=0.945
cc_59 N_GND_c_5_p N_B_M1014_g 0.00478641f $X=6.46 $Y=0.19 $X2=4.275 $Y2=0.945
cc_60 N_GND_M1009_b N_B_M1023_g 0.00794292f $X=-0.045 $Y=0 $X2=4.275 $Y2=3.825
cc_61 N_GND_M1009_b N_B_c_513_n 0.020418f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.5
cc_62 N_GND_M1009_b N_B_c_514_n 0.0408357f $X=-0.045 $Y=0 $X2=2.015 $Y2=2.17
cc_63 N_GND_M1009_b N_B_c_515_n 0.0261851f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.645
cc_64 N_GND_M1009_b N_B_c_516_n 0.0239449f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.33
cc_65 N_GND_M1009_b N_B_c_517_n 0.00747922f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.5
cc_66 N_GND_M1009_b N_B_c_518_n 0.00586424f $X=-0.045 $Y=0 $X2=2.305 $Y2=2.33
cc_67 N_GND_M1009_b N_B_c_519_n 0.00729369f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.645
cc_68 N_GND_M1009_b N_B_c_520_n 0.00316881f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.33
cc_69 N_GND_M1009_b N_B_c_521_n 0.00291156f $X=-0.045 $Y=0 $X2=0.485 $Y2=2.33
cc_70 N_GND_M1009_b N_B_c_522_n 0.00462048f $X=-0.045 $Y=0 $X2=2.015 $Y2=2.17
cc_71 N_GND_M1009_b N_B_c_523_n 0.0254763f $X=-0.045 $Y=0 $X2=2.16 $Y2=2.33
cc_72 N_GND_M1009_b N_B_c_524_n 0.0127164f $X=-0.045 $Y=0 $X2=0.63 $Y2=2.33
cc_73 N_GND_M1009_b N_B_c_525_n 0.011565f $X=-0.045 $Y=0 $X2=2.83 $Y2=2.33
cc_74 N_GND_M1009_b N_B_c_526_n 0.00467059f $X=-0.045 $Y=0 $X2=2.45 $Y2=2.33
cc_75 N_GND_M1009_b N_B_c_527_n 0.00762182f $X=-0.045 $Y=0 $X2=4.06 $Y2=2.332
cc_76 N_GND_M1009_b N_B_c_528_n 0.019513f $X=-0.045 $Y=0 $X2=3.67 $Y2=2.332
cc_77 N_GND_M1009_b N_CI_M1002_g 0.0366615f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.945
cc_78 N_GND_c_3_p N_CI_M1002_g 0.0063578f $X=2.255 $Y=0.152 $X2=1.335 $Y2=0.945
cc_79 N_GND_c_5_p N_CI_M1002_g 0.00478641f $X=6.46 $Y=0.19 $X2=1.335 $Y2=0.945
cc_80 N_GND_M1009_b N_CI_M1008_g 0.0255405f $X=-0.045 $Y=0 $X2=1.335 $Y2=3.825
cc_81 N_GND_M1009_b N_CI_M1012_g 0.0516995f $X=-0.045 $Y=0 $X2=3.415 $Y2=0.945
cc_82 N_GND_c_54_p N_CI_M1012_g 0.00385579f $X=3.2 $Y=0.74 $X2=3.415 $Y2=0.945
cc_83 N_GND_c_26_p N_CI_M1012_g 0.0063578f $X=5.225 $Y=0.152 $X2=3.415 $Y2=0.945
cc_84 N_GND_c_5_p N_CI_M1012_g 0.00478641f $X=6.46 $Y=0.19 $X2=3.415 $Y2=0.945
cc_85 N_GND_M1009_b N_CI_M1018_g 0.00805841f $X=-0.045 $Y=0 $X2=3.415 $Y2=3.825
cc_86 N_GND_M1009_b N_CI_M1005_g 0.0444321f $X=-0.045 $Y=0 $X2=4.685 $Y2=0.945
cc_87 N_GND_c_26_p N_CI_M1005_g 0.0063578f $X=5.225 $Y=0.152 $X2=4.685 $Y2=0.945
cc_88 N_GND_c_5_p N_CI_M1005_g 0.00478641f $X=6.46 $Y=0.19 $X2=4.685 $Y2=0.945
cc_89 N_GND_M1009_b N_CI_M1010_g 0.0180089f $X=-0.045 $Y=0 $X2=4.685 $Y2=3.825
cc_90 N_GND_M1009_b N_CI_c_737_n 0.0263087f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.96
cc_91 N_GND_M1009_b N_CI_c_738_n 0.0265765f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.33
cc_92 N_GND_M1009_b N_CI_c_739_n 0.027099f $X=-0.045 $Y=0 $X2=4.745 $Y2=2.14
cc_93 N_GND_M1009_b N_CI_c_740_n 4.344e-19 $X=-0.045 $Y=0 $X2=1.325 $Y2=1.96
cc_94 N_GND_M1009_b N_CI_c_741_n 0.0034786f $X=-0.045 $Y=0 $X2=3.415 $Y2=1.96
cc_95 N_GND_M1009_b N_CI_c_742_n 0.00482822f $X=-0.045 $Y=0 $X2=4.745 $Y2=1.96
cc_96 N_GND_M1009_b N_CI_c_743_n 0.00272047f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.33
cc_97 N_GND_M1009_b N_CI_c_744_n 0.0145621f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.96
cc_98 N_GND_M1009_b N_CI_c_745_n 0.00159337f $X=-0.045 $Y=0 $X2=1.47 $Y2=1.96
cc_99 N_GND_M1009_b N_CI_c_746_n 0.0148915f $X=-0.045 $Y=0 $X2=4.6 $Y2=1.96
cc_100 N_GND_M1009_b N_CI_c_747_n 0.00231544f $X=-0.045 $Y=0 $X2=3.56 $Y2=1.96
cc_101 N_GND_M1009_b CI 0.0120192f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.96
cc_102 N_GND_M1009_b N_CI_c_749_n 0.00618156f $X=-0.045 $Y=0 $X2=4.745 $Y2=1.96
cc_103 N_GND_M1009_b N_CON_c_907_n 0.0180088f $X=-0.045 $Y=0 $X2=3.845 $Y2=1.425
cc_104 N_GND_c_26_p N_CON_c_907_n 0.0063578f $X=5.225 $Y=0.152 $X2=3.845
+ $Y2=1.425
cc_105 N_GND_c_5_p N_CON_c_907_n 0.00478641f $X=6.46 $Y=0.19 $X2=3.845 $Y2=1.425
cc_106 N_GND_M1009_b N_CON_M1021_g 0.0372583f $X=-0.045 $Y=0 $X2=3.845 $Y2=3.825
cc_107 N_GND_M1009_b N_CON_M1020_g 0.105191f $X=-0.045 $Y=0 $X2=6.535 $Y2=0.835
cc_108 N_GND_c_108_p N_CON_M1020_g 0.0067724f $X=6.32 $Y=0.74 $X2=6.535
+ $Y2=0.835
cc_109 N_GND_c_5_p N_CON_M1020_g 0.00481485f $X=6.46 $Y=0.19 $X2=6.535 $Y2=0.835
cc_110 N_GND_M1009_b N_CON_c_914_n 0.0252876f $X=-0.045 $Y=0 $X2=3.845 $Y2=1.59
cc_111 N_GND_M1009_b N_CON_c_915_n 0.0356508f $X=-0.045 $Y=0 $X2=6.41 $Y2=2.48
cc_112 N_GND_M1009_b N_CON_c_916_n 0.00417041f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.74
cc_113 N_GND_c_3_p N_CON_c_916_n 0.00779312f $X=2.255 $Y=0.152 $X2=1.55 $Y2=0.74
cc_114 N_GND_c_4_p N_CON_c_916_n 0.00114036f $X=2.34 $Y=0.74 $X2=1.55 $Y2=0.74
cc_115 N_GND_c_5_p N_CON_c_916_n 0.00478039f $X=6.46 $Y=0.19 $X2=1.55 $Y2=0.74
cc_116 N_GND_M1009_b N_CON_c_920_n 0.00911049f $X=-0.045 $Y=0 $X2=1.665
+ $Y2=2.765
cc_117 N_GND_M1009_b N_CON_c_921_n 0.00107881f $X=-0.045 $Y=0 $X2=3.97 $Y2=1.22
cc_118 N_GND_M1009_b N_CON_c_922_n 0.0107538f $X=-0.045 $Y=0 $X2=6.41 $Y2=2.48
cc_119 N_GND_M1009_b N_CON_c_923_n 0.00462698f $X=-0.045 $Y=0 $X2=1.665
+ $Y2=1.505
cc_120 N_GND_M1009_b N_CON_c_924_n 0.00289677f $X=-0.045 $Y=0 $X2=3.97 $Y2=1.59
cc_121 N_GND_M1009_b N_CON_c_925_n 0.0123826f $X=-0.045 $Y=0 $X2=6.41 $Y2=1.22
cc_122 N_GND_c_108_p N_CON_c_925_n 0.0104315f $X=6.32 $Y=0.74 $X2=6.41 $Y2=1.22
cc_123 N_GND_M1025_d N_CON_c_927_n 0.00593744f $X=2.2 $Y=0.575 $X2=3.825
+ $Y2=1.22
cc_124 N_GND_M1022_d N_CON_c_927_n 0.00244115f $X=3.06 $Y=0.575 $X2=3.825
+ $Y2=1.22
cc_125 N_GND_c_4_p N_CON_c_927_n 0.0173894f $X=2.34 $Y=0.74 $X2=3.825 $Y2=1.22
cc_126 N_GND_c_54_p N_CON_c_927_n 0.00128152f $X=3.2 $Y=0.74 $X2=3.825 $Y2=1.22
cc_127 N_GND_M1009_b N_CON_c_931_n 5.54826e-19 $X=-0.045 $Y=0 $X2=1.695 $Y2=1.22
cc_128 N_GND_c_4_p N_CON_c_931_n 5.67165e-19 $X=2.34 $Y=0.74 $X2=1.695 $Y2=1.22
cc_129 N_GND_M1003_d N_CON_c_933_n 0.00887784f $X=5.17 $Y=0.575 $X2=5.995
+ $Y2=1.22
cc_130 N_GND_M1009_b N_CON_c_933_n 0.0146888f $X=-0.045 $Y=0 $X2=5.995 $Y2=1.22
cc_131 N_GND_c_24_p N_CON_c_933_n 0.0186277f $X=5.31 $Y=0.74 $X2=5.995 $Y2=1.22
cc_132 N_GND_M1009_b N_CON_c_936_n 4.50048e-19 $X=-0.045 $Y=0 $X2=4.115 $Y2=1.22
cc_133 N_GND_M1009_b CON 0.0206412f $X=-0.045 $Y=0 $X2=6.14 $Y2=1.22
cc_134 N_GND_c_108_p CON 0.00140294f $X=6.32 $Y=0.74 $X2=6.14 $Y2=1.22
cc_135 N_GND_M1009_b N_A_784_115#_M1015_g 0.0861907f $X=-0.045 $Y=0 $X2=5.585
+ $Y2=0.835
cc_136 N_GND_c_24_p N_A_784_115#_M1015_g 0.00981172f $X=5.31 $Y=0.74 $X2=5.585
+ $Y2=0.835
cc_137 N_GND_c_137_p N_A_784_115#_M1015_g 0.00644441f $X=6.235 $Y=0.152
+ $X2=5.585 $Y2=0.835
cc_138 N_GND_c_108_p N_A_784_115#_M1015_g 0.00460621f $X=6.32 $Y=0.74 $X2=5.585
+ $Y2=0.835
cc_139 N_GND_c_5_p N_A_784_115#_M1015_g 0.00481485f $X=6.46 $Y=0.19 $X2=5.585
+ $Y2=0.835
cc_140 N_GND_M1009_b N_A_784_115#_c_1098_n 0.0268831f $X=-0.045 $Y=0 $X2=5.585
+ $Y2=2.495
cc_141 N_GND_M1009_b N_A_784_115#_c_1099_n 0.00887593f $X=-0.045 $Y=0 $X2=3.845
+ $Y2=2.77
cc_142 N_GND_M1009_b N_A_784_115#_c_1100_n 0.00593307f $X=-0.045 $Y=0 $X2=4.225
+ $Y2=1.96
cc_143 N_GND_M1009_b N_A_784_115#_c_1101_n 9.19767e-19 $X=-0.045 $Y=0 $X2=3.93
+ $Y2=1.96
cc_144 N_GND_M1009_b N_A_784_115#_c_1102_n 0.00483243f $X=-0.045 $Y=0 $X2=4.31
+ $Y2=1.875
cc_145 N_GND_M1009_b N_A_784_115#_c_1103_n 0.00155336f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=0.74
cc_146 N_GND_c_26_p N_A_784_115#_c_1103_n 0.0140069f $X=5.225 $Y=0.152 $X2=4.06
+ $Y2=0.74
cc_147 N_GND_c_5_p N_A_784_115#_c_1103_n 0.0112943f $X=6.46 $Y=0.19 $X2=4.06
+ $Y2=0.74
cc_148 N_GND_M1009_b N_A_784_115#_c_1106_n 0.00798748f $X=-0.045 $Y=0 $X2=5.415
+ $Y2=2.495
cc_149 N_GND_M1009_b N_S_c_1244_n 0.0198074f $X=-0.045 $Y=0 $X2=5.8 $Y2=0.74
cc_150 N_GND_c_24_p N_S_c_1244_n 0.0175944f $X=5.31 $Y=0.74 $X2=5.8 $Y2=0.74
cc_151 N_GND_c_137_p N_S_c_1244_n 0.00736239f $X=6.235 $Y=0.152 $X2=5.8 $Y2=0.74
cc_152 N_GND_c_108_p N_S_c_1244_n 0.0140971f $X=6.32 $Y=0.74 $X2=5.8 $Y2=0.74
cc_153 N_GND_c_5_p N_S_c_1244_n 0.00476261f $X=6.46 $Y=0.19 $X2=5.8 $Y2=0.74
cc_154 N_GND_M1009_b N_S_c_1249_n 0.0135159f $X=-0.045 $Y=0 $X2=5.925 $Y2=2.905
cc_155 N_GND_M1009_b N_S_c_1250_n 0.0121999f $X=-0.045 $Y=0 $X2=5.925 $Y2=1.96
cc_156 N_GND_M1009_b N_CO_c_1296_n 0.0789044f $X=-0.045 $Y=0 $X2=6.75 $Y2=0.74
cc_157 N_GND_c_5_p N_CO_c_1296_n 0.00476261f $X=6.46 $Y=0.19 $X2=6.75 $Y2=0.74
cc_158 N_GND_M1009_b CO 0.00667411f $X=-0.045 $Y=0 $X2=6.75 $Y2=2.7
cc_159 N_GND_M1009_b N_A_27_115#_c_1313_n 0.00156074f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_160 N_GND_c_14_p N_A_27_115#_c_1313_n 0.00736644f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_161 N_GND_c_5_p N_A_27_115#_c_1313_n 0.00476377f $X=6.46 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_162 N_GND_M1009_d N_A_27_115#_c_1316_n 0.00400988f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.175
cc_163 N_GND_c_15_p N_A_27_115#_c_1316_n 0.012242f $X=0.69 $Y=0.74 $X2=1.035
+ $Y2=1.175
cc_164 N_GND_M1009_b N_A_27_115#_c_1318_n 0.00158657f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.74
cc_165 N_GND_c_15_p N_A_27_115#_c_1318_n 2.23682e-19 $X=0.69 $Y=0.74 $X2=1.12
+ $Y2=0.74
cc_166 N_GND_c_3_p N_A_27_115#_c_1318_n 0.00776503f $X=2.255 $Y=0.152 $X2=1.12
+ $Y2=0.74
cc_167 N_GND_c_5_p N_A_27_115#_c_1318_n 0.00478269f $X=6.46 $Y=0.19 $X2=1.12
+ $Y2=0.74
cc_168 N_GND_M1009_b N_A_526_115#_c_1333_n 0.00158657f $X=-0.045 $Y=0 $X2=2.77
+ $Y2=0.74
cc_169 N_GND_c_4_p N_A_526_115#_c_1333_n 2.23682e-19 $X=2.34 $Y=0.74 $X2=2.77
+ $Y2=0.74
cc_170 N_GND_c_20_p N_A_526_115#_c_1333_n 0.00797933f $X=3.115 $Y=0.152 $X2=2.77
+ $Y2=0.74
cc_171 N_GND_c_54_p N_A_526_115#_c_1333_n 2.23682e-19 $X=3.2 $Y=0.74 $X2=2.77
+ $Y2=0.74
cc_172 N_GND_c_5_p N_A_526_115#_c_1333_n 0.00478269f $X=6.46 $Y=0.19 $X2=2.77
+ $Y2=0.74
cc_173 N_GND_M1022_d N_A_526_115#_c_1338_n 0.00465706f $X=3.06 $Y=0.575
+ $X2=3.545 $Y2=1.175
cc_174 N_GND_c_54_p N_A_526_115#_c_1338_n 0.011349f $X=3.2 $Y=0.74 $X2=3.545
+ $Y2=1.175
cc_175 N_GND_c_4_p N_A_526_115#_c_1340_n 0.00262623f $X=2.34 $Y=0.74 $X2=2.855
+ $Y2=1.175
cc_176 N_GND_M1009_b N_A_526_115#_c_1341_n 0.00158657f $X=-0.045 $Y=0 $X2=3.63
+ $Y2=0.74
cc_177 N_GND_c_54_p N_A_526_115#_c_1341_n 2.23682e-19 $X=3.2 $Y=0.74 $X2=3.63
+ $Y2=0.74
cc_178 N_GND_c_26_p N_A_526_115#_c_1341_n 0.00776503f $X=5.225 $Y=0.152 $X2=3.63
+ $Y2=0.74
cc_179 N_GND_c_5_p N_A_526_115#_c_1341_n 0.00478269f $X=6.46 $Y=0.19 $X2=3.63
+ $Y2=0.74
cc_180 N_VDD_M1017_b N_A_M1017_g 0.0296275f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_181 N_VDD_c_181_p N_A_M1017_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_182 N_VDD_c_182_p N_A_M1017_g 0.00354579f $X=0.69 $Y=3.895 $X2=0.475
+ $Y2=3.825
cc_183 N_VDD_c_183_p N_A_M1017_g 0.00429146f $X=6.46 $Y=5.36 $X2=0.475 $Y2=3.825
cc_184 N_VDD_M1017_b N_A_c_334_n 0.0168245f $X=-0.045 $Y=2.645 $X2=2.125 $Y2=2.7
cc_185 N_VDD_c_185_p N_A_c_334_n 0.00496961f $X=2.255 $Y=5.397 $X2=2.125 $Y2=2.7
cc_186 N_VDD_c_186_p N_A_c_334_n 0.00354579f $X=2.34 $Y=3.555 $X2=2.125 $Y2=2.7
cc_187 N_VDD_c_183_p N_A_c_334_n 0.00429146f $X=6.46 $Y=5.36 $X2=2.125 $Y2=2.7
cc_188 N_VDD_M1017_b N_A_c_295_n 0.00301031f $X=-0.045 $Y=2.645 $X2=2.36
+ $Y2=2.625
cc_189 N_VDD_c_186_p N_A_c_295_n 0.00274574f $X=2.34 $Y=3.555 $X2=2.36 $Y2=2.625
cc_190 N_VDD_M1017_b N_A_c_296_n 0.00180595f $X=-0.045 $Y=2.645 $X2=2.2
+ $Y2=2.625
cc_191 N_VDD_M1017_b N_A_c_341_n 0.0175567f $X=-0.045 $Y=2.645 $X2=2.555 $Y2=2.7
cc_192 N_VDD_c_186_p N_A_c_341_n 0.00354579f $X=2.34 $Y=3.555 $X2=2.555 $Y2=2.7
cc_193 N_VDD_c_193_p N_A_c_341_n 0.00496961f $X=3.115 $Y=5.397 $X2=2.555 $Y2=2.7
cc_194 N_VDD_c_183_p N_A_c_341_n 0.00429146f $X=6.46 $Y=5.36 $X2=2.555 $Y2=2.7
cc_195 N_VDD_M1017_b N_A_M1007_g 0.0207392f $X=-0.045 $Y=2.645 $X2=5.095
+ $Y2=3.825
cc_196 N_VDD_c_196_p N_A_M1007_g 0.00503522f $X=5.225 $Y=5.397 $X2=5.095
+ $Y2=3.825
cc_197 N_VDD_c_197_p N_A_M1007_g 0.0039779f $X=5.31 $Y=3.895 $X2=5.095 $Y2=3.825
cc_198 N_VDD_c_183_p N_A_M1007_g 0.00431676f $X=6.46 $Y=5.36 $X2=5.095 $Y2=3.825
cc_199 N_VDD_M1017_b N_A_c_308_n 0.0037377f $X=-0.045 $Y=2.645 $X2=2.555
+ $Y2=2.625
cc_200 N_VDD_M1017_b N_A_c_316_n 0.0032155f $X=-0.045 $Y=2.645 $X2=5.13
+ $Y2=2.665
cc_201 N_VDD_M1017_b N_B_M1006_g 0.0198657f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_202 N_VDD_c_182_p N_B_M1006_g 0.00354579f $X=0.69 $Y=3.895 $X2=0.905
+ $Y2=3.825
cc_203 N_VDD_c_185_p N_B_M1006_g 0.00496961f $X=2.255 $Y=5.397 $X2=0.905
+ $Y2=3.825
cc_204 N_VDD_c_183_p N_B_M1006_g 0.00429146f $X=6.46 $Y=5.36 $X2=0.905 $Y2=3.825
cc_205 N_VDD_M1017_b N_B_M1000_g 0.0197066f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=3.825
cc_206 N_VDD_c_185_p N_B_M1000_g 0.00503522f $X=2.255 $Y=5.397 $X2=1.765
+ $Y2=3.825
cc_207 N_VDD_c_186_p N_B_M1000_g 0.00294885f $X=2.34 $Y=3.555 $X2=1.765
+ $Y2=3.825
cc_208 N_VDD_c_183_p N_B_M1000_g 0.00431676f $X=6.46 $Y=5.36 $X2=1.765 $Y2=3.825
cc_209 N_VDD_M1017_b N_B_M1027_g 0.0216181f $X=-0.045 $Y=2.645 $X2=2.985
+ $Y2=3.825
cc_210 N_VDD_c_186_p N_B_M1027_g 4.9048e-19 $X=2.34 $Y=3.555 $X2=2.985 $Y2=3.825
cc_211 N_VDD_c_193_p N_B_M1027_g 0.00503522f $X=3.115 $Y=5.397 $X2=2.985
+ $Y2=3.825
cc_212 N_VDD_c_212_p N_B_M1027_g 0.00378444f $X=3.2 $Y=3.895 $X2=2.985 $Y2=3.825
cc_213 N_VDD_c_183_p N_B_M1027_g 0.00431676f $X=6.46 $Y=5.36 $X2=2.985 $Y2=3.825
cc_214 N_VDD_M1017_b N_B_M1023_g 0.0212968f $X=-0.045 $Y=2.645 $X2=4.275
+ $Y2=3.825
cc_215 N_VDD_c_196_p N_B_M1023_g 0.00503522f $X=5.225 $Y=5.397 $X2=4.275
+ $Y2=3.825
cc_216 N_VDD_c_183_p N_B_M1023_g 0.00431675f $X=6.46 $Y=5.36 $X2=4.275 $Y2=3.825
cc_217 N_VDD_M1017_b N_B_c_513_n 0.00479818f $X=-0.045 $Y=2.645 $X2=0.895
+ $Y2=2.5
cc_218 N_VDD_M1017_b N_CI_M1008_g 0.0215563f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=3.825
cc_219 N_VDD_c_182_p N_CI_M1008_g 4.9048e-19 $X=0.69 $Y=3.895 $X2=1.335
+ $Y2=3.825
cc_220 N_VDD_c_185_p N_CI_M1008_g 0.00503522f $X=2.255 $Y=5.397 $X2=1.335
+ $Y2=3.825
cc_221 N_VDD_c_183_p N_CI_M1008_g 0.00431676f $X=6.46 $Y=5.36 $X2=1.335
+ $Y2=3.825
cc_222 N_VDD_M1017_b N_CI_M1018_g 0.0215058f $X=-0.045 $Y=2.645 $X2=3.415
+ $Y2=3.825
cc_223 N_VDD_c_212_p N_CI_M1018_g 0.00378444f $X=3.2 $Y=3.895 $X2=3.415
+ $Y2=3.825
cc_224 N_VDD_c_196_p N_CI_M1018_g 0.00503522f $X=5.225 $Y=5.397 $X2=3.415
+ $Y2=3.825
cc_225 N_VDD_c_183_p N_CI_M1018_g 0.00431676f $X=6.46 $Y=5.36 $X2=3.415
+ $Y2=3.825
cc_226 N_VDD_M1017_b N_CI_M1010_g 0.021076f $X=-0.045 $Y=2.645 $X2=4.685
+ $Y2=3.825
cc_227 N_VDD_c_196_p N_CI_M1010_g 0.00503522f $X=5.225 $Y=5.397 $X2=4.685
+ $Y2=3.825
cc_228 N_VDD_c_183_p N_CI_M1010_g 0.00431675f $X=6.46 $Y=5.36 $X2=4.685
+ $Y2=3.825
cc_229 N_VDD_M1017_b N_CON_M1021_g 0.0194185f $X=-0.045 $Y=2.645 $X2=3.845
+ $Y2=3.825
cc_230 N_VDD_c_196_p N_CON_M1021_g 0.00503522f $X=5.225 $Y=5.397 $X2=3.845
+ $Y2=3.825
cc_231 N_VDD_c_183_p N_CON_M1021_g 0.00431676f $X=6.46 $Y=5.36 $X2=3.845
+ $Y2=3.825
cc_232 N_VDD_M1017_b N_CON_M1016_g 0.0785026f $X=-0.045 $Y=2.645 $X2=6.535
+ $Y2=4.195
cc_233 N_VDD_c_233_p N_CON_M1016_g 0.00752104f $X=6.32 $Y=4.235 $X2=6.535
+ $Y2=4.195
cc_234 N_VDD_c_234_p N_CON_M1016_g 0.00503522f $X=6.46 $Y=5.33 $X2=6.535
+ $Y2=4.195
cc_235 N_VDD_c_183_p N_CON_M1016_g 0.00431676f $X=6.46 $Y=5.36 $X2=6.535
+ $Y2=4.195
cc_236 N_VDD_M1017_b N_CON_c_915_n 0.00643378f $X=-0.045 $Y=2.645 $X2=6.41
+ $Y2=2.48
cc_237 N_VDD_M1017_b N_CON_c_947_n 0.00198641f $X=-0.045 $Y=2.645 $X2=1.55
+ $Y2=3.555
cc_238 N_VDD_c_185_p N_CON_c_947_n 0.00455459f $X=2.255 $Y=5.397 $X2=1.55
+ $Y2=3.555
cc_239 N_VDD_c_183_p N_CON_c_947_n 0.00434939f $X=6.46 $Y=5.36 $X2=1.55
+ $Y2=3.555
cc_240 N_VDD_M1017_b N_CON_c_920_n 0.00146295f $X=-0.045 $Y=2.645 $X2=1.665
+ $Y2=2.765
cc_241 N_VDD_M1017_b N_CON_c_922_n 0.00545748f $X=-0.045 $Y=2.645 $X2=6.41
+ $Y2=2.48
cc_242 N_VDD_M1017_b N_CON_c_952_n 0.00251676f $X=-0.045 $Y=2.645 $X2=1.665
+ $Y2=2.857
cc_243 N_VDD_M1017_b N_A_784_115#_M1011_g 0.0692472f $X=-0.045 $Y=2.645
+ $X2=5.585 $Y2=4.195
cc_244 N_VDD_c_197_p N_A_784_115#_M1011_g 0.0135052f $X=5.31 $Y=3.895 $X2=5.585
+ $Y2=4.195
cc_245 N_VDD_c_245_p N_A_784_115#_M1011_g 0.00503522f $X=6.235 $Y=5.397
+ $X2=5.585 $Y2=4.195
cc_246 N_VDD_c_233_p N_A_784_115#_M1011_g 0.00486385f $X=6.32 $Y=4.235 $X2=5.585
+ $Y2=4.195
cc_247 N_VDD_c_183_p N_A_784_115#_M1011_g 0.00431675f $X=6.46 $Y=5.36 $X2=5.585
+ $Y2=4.195
cc_248 N_VDD_M1017_b N_A_784_115#_c_1098_n 0.00469272f $X=-0.045 $Y=2.645
+ $X2=5.585 $Y2=2.495
cc_249 N_VDD_M1017_b N_A_784_115#_c_1099_n 0.00257504f $X=-0.045 $Y=2.645
+ $X2=3.845 $Y2=2.77
cc_250 N_VDD_M1017_b N_A_784_115#_c_1114_n 0.00427075f $X=-0.045 $Y=2.645
+ $X2=4.06 $Y2=3.16
cc_251 N_VDD_M1017_b N_A_784_115#_c_1115_n 0.00198641f $X=-0.045 $Y=2.645
+ $X2=4.06 $Y2=3.555
cc_252 N_VDD_c_196_p N_A_784_115#_c_1115_n 0.00475585f $X=5.225 $Y=5.397
+ $X2=4.06 $Y2=3.555
cc_253 N_VDD_c_183_p N_A_784_115#_c_1115_n 0.00434939f $X=6.46 $Y=5.36 $X2=4.06
+ $Y2=3.555
cc_254 N_VDD_M1007_d N_A_784_115#_c_1118_n 0.00919791f $X=5.17 $Y=2.825 $X2=5.33
+ $Y2=3.075
cc_255 N_VDD_M1017_b N_A_784_115#_c_1118_n 0.00388557f $X=-0.045 $Y=2.645
+ $X2=5.33 $Y2=3.075
cc_256 N_VDD_c_197_p N_A_784_115#_c_1118_n 0.0064526f $X=5.31 $Y=3.895 $X2=5.33
+ $Y2=3.075
cc_257 N_VDD_M1007_d N_A_784_115#_c_1121_n 0.00259083f $X=5.17 $Y=2.825
+ $X2=5.415 $Y2=2.99
cc_258 N_VDD_M1017_b N_A_784_115#_c_1121_n 0.00416996f $X=-0.045 $Y=2.645
+ $X2=5.415 $Y2=2.99
cc_259 N_VDD_M1017_b N_A_784_115#_c_1106_n 6.65464e-19 $X=-0.045 $Y=2.645
+ $X2=5.415 $Y2=2.495
cc_260 N_VDD_M1017_b N_A_27_565#_c_1217_n 0.00199838f $X=-0.045 $Y=2.645
+ $X2=0.26 $Y2=3.555
cc_261 N_VDD_c_181_p N_A_27_565#_c_1217_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.555
cc_262 N_VDD_c_183_p N_A_27_565#_c_1217_n 0.00435496f $X=6.46 $Y=5.36 $X2=0.26
+ $Y2=3.555
cc_263 N_VDD_M1017_d N_A_27_565#_c_1220_n 0.005567f $X=0.55 $Y=2.825 $X2=1.035
+ $Y2=3.2
cc_264 N_VDD_c_182_p N_A_27_565#_c_1220_n 0.0077616f $X=0.69 $Y=3.895 $X2=1.035
+ $Y2=3.2
cc_265 N_VDD_M1017_b N_A_27_565#_c_1222_n 0.00198641f $X=-0.045 $Y=2.645
+ $X2=1.12 $Y2=3.555
cc_266 N_VDD_c_185_p N_A_27_565#_c_1222_n 0.0045126f $X=2.255 $Y=5.397 $X2=1.12
+ $Y2=3.555
cc_267 N_VDD_c_183_p N_A_27_565#_c_1222_n 0.00434939f $X=6.46 $Y=5.36 $X2=1.12
+ $Y2=3.555
cc_268 N_VDD_M1017_b N_A_526_565#_c_1230_n 0.00198641f $X=-0.045 $Y=2.645
+ $X2=2.77 $Y2=3.555
cc_269 N_VDD_c_193_p N_A_526_565#_c_1230_n 0.00475585f $X=3.115 $Y=5.397
+ $X2=2.77 $Y2=3.555
cc_270 N_VDD_c_183_p N_A_526_565#_c_1230_n 0.00434939f $X=6.46 $Y=5.36 $X2=2.77
+ $Y2=3.555
cc_271 N_VDD_M1027_d N_A_526_565#_c_1233_n 0.00875443f $X=3.06 $Y=2.825
+ $X2=3.545 $Y2=3.195
cc_272 N_VDD_c_212_p N_A_526_565#_c_1233_n 0.00768266f $X=3.2 $Y=3.895 $X2=3.545
+ $Y2=3.195
cc_273 N_VDD_M1017_b N_A_526_565#_c_1235_n 0.00198641f $X=-0.045 $Y=2.645
+ $X2=3.63 $Y2=3.555
cc_274 N_VDD_c_196_p N_A_526_565#_c_1235_n 0.0045126f $X=5.225 $Y=5.397 $X2=3.63
+ $Y2=3.555
cc_275 N_VDD_c_183_p N_A_526_565#_c_1235_n 0.00434939f $X=6.46 $Y=5.36 $X2=3.63
+ $Y2=3.555
cc_276 N_VDD_M1017_b N_S_c_1251_n 0.0158717f $X=-0.045 $Y=2.645 $X2=5.8
+ $Y2=3.105
cc_277 N_VDD_c_245_p N_S_c_1251_n 0.00452684f $X=6.235 $Y=5.397 $X2=5.8
+ $Y2=3.105
cc_278 N_VDD_c_233_p N_S_c_1251_n 0.0358835f $X=6.32 $Y=4.235 $X2=5.8 $Y2=3.105
cc_279 N_VDD_c_183_p N_S_c_1251_n 0.00435496f $X=6.46 $Y=5.36 $X2=5.8 $Y2=3.105
cc_280 N_VDD_M1017_b N_S_c_1249_n 0.00671597f $X=-0.045 $Y=2.645 $X2=5.925
+ $Y2=2.905
cc_281 N_VDD_M1017_b N_S_c_1256_n 0.0123513f $X=-0.045 $Y=2.645 $X2=5.925
+ $Y2=2.99
cc_282 N_VDD_M1017_b S 0.00760382f $X=-0.045 $Y=2.645 $X2=5.8 $Y2=3.105
cc_283 N_VDD_M1017_b N_CO_c_1296_n 0.0440481f $X=-0.045 $Y=2.645 $X2=6.75
+ $Y2=0.74
cc_284 N_VDD_c_234_p N_CO_c_1296_n 0.00477009f $X=6.46 $Y=5.33 $X2=6.75 $Y2=0.74
cc_285 N_VDD_c_183_p N_CO_c_1296_n 0.00435496f $X=6.46 $Y=5.36 $X2=6.75 $Y2=0.74
cc_286 N_VDD_M1017_b CO 0.0109934f $X=-0.045 $Y=2.645 $X2=6.75 $Y2=2.7
cc_287 N_A_M1017_g N_B_M1001_g 0.0285181f $X=0.475 $Y=3.825 $X2=0.905 $Y2=0.945
cc_288 N_A_c_298_n N_B_M1001_g 0.0223074f $X=0.485 $Y=1.59 $X2=0.905 $Y2=0.945
cc_289 N_A_c_299_n N_B_M1001_g 0.0282855f $X=0.485 $Y=1.425 $X2=0.905 $Y2=0.945
cc_290 N_A_c_317_n N_B_M1001_g 0.00278747f $X=0.485 $Y=1.59 $X2=0.905 $Y2=0.945
cc_291 N_A_c_322_n N_B_M1001_g 0.006033f $X=2.35 $Y=1.59 $X2=0.905 $Y2=0.945
cc_292 N_A_c_324_n N_B_M1001_g 8.6716e-19 $X=0.63 $Y=1.59 $X2=0.905 $Y2=0.945
cc_293 N_A_M1017_g N_B_M1006_g 0.0539782f $X=0.475 $Y=3.825 $X2=0.905 $Y2=3.825
cc_294 N_A_c_288_n N_B_M1024_g 0.0723172f $X=2.125 $Y=1.425 $X2=1.765 $Y2=0.945
cc_295 N_A_c_303_n N_B_M1024_g 0.00810048f $X=2.495 $Y=1.5 $X2=1.765 $Y2=0.945
cc_296 N_A_c_318_n N_B_M1024_g 0.00113262f $X=2.495 $Y=1.59 $X2=1.765 $Y2=0.945
cc_297 N_A_c_322_n N_B_M1024_g 0.0037004f $X=2.35 $Y=1.59 $X2=1.765 $Y2=0.945
cc_298 N_A_c_326_n N_B_M1024_g 5.04344e-19 $X=2.64 $Y=1.59 $X2=1.765 $Y2=0.945
cc_299 N_A_c_296_n N_B_M1000_g 0.143904f $X=2.2 $Y=2.625 $X2=1.765 $Y2=3.825
cc_300 N_A_c_297_n N_B_M1000_g 0.00269561f $X=2.435 $Y=2.55 $X2=1.765 $Y2=3.825
cc_301 N_A_c_304_n N_B_M1022_g 0.0175139f $X=2.495 $Y=1.425 $X2=2.985 $Y2=0.945
cc_302 N_A_c_297_n N_B_M1027_g 0.0223254f $X=2.435 $Y=2.55 $X2=2.985 $Y2=3.825
cc_303 N_A_c_308_n N_B_M1027_g 0.0462588f $X=2.555 $Y=2.625 $X2=2.985 $Y2=3.825
cc_304 N_A_c_325_n N_B_M1014_g 0.00122134f $X=5.01 $Y=1.59 $X2=4.275 $Y2=0.945
cc_305 N_A_M1017_g N_B_c_513_n 0.0218907f $X=0.475 $Y=3.825 $X2=0.895 $Y2=2.5
cc_306 N_A_c_294_n N_B_c_514_n 0.00301833f $X=2.2 $Y=1.5 $X2=2.015 $Y2=2.17
cc_307 N_A_c_296_n N_B_c_514_n 0.00640881f $X=2.2 $Y=2.625 $X2=2.015 $Y2=2.17
cc_308 N_A_c_297_n N_B_c_514_n 0.022133f $X=2.435 $Y=2.55 $X2=2.015 $Y2=2.17
cc_309 N_A_c_322_n N_B_c_514_n 5.24163e-19 $X=2.35 $Y=1.59 $X2=2.015 $Y2=2.17
cc_310 N_A_c_297_n N_B_c_515_n 0.00217946f $X=2.435 $Y=2.55 $X2=2.975 $Y2=1.645
cc_311 N_A_c_303_n N_B_c_515_n 0.0187158f $X=2.495 $Y=1.5 $X2=2.975 $Y2=1.645
cc_312 N_A_c_318_n N_B_c_515_n 7.65216e-19 $X=2.495 $Y=1.59 $X2=2.975 $Y2=1.645
cc_313 N_A_c_325_n N_B_c_515_n 0.0026048f $X=5.01 $Y=1.59 $X2=2.975 $Y2=1.645
cc_314 N_A_c_326_n N_B_c_515_n 8.1198e-19 $X=2.64 $Y=1.59 $X2=2.975 $Y2=1.645
cc_315 N_A_M1017_g N_B_c_517_n 4.31631e-19 $X=0.475 $Y=3.825 $X2=0.895 $Y2=2.5
cc_316 N_A_c_298_n N_B_c_517_n 8.97793e-19 $X=0.485 $Y=1.59 $X2=0.895 $Y2=2.5
cc_317 N_A_c_294_n N_B_c_518_n 0.00243929f $X=2.2 $Y=1.5 $X2=2.305 $Y2=2.33
cc_318 N_A_c_296_n N_B_c_518_n 0.00867832f $X=2.2 $Y=2.625 $X2=2.305 $Y2=2.33
cc_319 N_A_c_297_n N_B_c_518_n 0.00530786f $X=2.435 $Y=2.55 $X2=2.305 $Y2=2.33
cc_320 N_A_c_318_n N_B_c_518_n 9.1275e-19 $X=2.495 $Y=1.59 $X2=2.305 $Y2=2.33
cc_321 N_A_c_297_n N_B_c_519_n 0.00783283f $X=2.435 $Y=2.55 $X2=2.975 $Y2=1.645
cc_322 N_A_c_303_n N_B_c_519_n 9.28573e-19 $X=2.495 $Y=1.5 $X2=2.975 $Y2=1.645
cc_323 N_A_c_318_n N_B_c_519_n 0.00843011f $X=2.495 $Y=1.59 $X2=2.975 $Y2=1.645
cc_324 N_A_c_325_n N_B_c_519_n 0.0127134f $X=5.01 $Y=1.59 $X2=2.975 $Y2=1.645
cc_325 N_A_c_326_n N_B_c_519_n 0.00227634f $X=2.64 $Y=1.59 $X2=2.975 $Y2=1.645
cc_326 N_A_M1017_g N_B_c_521_n 0.0206591f $X=0.475 $Y=3.825 $X2=0.485 $Y2=2.33
cc_327 N_A_c_298_n N_B_c_521_n 3.21671e-19 $X=0.485 $Y=1.59 $X2=0.485 $Y2=2.33
cc_328 N_A_c_317_n N_B_c_521_n 0.00208589f $X=0.485 $Y=1.59 $X2=0.485 $Y2=2.33
cc_329 N_A_c_294_n N_B_c_522_n 4.19356e-19 $X=2.2 $Y=1.5 $X2=2.015 $Y2=2.17
cc_330 N_A_c_296_n N_B_c_522_n 9.92874e-19 $X=2.2 $Y=2.625 $X2=2.015 $Y2=2.17
cc_331 N_A_c_297_n N_B_c_522_n 0.00170298f $X=2.435 $Y=2.55 $X2=2.015 $Y2=2.17
cc_332 N_A_c_322_n N_B_c_522_n 0.00231345f $X=2.35 $Y=1.59 $X2=2.015 $Y2=2.17
cc_333 N_A_c_296_n N_B_c_523_n 0.00100445f $X=2.2 $Y=2.625 $X2=2.16 $Y2=2.33
cc_334 N_A_M1017_g N_B_c_524_n 0.00322062f $X=0.475 $Y=3.825 $X2=0.63 $Y2=2.33
cc_335 N_A_c_298_n N_B_c_524_n 7.14347e-19 $X=0.485 $Y=1.59 $X2=0.63 $Y2=2.33
cc_336 N_A_c_317_n N_B_c_524_n 9.8095e-19 $X=0.485 $Y=1.59 $X2=0.63 $Y2=2.33
cc_337 N_A_c_324_n N_B_c_524_n 0.003172f $X=0.63 $Y=1.59 $X2=0.63 $Y2=2.33
cc_338 N_A_c_297_n N_B_c_525_n 0.00451179f $X=2.435 $Y=2.55 $X2=2.83 $Y2=2.33
cc_339 N_A_c_308_n N_B_c_525_n 0.00349205f $X=2.555 $Y=2.625 $X2=2.83 $Y2=2.33
cc_340 N_A_c_296_n N_B_c_526_n 0.00563612f $X=2.2 $Y=2.625 $X2=2.45 $Y2=2.33
cc_341 N_A_c_297_n N_B_c_526_n 0.0049099f $X=2.435 $Y=2.55 $X2=2.45 $Y2=2.33
cc_342 N_A_c_297_n N_B_c_528_n 3.06713e-19 $X=2.435 $Y=2.55 $X2=3.67 $Y2=2.332
cc_343 N_A_c_322_n N_CI_M1002_g 0.00986519f $X=2.35 $Y=1.59 $X2=1.335 $Y2=0.945
cc_344 N_A_c_325_n N_CI_M1012_g 0.00474173f $X=5.01 $Y=1.59 $X2=3.415 $Y2=0.945
cc_345 N_A_c_311_n N_CI_M1005_g 0.0676079f $X=5.155 $Y=1.425 $X2=4.685 $Y2=0.945
cc_346 N_A_c_315_n N_CI_M1005_g 0.00809446f $X=5.13 $Y=2.515 $X2=4.685 $Y2=0.945
cc_347 N_A_c_320_n N_CI_M1005_g 0.00116181f $X=5.155 $Y=1.59 $X2=4.685 $Y2=0.945
cc_348 N_A_c_325_n N_CI_M1005_g 0.00570385f $X=5.01 $Y=1.59 $X2=4.685 $Y2=0.945
cc_349 N_A_c_328_n N_CI_M1005_g 8.57008e-19 $X=5.155 $Y=1.59 $X2=4.685 $Y2=0.945
cc_350 N_A_c_315_n N_CI_M1010_g 0.00831744f $X=5.13 $Y=2.515 $X2=4.685 $Y2=3.825
cc_351 N_A_c_316_n N_CI_M1010_g 0.125125f $X=5.13 $Y=2.665 $X2=4.685 $Y2=3.825
cc_352 N_A_c_322_n N_CI_c_737_n 0.00157267f $X=2.35 $Y=1.59 $X2=1.325 $Y2=1.96
cc_353 N_A_c_315_n N_CI_c_739_n 0.0209004f $X=5.13 $Y=2.515 $X2=4.745 $Y2=2.14
cc_354 N_A_c_325_n N_CI_c_739_n 2.31739e-19 $X=5.01 $Y=1.59 $X2=4.745 $Y2=2.14
cc_355 N_A_c_322_n N_CI_c_740_n 0.00446594f $X=2.35 $Y=1.59 $X2=1.325 $Y2=1.96
cc_356 N_A_c_325_n N_CI_c_741_n 0.00121378f $X=5.01 $Y=1.59 $X2=3.415 $Y2=1.96
cc_357 N_A_c_315_n N_CI_c_742_n 0.00385032f $X=5.13 $Y=2.515 $X2=4.745 $Y2=1.96
cc_358 N_A_c_325_n N_CI_c_742_n 0.00203847f $X=5.01 $Y=1.59 $X2=4.745 $Y2=1.96
cc_359 N_A_c_294_n N_CI_c_744_n 0.00109073f $X=2.2 $Y=1.5 $X2=3.27 $Y2=1.96
cc_360 N_A_c_297_n N_CI_c_744_n 0.00626944f $X=2.435 $Y=2.55 $X2=3.27 $Y2=1.96
cc_361 N_A_c_303_n N_CI_c_744_n 0.00232838f $X=2.495 $Y=1.5 $X2=3.27 $Y2=1.96
cc_362 N_A_c_318_n N_CI_c_744_n 0.00394572f $X=2.495 $Y=1.59 $X2=3.27 $Y2=1.96
cc_363 N_A_c_322_n N_CI_c_744_n 0.0733404f $X=2.35 $Y=1.59 $X2=3.27 $Y2=1.96
cc_364 N_A_c_325_n N_CI_c_744_n 0.0520179f $X=5.01 $Y=1.59 $X2=3.27 $Y2=1.96
cc_365 N_A_c_326_n N_CI_c_744_n 0.0266076f $X=2.64 $Y=1.59 $X2=3.27 $Y2=1.96
cc_366 N_A_c_322_n N_CI_c_745_n 0.0259568f $X=2.35 $Y=1.59 $X2=1.47 $Y2=1.96
cc_367 N_A_c_325_n N_CI_c_746_n 0.0858958f $X=5.01 $Y=1.59 $X2=4.6 $Y2=1.96
cc_368 N_A_c_325_n N_CI_c_747_n 0.0268168f $X=5.01 $Y=1.59 $X2=3.56 $Y2=1.96
cc_369 N_A_M1017_g CI 0.00555516f $X=0.475 $Y=3.825 $X2=1.325 $Y2=1.96
cc_370 N_A_c_298_n CI 0.00108997f $X=0.485 $Y=1.59 $X2=1.325 $Y2=1.96
cc_371 N_A_c_317_n CI 0.00205922f $X=0.485 $Y=1.59 $X2=1.325 $Y2=1.96
cc_372 N_A_c_322_n CI 0.0466592f $X=2.35 $Y=1.59 $X2=1.325 $Y2=1.96
cc_373 N_A_c_324_n CI 0.0210627f $X=0.63 $Y=1.59 $X2=1.325 $Y2=1.96
cc_374 N_A_c_315_n N_CI_c_749_n 0.00413683f $X=5.13 $Y=2.515 $X2=4.745 $Y2=1.96
cc_375 N_A_c_325_n N_CI_c_749_n 0.0268056f $X=5.01 $Y=1.59 $X2=4.745 $Y2=1.96
cc_376 N_A_c_325_n N_CON_c_914_n 0.00283634f $X=5.01 $Y=1.59 $X2=3.845 $Y2=1.59
cc_377 N_A_c_296_n N_CON_c_920_n 0.00127956f $X=2.2 $Y=2.625 $X2=1.665 $Y2=2.765
cc_378 N_A_c_303_n N_CON_c_920_n 0.00171426f $X=2.495 $Y=1.5 $X2=1.665 $Y2=2.765
cc_379 N_A_c_318_n N_CON_c_920_n 0.00126357f $X=2.495 $Y=1.59 $X2=1.665
+ $Y2=2.765
cc_380 N_A_c_322_n N_CON_c_920_n 0.00898724f $X=2.35 $Y=1.59 $X2=1.665 $Y2=2.765
cc_381 N_A_c_326_n N_CON_c_920_n 8.75747e-19 $X=2.64 $Y=1.59 $X2=1.665 $Y2=2.765
cc_382 N_A_c_325_n N_CON_c_921_n 6.93264e-19 $X=5.01 $Y=1.59 $X2=3.97 $Y2=1.22
cc_383 N_A_c_288_n N_CON_c_923_n 8.12393e-19 $X=2.125 $Y=1.425 $X2=1.665
+ $Y2=1.505
cc_384 N_A_c_318_n N_CON_c_923_n 0.00101586f $X=2.495 $Y=1.59 $X2=1.665
+ $Y2=1.505
cc_385 N_A_c_322_n N_CON_c_923_n 0.0122304f $X=2.35 $Y=1.59 $X2=1.665 $Y2=1.505
cc_386 N_A_c_326_n N_CON_c_923_n 8.13159e-19 $X=2.64 $Y=1.59 $X2=1.665 $Y2=1.505
cc_387 N_A_c_334_n N_CON_c_952_n 9.92167e-19 $X=2.125 $Y=2.7 $X2=1.665 $Y2=2.857
cc_388 N_A_c_325_n N_CON_c_924_n 0.0171196f $X=5.01 $Y=1.59 $X2=3.97 $Y2=1.59
cc_389 N_A_c_288_n N_CON_c_927_n 0.00956968f $X=2.125 $Y=1.425 $X2=3.825
+ $Y2=1.22
cc_390 N_A_c_292_n N_CON_c_927_n 0.00146289f $X=2.36 $Y=1.5 $X2=3.825 $Y2=1.22
cc_391 N_A_c_304_n N_CON_c_927_n 0.00790627f $X=2.495 $Y=1.425 $X2=3.825
+ $Y2=1.22
cc_392 N_A_c_318_n N_CON_c_927_n 0.00357434f $X=2.495 $Y=1.59 $X2=3.825 $Y2=1.22
cc_393 N_A_c_322_n N_CON_c_927_n 0.0546702f $X=2.35 $Y=1.59 $X2=3.825 $Y2=1.22
cc_394 N_A_c_325_n N_CON_c_927_n 0.0990817f $X=5.01 $Y=1.59 $X2=3.825 $Y2=1.22
cc_395 N_A_c_326_n N_CON_c_927_n 0.0264994f $X=2.64 $Y=1.59 $X2=3.825 $Y2=1.22
cc_396 N_A_c_288_n N_CON_c_931_n 2.65615e-19 $X=2.125 $Y=1.425 $X2=1.695
+ $Y2=1.22
cc_397 N_A_c_322_n N_CON_c_931_n 0.0250774f $X=2.35 $Y=1.59 $X2=1.695 $Y2=1.22
cc_398 N_A_c_309_n N_CON_c_933_n 0.00213677f $X=5.155 $Y=1.59 $X2=5.995 $Y2=1.22
cc_399 N_A_c_311_n N_CON_c_933_n 0.00914791f $X=5.155 $Y=1.425 $X2=5.995
+ $Y2=1.22
cc_400 N_A_c_320_n N_CON_c_933_n 0.00398656f $X=5.155 $Y=1.59 $X2=5.995 $Y2=1.22
cc_401 N_A_c_325_n N_CON_c_933_n 0.0740953f $X=5.01 $Y=1.59 $X2=5.995 $Y2=1.22
cc_402 N_A_c_328_n N_CON_c_933_n 0.026558f $X=5.155 $Y=1.59 $X2=5.995 $Y2=1.22
cc_403 N_A_c_325_n N_CON_c_936_n 0.0252794f $X=5.01 $Y=1.59 $X2=4.115 $Y2=1.22
cc_404 N_A_c_309_n N_A_784_115#_M1015_g 0.0195004f $X=5.155 $Y=1.59 $X2=5.585
+ $Y2=0.835
cc_405 N_A_c_311_n N_A_784_115#_M1015_g 0.0204525f $X=5.155 $Y=1.425 $X2=5.585
+ $Y2=0.835
cc_406 N_A_c_315_n N_A_784_115#_M1015_g 0.0266804f $X=5.13 $Y=2.515 $X2=5.585
+ $Y2=0.835
cc_407 N_A_c_320_n N_A_784_115#_M1015_g 0.00131152f $X=5.155 $Y=1.59 $X2=5.585
+ $Y2=0.835
cc_408 N_A_c_328_n N_A_784_115#_M1015_g 9.02444e-19 $X=5.155 $Y=1.59 $X2=5.585
+ $Y2=0.835
cc_409 N_A_M1007_g N_A_784_115#_M1011_g 0.0532145f $X=5.095 $Y=3.825 $X2=5.585
+ $Y2=4.195
cc_410 N_A_c_315_n N_A_784_115#_c_1098_n 0.0199271f $X=5.13 $Y=2.515 $X2=5.585
+ $Y2=2.495
cc_411 N_A_c_325_n N_A_784_115#_c_1100_n 0.0018868f $X=5.01 $Y=1.59 $X2=4.225
+ $Y2=1.96
cc_412 N_A_c_325_n N_A_784_115#_c_1101_n 7.77654e-19 $X=5.01 $Y=1.59 $X2=3.93
+ $Y2=1.96
cc_413 N_A_M1007_g N_A_784_115#_c_1118_n 0.0193311f $X=5.095 $Y=3.825 $X2=5.33
+ $Y2=3.075
cc_414 N_A_c_316_n N_A_784_115#_c_1118_n 0.0016251f $X=5.13 $Y=2.665 $X2=5.33
+ $Y2=3.075
cc_415 N_A_c_320_n N_A_784_115#_c_1102_n 0.00296302f $X=5.155 $Y=1.59 $X2=4.31
+ $Y2=1.875
cc_416 N_A_c_325_n N_A_784_115#_c_1102_n 0.0140552f $X=5.01 $Y=1.59 $X2=4.31
+ $Y2=1.875
cc_417 N_A_c_328_n N_A_784_115#_c_1102_n 0.00192851f $X=5.155 $Y=1.59 $X2=4.31
+ $Y2=1.875
cc_418 N_A_M1007_g N_A_784_115#_c_1121_n 0.00698879f $X=5.095 $Y=3.825 $X2=5.415
+ $Y2=2.99
cc_419 N_A_c_315_n N_A_784_115#_c_1106_n 0.00675793f $X=5.13 $Y=2.515 $X2=5.415
+ $Y2=2.495
cc_420 N_A_M1017_g N_A_27_565#_c_1220_n 0.0179393f $X=0.475 $Y=3.825 $X2=1.035
+ $Y2=3.2
cc_421 N_A_c_320_n N_S_c_1244_n 0.00615434f $X=5.155 $Y=1.59 $X2=5.8 $Y2=0.74
cc_422 N_A_c_328_n N_S_c_1244_n 0.00346849f $X=5.155 $Y=1.59 $X2=5.8 $Y2=0.74
cc_423 N_A_M1007_g S 2.86673e-19 $X=5.095 $Y=3.825 $X2=5.8 $Y2=3.105
cc_424 N_A_c_298_n N_A_27_115#_c_1316_n 0.00146373f $X=0.485 $Y=1.59 $X2=1.035
+ $Y2=1.175
cc_425 N_A_c_299_n N_A_27_115#_c_1316_n 0.0132827f $X=0.485 $Y=1.425 $X2=1.035
+ $Y2=1.175
cc_426 N_A_c_317_n N_A_27_115#_c_1316_n 0.0102023f $X=0.485 $Y=1.59 $X2=1.035
+ $Y2=1.175
cc_427 N_A_c_322_n N_A_27_115#_c_1316_n 0.0241923f $X=2.35 $Y=1.59 $X2=1.035
+ $Y2=1.175
cc_428 N_A_c_324_n N_A_27_115#_c_1316_n 0.00663062f $X=0.63 $Y=1.59 $X2=1.035
+ $Y2=1.175
cc_429 N_A_c_317_n N_A_27_115#_c_1327_n 0.00146727f $X=0.485 $Y=1.59 $X2=0.345
+ $Y2=1.175
cc_430 N_A_c_325_n N_A_526_115#_c_1338_n 0.00468444f $X=5.01 $Y=1.59 $X2=3.545
+ $Y2=1.175
cc_431 N_A_c_325_n N_A_526_115#_c_1340_n 0.00107807f $X=5.01 $Y=1.59 $X2=2.855
+ $Y2=1.175
cc_432 N_B_M1001_g N_CI_M1002_g 0.03238f $X=0.905 $Y=0.945 $X2=1.335 $Y2=0.945
cc_433 N_B_M1024_g N_CI_M1002_g 0.0306611f $X=1.765 $Y=0.945 $X2=1.335 $Y2=0.945
cc_434 N_B_M1001_g N_CI_M1008_g 0.0101134f $X=0.905 $Y=0.945 $X2=1.335 $Y2=3.825
cc_435 N_B_M1006_g N_CI_M1008_g 0.0383066f $X=0.905 $Y=3.825 $X2=1.335 $Y2=3.825
cc_436 N_B_c_513_n N_CI_M1008_g 0.0188528f $X=0.895 $Y=2.5 $X2=1.335 $Y2=3.825
cc_437 N_B_c_514_n N_CI_M1008_g 0.057975f $X=2.015 $Y=2.17 $X2=1.335 $Y2=3.825
cc_438 N_B_c_517_n N_CI_M1008_g 0.00162835f $X=0.895 $Y=2.5 $X2=1.335 $Y2=3.825
cc_439 N_B_c_523_n N_CI_M1008_g 0.0102981f $X=2.16 $Y=2.33 $X2=1.335 $Y2=3.825
cc_440 N_B_M1022_g N_CI_M1012_g 0.0310575f $X=2.985 $Y=0.945 $X2=3.415 $Y2=0.945
cc_441 N_B_M1027_g N_CI_M1012_g 0.0160293f $X=2.985 $Y=3.825 $X2=3.415 $Y2=0.945
cc_442 N_B_c_515_n N_CI_M1012_g 0.0199829f $X=2.975 $Y=1.645 $X2=3.415 $Y2=0.945
cc_443 N_B_c_519_n N_CI_M1012_g 0.00255874f $X=2.975 $Y=1.645 $X2=3.415
+ $Y2=0.945
cc_444 N_B_M1027_g N_CI_M1018_g 0.0624306f $X=2.985 $Y=3.825 $X2=3.415 $Y2=3.825
cc_445 N_B_M1014_g N_CI_M1005_g 0.0851559f $X=4.275 $Y=0.945 $X2=4.685 $Y2=0.945
cc_446 N_B_M1023_g N_CI_M1010_g 0.124421f $X=4.275 $Y=3.825 $X2=4.685 $Y2=3.825
cc_447 N_B_M1001_g N_CI_c_737_n 0.0219985f $X=0.905 $Y=0.945 $X2=1.325 $Y2=1.96
cc_448 N_B_M1024_g N_CI_c_737_n 0.0193664f $X=1.765 $Y=0.945 $X2=1.325 $Y2=1.96
cc_449 N_B_c_523_n N_CI_c_737_n 0.00157267f $X=2.16 $Y=2.33 $X2=1.325 $Y2=1.96
cc_450 N_B_M1027_g N_CI_c_738_n 0.0204315f $X=2.985 $Y=3.825 $X2=3.415 $Y2=2.33
cc_451 N_B_c_519_n N_CI_c_738_n 9.41528e-19 $X=2.975 $Y=1.645 $X2=3.415 $Y2=2.33
cc_452 N_B_c_528_n N_CI_c_738_n 0.0120043f $X=3.67 $Y=2.332 $X2=3.415 $Y2=2.33
cc_453 N_B_c_516_n N_CI_c_739_n 0.0208261f $X=4.265 $Y=2.33 $X2=4.745 $Y2=2.14
cc_454 N_B_c_520_n N_CI_c_739_n 0.00282159f $X=4.265 $Y=2.33 $X2=4.745 $Y2=2.14
cc_455 N_B_c_527_n N_CI_c_739_n 9.10645e-19 $X=4.06 $Y=2.332 $X2=4.745 $Y2=2.14
cc_456 N_B_M1001_g N_CI_c_740_n 0.00277751f $X=0.905 $Y=0.945 $X2=1.325 $Y2=1.96
cc_457 N_B_M1024_g N_CI_c_740_n 4.162e-19 $X=1.765 $Y=0.945 $X2=1.325 $Y2=1.96
cc_458 N_B_c_523_n N_CI_c_740_n 0.00446594f $X=2.16 $Y=2.33 $X2=1.325 $Y2=1.96
cc_459 N_B_M1027_g N_CI_c_741_n 0.00154506f $X=2.985 $Y=3.825 $X2=3.415 $Y2=1.96
cc_460 N_B_c_519_n N_CI_c_741_n 0.016155f $X=2.975 $Y=1.645 $X2=3.415 $Y2=1.96
cc_461 N_B_c_528_n N_CI_c_741_n 8.40427e-19 $X=3.67 $Y=2.332 $X2=3.415 $Y2=1.96
cc_462 N_B_M1014_g N_CI_c_742_n 0.00109484f $X=4.275 $Y=0.945 $X2=4.745 $Y2=1.96
cc_463 N_B_c_516_n N_CI_c_742_n 5.51285e-19 $X=4.265 $Y=2.33 $X2=4.745 $Y2=1.96
cc_464 N_B_c_520_n N_CI_c_742_n 0.00317294f $X=4.265 $Y=2.33 $X2=4.745 $Y2=1.96
cc_465 N_B_c_527_n N_CI_c_742_n 0.00164652f $X=4.06 $Y=2.332 $X2=4.745 $Y2=1.96
cc_466 N_B_M1027_g N_CI_c_743_n 6.79377e-19 $X=2.985 $Y=3.825 $X2=3.415 $Y2=2.33
cc_467 N_B_c_519_n N_CI_c_743_n 0.0103583f $X=2.975 $Y=1.645 $X2=3.415 $Y2=2.33
cc_468 N_B_c_528_n N_CI_c_743_n 0.0188576f $X=3.67 $Y=2.332 $X2=3.415 $Y2=2.33
cc_469 N_B_M1024_g N_CI_c_744_n 0.00219877f $X=1.765 $Y=0.945 $X2=3.27 $Y2=1.96
cc_470 N_B_M1027_g N_CI_c_744_n 0.00107346f $X=2.985 $Y=3.825 $X2=3.27 $Y2=1.96
cc_471 N_B_c_514_n N_CI_c_744_n 0.00482273f $X=2.015 $Y=2.17 $X2=3.27 $Y2=1.96
cc_472 N_B_c_515_n N_CI_c_744_n 0.00166027f $X=2.975 $Y=1.645 $X2=3.27 $Y2=1.96
cc_473 N_B_c_518_n N_CI_c_744_n 0.0023297f $X=2.305 $Y=2.33 $X2=3.27 $Y2=1.96
cc_474 N_B_c_519_n N_CI_c_744_n 0.0163564f $X=2.975 $Y=1.645 $X2=3.27 $Y2=1.96
cc_475 N_B_c_522_n N_CI_c_744_n 0.00748189f $X=2.015 $Y=2.17 $X2=3.27 $Y2=1.96
cc_476 N_B_c_523_n N_CI_c_744_n 0.055048f $X=2.16 $Y=2.33 $X2=3.27 $Y2=1.96
cc_477 N_B_c_525_n N_CI_c_744_n 0.0323265f $X=2.83 $Y=2.33 $X2=3.27 $Y2=1.96
cc_478 N_B_c_526_n N_CI_c_744_n 0.0269315f $X=2.45 $Y=2.33 $X2=3.27 $Y2=1.96
cc_479 N_B_c_528_n N_CI_c_744_n 0.0380655f $X=3.67 $Y=2.332 $X2=3.27 $Y2=1.96
cc_480 N_B_M1001_g N_CI_c_745_n 8.6716e-19 $X=0.905 $Y=0.945 $X2=1.47 $Y2=1.96
cc_481 N_B_c_523_n N_CI_c_745_n 0.0259579f $X=2.16 $Y=2.33 $X2=1.47 $Y2=1.96
cc_482 N_B_M1014_g N_CI_c_746_n 0.00112864f $X=4.275 $Y=0.945 $X2=4.6 $Y2=1.96
cc_483 N_B_c_516_n N_CI_c_746_n 0.00116782f $X=4.265 $Y=2.33 $X2=4.6 $Y2=1.96
cc_484 N_B_c_520_n N_CI_c_746_n 0.00192504f $X=4.265 $Y=2.33 $X2=4.6 $Y2=1.96
cc_485 N_B_c_527_n N_CI_c_746_n 0.062156f $X=4.06 $Y=2.332 $X2=4.6 $Y2=1.96
cc_486 N_B_c_528_n N_CI_c_746_n 0.0092809f $X=3.67 $Y=2.332 $X2=4.6 $Y2=1.96
cc_487 N_B_M1027_g N_CI_c_747_n 8.88888e-19 $X=2.985 $Y=3.825 $X2=3.56 $Y2=1.96
cc_488 N_B_c_519_n N_CI_c_747_n 0.00213923f $X=2.975 $Y=1.645 $X2=3.56 $Y2=1.96
cc_489 N_B_c_528_n N_CI_c_747_n 0.0247742f $X=3.67 $Y=2.332 $X2=3.56 $Y2=1.96
cc_490 N_B_M1001_g CI 0.00535234f $X=0.905 $Y=0.945 $X2=1.325 $Y2=1.96
cc_491 N_B_c_513_n CI 5.74814e-19 $X=0.895 $Y=2.5 $X2=1.325 $Y2=1.96
cc_492 N_B_c_517_n CI 2.90821e-19 $X=0.895 $Y=2.5 $X2=1.325 $Y2=1.96
cc_493 N_B_c_521_n CI 0.00110643f $X=0.485 $Y=2.33 $X2=1.325 $Y2=1.96
cc_494 N_B_c_523_n CI 0.0466415f $X=2.16 $Y=2.33 $X2=1.325 $Y2=1.96
cc_495 N_B_c_524_n CI 0.0211771f $X=0.63 $Y=2.33 $X2=1.325 $Y2=1.96
cc_496 N_B_M1014_g N_CI_c_749_n 4.28504e-19 $X=4.275 $Y=0.945 $X2=4.745 $Y2=1.96
cc_497 N_B_M1014_g N_CON_c_907_n 0.0294515f $X=4.275 $Y=0.945 $X2=3.845
+ $Y2=1.425
cc_498 N_B_M1014_g N_CON_M1021_g 0.0179106f $X=4.275 $Y=0.945 $X2=3.845
+ $Y2=3.825
cc_499 N_B_M1023_g N_CON_M1021_g 0.042769f $X=4.275 $Y=3.825 $X2=3.845 $Y2=3.825
cc_500 N_B_c_516_n N_CON_M1021_g 0.0211897f $X=4.265 $Y=2.33 $X2=3.845 $Y2=3.825
cc_501 N_B_c_520_n N_CON_M1021_g 4.28168e-19 $X=4.265 $Y=2.33 $X2=3.845
+ $Y2=3.825
cc_502 N_B_M1014_g N_CON_c_914_n 0.0200025f $X=4.275 $Y=0.945 $X2=3.845 $Y2=1.59
cc_503 N_B_M1024_g N_CON_c_916_n 0.00370639f $X=1.765 $Y=0.945 $X2=1.55 $Y2=0.74
cc_504 N_B_M1024_g N_CON_c_920_n 0.0112485f $X=1.765 $Y=0.945 $X2=1.665
+ $Y2=2.765
cc_505 N_B_M1000_g N_CON_c_920_n 0.0123615f $X=1.765 $Y=3.825 $X2=1.665
+ $Y2=2.765
cc_506 N_B_c_514_n N_CON_c_920_n 0.00754141f $X=2.015 $Y=2.17 $X2=1.665
+ $Y2=2.765
cc_507 N_B_c_517_n N_CON_c_920_n 0.00630121f $X=0.895 $Y=2.5 $X2=1.665 $Y2=2.765
cc_508 N_B_c_522_n N_CON_c_920_n 0.0257712f $X=2.015 $Y=2.17 $X2=1.665 $Y2=2.765
cc_509 N_B_c_523_n N_CON_c_920_n 0.0157763f $X=2.16 $Y=2.33 $X2=1.665 $Y2=2.765
cc_510 N_B_c_526_n N_CON_c_920_n 0.00105333f $X=2.45 $Y=2.33 $X2=1.665 $Y2=2.765
cc_511 N_B_M1014_g N_CON_c_921_n 0.0018911f $X=4.275 $Y=0.945 $X2=3.97 $Y2=1.22
cc_512 N_B_M1024_g N_CON_c_923_n 0.00525936f $X=1.765 $Y=0.945 $X2=1.665
+ $Y2=1.505
cc_513 N_B_M1000_g N_CON_c_952_n 0.00812165f $X=1.765 $Y=3.825 $X2=1.665
+ $Y2=2.857
cc_514 N_B_c_523_n N_CON_c_952_n 0.00503431f $X=2.16 $Y=2.33 $X2=1.665 $Y2=2.857
cc_515 N_B_M1014_g N_CON_c_924_n 7.2637e-19 $X=4.275 $Y=0.945 $X2=3.97 $Y2=1.59
cc_516 N_B_c_519_n N_CON_c_924_n 0.0022487f $X=2.975 $Y=1.645 $X2=3.97 $Y2=1.59
cc_517 N_B_M1024_g N_CON_c_927_n 0.00888363f $X=1.765 $Y=0.945 $X2=3.825
+ $Y2=1.22
cc_518 N_B_M1022_g N_CON_c_927_n 0.00137389f $X=2.985 $Y=0.945 $X2=3.825
+ $Y2=1.22
cc_519 N_B_c_515_n N_CON_c_927_n 0.00153777f $X=2.975 $Y=1.645 $X2=3.825
+ $Y2=1.22
cc_520 N_B_c_519_n N_CON_c_927_n 0.00117917f $X=2.975 $Y=1.645 $X2=3.825
+ $Y2=1.22
cc_521 N_B_M1001_g N_CON_c_931_n 3.1812e-19 $X=0.905 $Y=0.945 $X2=1.695 $Y2=1.22
cc_522 N_B_M1024_g N_CON_c_931_n 0.00131762f $X=1.765 $Y=0.945 $X2=1.695
+ $Y2=1.22
cc_523 N_B_M1014_g N_CON_c_933_n 0.00151809f $X=4.275 $Y=0.945 $X2=5.995
+ $Y2=1.22
cc_524 N_B_M1014_g N_CON_c_936_n 9.72315e-19 $X=4.275 $Y=0.945 $X2=4.115
+ $Y2=1.22
cc_525 N_B_M1014_g N_A_784_115#_c_1099_n 0.00218215f $X=4.275 $Y=0.945 $X2=3.845
+ $Y2=2.77
cc_526 N_B_M1023_g N_A_784_115#_c_1099_n 0.00502446f $X=4.275 $Y=3.825 $X2=3.845
+ $Y2=2.77
cc_527 N_B_c_516_n N_A_784_115#_c_1099_n 0.003498f $X=4.265 $Y=2.33 $X2=3.845
+ $Y2=2.77
cc_528 N_B_c_520_n N_A_784_115#_c_1099_n 0.0120274f $X=4.265 $Y=2.33 $X2=3.845
+ $Y2=2.77
cc_529 N_B_c_527_n N_A_784_115#_c_1099_n 0.0204781f $X=4.06 $Y=2.332 $X2=3.845
+ $Y2=2.77
cc_530 N_B_M1014_g N_A_784_115#_c_1100_n 0.00690261f $X=4.275 $Y=0.945 $X2=4.225
+ $Y2=1.96
cc_531 N_B_c_516_n N_A_784_115#_c_1100_n 0.00274037f $X=4.265 $Y=2.33 $X2=4.225
+ $Y2=1.96
cc_532 N_B_c_520_n N_A_784_115#_c_1100_n 0.016625f $X=4.265 $Y=2.33 $X2=4.225
+ $Y2=1.96
cc_533 N_B_c_527_n N_A_784_115#_c_1100_n 0.00247487f $X=4.06 $Y=2.332 $X2=4.225
+ $Y2=1.96
cc_534 N_B_M1023_g N_A_784_115#_c_1114_n 0.00221174f $X=4.275 $Y=3.825 $X2=4.06
+ $Y2=3.16
cc_535 N_B_c_516_n N_A_784_115#_c_1114_n 3.44204e-19 $X=4.265 $Y=2.33 $X2=4.06
+ $Y2=3.16
cc_536 N_B_c_520_n N_A_784_115#_c_1114_n 0.0015127f $X=4.265 $Y=2.33 $X2=4.06
+ $Y2=3.16
cc_537 N_B_c_527_n N_A_784_115#_c_1114_n 0.00840219f $X=4.06 $Y=2.332 $X2=4.06
+ $Y2=3.16
cc_538 N_B_M1023_g N_A_784_115#_c_1118_n 0.0162839f $X=4.275 $Y=3.825 $X2=5.33
+ $Y2=3.075
cc_539 N_B_c_520_n N_A_784_115#_c_1118_n 0.00328494f $X=4.265 $Y=2.33 $X2=5.33
+ $Y2=3.075
cc_540 N_B_c_527_n N_A_784_115#_c_1118_n 0.00471773f $X=4.06 $Y=2.332 $X2=5.33
+ $Y2=3.075
cc_541 N_B_M1014_g N_A_784_115#_c_1102_n 0.0218215f $X=4.275 $Y=0.945 $X2=4.31
+ $Y2=1.875
cc_542 N_B_M1014_g N_A_784_115#_c_1103_n 0.00727511f $X=4.275 $Y=0.945 $X2=4.06
+ $Y2=0.74
cc_543 N_B_M1006_g N_A_27_565#_c_1220_n 0.0163254f $X=0.905 $Y=3.825 $X2=1.035
+ $Y2=3.2
cc_544 N_B_c_513_n N_A_27_565#_c_1220_n 0.00110112f $X=0.895 $Y=2.5 $X2=1.035
+ $Y2=3.2
cc_545 N_B_c_517_n N_A_27_565#_c_1220_n 0.0124135f $X=0.895 $Y=2.5 $X2=1.035
+ $Y2=3.2
cc_546 N_B_c_521_n N_A_27_565#_c_1220_n 0.00457576f $X=0.485 $Y=2.33 $X2=1.035
+ $Y2=3.2
cc_547 N_B_M1027_g N_A_526_565#_c_1233_n 0.0167311f $X=2.985 $Y=3.825 $X2=3.545
+ $Y2=3.195
cc_548 N_B_c_519_n N_A_526_565#_c_1233_n 0.00240309f $X=2.975 $Y=1.645 $X2=3.545
+ $Y2=3.195
cc_549 N_B_M1001_g N_A_27_115#_c_1316_n 0.0134206f $X=0.905 $Y=0.945 $X2=1.035
+ $Y2=1.175
cc_550 N_B_M1022_g N_A_526_115#_c_1338_n 0.0123452f $X=2.985 $Y=0.945 $X2=3.545
+ $Y2=1.175
cc_551 N_B_c_515_n N_A_526_115#_c_1338_n 0.0022776f $X=2.975 $Y=1.645 $X2=3.545
+ $Y2=1.175
cc_552 N_B_c_519_n N_A_526_115#_c_1338_n 0.00811365f $X=2.975 $Y=1.645 $X2=3.545
+ $Y2=1.175
cc_553 N_B_c_515_n N_A_526_115#_c_1340_n 5.11238e-19 $X=2.975 $Y=1.645 $X2=2.855
+ $Y2=1.175
cc_554 N_CI_M1012_g N_CON_c_907_n 0.0145387f $X=3.415 $Y=0.945 $X2=3.845
+ $Y2=1.425
cc_555 N_CI_M1012_g N_CON_M1021_g 0.0190239f $X=3.415 $Y=0.945 $X2=3.845
+ $Y2=3.825
cc_556 N_CI_M1018_g N_CON_M1021_g 0.0442742f $X=3.415 $Y=3.825 $X2=3.845
+ $Y2=3.825
cc_557 N_CI_c_738_n N_CON_M1021_g 0.0196718f $X=3.415 $Y=2.33 $X2=3.845
+ $Y2=3.825
cc_558 N_CI_c_741_n N_CON_M1021_g 9.22089e-19 $X=3.415 $Y=1.96 $X2=3.845
+ $Y2=3.825
cc_559 N_CI_c_743_n N_CON_M1021_g 4.41794e-19 $X=3.415 $Y=2.33 $X2=3.845
+ $Y2=3.825
cc_560 N_CI_c_746_n N_CON_M1021_g 9.30638e-19 $X=4.6 $Y=1.96 $X2=3.845 $Y2=3.825
cc_561 N_CI_c_747_n N_CON_M1021_g 4.44444e-19 $X=3.56 $Y=1.96 $X2=3.845
+ $Y2=3.825
cc_562 N_CI_M1012_g N_CON_c_914_n 0.0207719f $X=3.415 $Y=0.945 $X2=3.845
+ $Y2=1.59
cc_563 N_CI_c_746_n N_CON_c_914_n 0.00158152f $X=4.6 $Y=1.96 $X2=3.845 $Y2=1.59
cc_564 N_CI_M1002_g N_CON_c_916_n 0.00333583f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=0.74
cc_565 N_CI_M1002_g N_CON_c_920_n 0.00386404f $X=1.335 $Y=0.945 $X2=1.665
+ $Y2=2.765
cc_566 N_CI_M1008_g N_CON_c_920_n 0.010554f $X=1.335 $Y=3.825 $X2=1.665
+ $Y2=2.765
cc_567 N_CI_c_737_n N_CON_c_920_n 0.00170665f $X=1.325 $Y=1.96 $X2=1.665
+ $Y2=2.765
cc_568 N_CI_c_740_n N_CON_c_920_n 0.0223962f $X=1.325 $Y=1.96 $X2=1.665
+ $Y2=2.765
cc_569 N_CI_c_744_n N_CON_c_920_n 0.0138278f $X=3.27 $Y=1.96 $X2=1.665 $Y2=2.765
cc_570 N_CI_c_745_n N_CON_c_920_n 0.00183606f $X=1.47 $Y=1.96 $X2=1.665
+ $Y2=2.765
cc_571 N_CI_M1012_g N_CON_c_921_n 0.00137601f $X=3.415 $Y=0.945 $X2=3.97
+ $Y2=1.22
cc_572 N_CI_M1002_g N_CON_c_923_n 0.00402444f $X=1.335 $Y=0.945 $X2=1.665
+ $Y2=1.505
cc_573 N_CI_c_744_n N_CON_c_923_n 7.55969e-19 $X=3.27 $Y=1.96 $X2=1.665
+ $Y2=1.505
cc_574 N_CI_M1008_g N_CON_c_952_n 0.00205937f $X=1.335 $Y=3.825 $X2=1.665
+ $Y2=2.857
cc_575 N_CI_M1012_g N_CON_c_924_n 0.00127353f $X=3.415 $Y=0.945 $X2=3.97
+ $Y2=1.59
cc_576 N_CI_c_746_n N_CON_c_924_n 0.00187655f $X=4.6 $Y=1.96 $X2=3.97 $Y2=1.59
cc_577 N_CI_M1012_g N_CON_c_927_n 0.00167509f $X=3.415 $Y=0.945 $X2=3.825
+ $Y2=1.22
cc_578 N_CI_M1002_g N_CON_c_931_n 0.00317242f $X=1.335 $Y=0.945 $X2=1.695
+ $Y2=1.22
cc_579 N_CI_M1005_g N_CON_c_933_n 0.0107454f $X=4.685 $Y=0.945 $X2=5.995
+ $Y2=1.22
cc_580 N_CI_M1012_g N_A_784_115#_c_1099_n 3.97727e-19 $X=3.415 $Y=0.945
+ $X2=3.845 $Y2=2.77
cc_581 N_CI_M1018_g N_A_784_115#_c_1099_n 0.00502446f $X=3.415 $Y=3.825
+ $X2=3.845 $Y2=2.77
cc_582 N_CI_c_738_n N_A_784_115#_c_1099_n 0.00241496f $X=3.415 $Y=2.33 $X2=3.845
+ $Y2=2.77
cc_583 N_CI_c_741_n N_A_784_115#_c_1099_n 0.0104334f $X=3.415 $Y=1.96 $X2=3.845
+ $Y2=2.77
cc_584 N_CI_c_743_n N_A_784_115#_c_1099_n 0.0114194f $X=3.415 $Y=2.33 $X2=3.845
+ $Y2=2.77
cc_585 N_CI_c_747_n N_A_784_115#_c_1099_n 8.66056e-19 $X=3.56 $Y=1.96 $X2=3.845
+ $Y2=2.77
cc_586 N_CI_M1005_g N_A_784_115#_c_1100_n 8.45664e-19 $X=4.685 $Y=0.945
+ $X2=4.225 $Y2=1.96
cc_587 N_CI_c_742_n N_A_784_115#_c_1100_n 0.00742016f $X=4.745 $Y=1.96 $X2=4.225
+ $Y2=1.96
cc_588 N_CI_c_746_n N_A_784_115#_c_1100_n 0.0202332f $X=4.6 $Y=1.96 $X2=4.225
+ $Y2=1.96
cc_589 N_CI_M1012_g N_A_784_115#_c_1101_n 5.06918e-19 $X=3.415 $Y=0.945 $X2=3.93
+ $Y2=1.96
cc_590 N_CI_c_741_n N_A_784_115#_c_1101_n 0.00810858f $X=3.415 $Y=1.96 $X2=3.93
+ $Y2=1.96
cc_591 N_CI_c_746_n N_A_784_115#_c_1101_n 0.00872498f $X=4.6 $Y=1.96 $X2=3.93
+ $Y2=1.96
cc_592 N_CI_M1018_g N_A_784_115#_c_1114_n 0.00150127f $X=3.415 $Y=3.825 $X2=4.06
+ $Y2=3.16
cc_593 N_CI_M1010_g N_A_784_115#_c_1118_n 0.0193185f $X=4.685 $Y=3.825 $X2=5.33
+ $Y2=3.075
cc_594 N_CI_c_739_n N_A_784_115#_c_1118_n 0.00136691f $X=4.745 $Y=2.14 $X2=5.33
+ $Y2=3.075
cc_595 N_CI_M1005_g N_A_784_115#_c_1102_n 0.0108085f $X=4.685 $Y=0.945 $X2=4.31
+ $Y2=1.875
cc_596 N_CI_c_749_n N_A_784_115#_c_1102_n 0.00139142f $X=4.745 $Y=1.96 $X2=4.31
+ $Y2=1.875
cc_597 N_CI_M1018_g N_A_526_565#_c_1233_n 0.0191262f $X=3.415 $Y=3.825 $X2=3.545
+ $Y2=3.195
cc_598 N_CI_c_738_n N_A_526_565#_c_1233_n 9.07588e-19 $X=3.415 $Y=2.33 $X2=3.545
+ $Y2=3.195
cc_599 N_CI_c_737_n N_A_27_115#_c_1316_n 4.20092e-19 $X=1.325 $Y=1.96 $X2=1.035
+ $Y2=1.175
cc_600 N_CI_M1012_g N_A_526_115#_c_1338_n 0.0138088f $X=3.415 $Y=0.945 $X2=3.545
+ $Y2=1.175
cc_601 N_CI_c_741_n N_A_526_115#_c_1338_n 0.00177004f $X=3.415 $Y=1.96 $X2=3.545
+ $Y2=1.175
cc_602 N_CON_c_921_n N_A_784_115#_M1013_d 0.00133743f $X=3.97 $Y=1.22 $X2=3.92
+ $Y2=0.575
cc_603 N_CON_c_933_n N_A_784_115#_M1013_d 0.00128403f $X=5.995 $Y=1.22 $X2=3.92
+ $Y2=0.575
cc_604 N_CON_c_936_n N_A_784_115#_M1013_d 0.0037089f $X=4.115 $Y=1.22 $X2=3.92
+ $Y2=0.575
cc_605 N_CON_c_922_n N_A_784_115#_M1015_g 0.00198469f $X=6.41 $Y=2.48 $X2=5.585
+ $Y2=0.835
cc_606 N_CON_c_933_n N_A_784_115#_M1015_g 0.0170447f $X=5.995 $Y=1.22 $X2=5.585
+ $Y2=0.835
cc_607 N_CON_c_915_n N_A_784_115#_c_1098_n 0.00451843f $X=6.41 $Y=2.48 $X2=5.585
+ $Y2=2.495
cc_608 N_CON_M1021_g N_A_784_115#_c_1099_n 0.0136798f $X=3.845 $Y=3.825
+ $X2=3.845 $Y2=2.77
cc_609 N_CON_c_914_n N_A_784_115#_c_1100_n 0.00118003f $X=3.845 $Y=1.59
+ $X2=4.225 $Y2=1.96
cc_610 N_CON_c_924_n N_A_784_115#_c_1100_n 0.00732851f $X=3.97 $Y=1.59 $X2=4.225
+ $Y2=1.96
cc_611 N_CON_M1021_g N_A_784_115#_c_1101_n 0.00624765f $X=3.845 $Y=3.825
+ $X2=3.93 $Y2=1.96
cc_612 N_CON_c_914_n N_A_784_115#_c_1101_n 4.82273e-19 $X=3.845 $Y=1.59 $X2=3.93
+ $Y2=1.96
cc_613 N_CON_c_924_n N_A_784_115#_c_1101_n 0.00939629f $X=3.97 $Y=1.59 $X2=3.93
+ $Y2=1.96
cc_614 N_CON_M1021_g N_A_784_115#_c_1114_n 0.0124031f $X=3.845 $Y=3.825 $X2=4.06
+ $Y2=3.16
cc_615 N_CON_c_907_n N_A_784_115#_c_1102_n 0.0010862f $X=3.845 $Y=1.425 $X2=4.31
+ $Y2=1.875
cc_616 N_CON_M1021_g N_A_784_115#_c_1102_n 7.13673e-19 $X=3.845 $Y=3.825
+ $X2=4.31 $Y2=1.875
cc_617 N_CON_c_914_n N_A_784_115#_c_1102_n 8.78503e-19 $X=3.845 $Y=1.59 $X2=4.31
+ $Y2=1.875
cc_618 N_CON_c_921_n N_A_784_115#_c_1102_n 0.0253848f $X=3.97 $Y=1.22 $X2=4.31
+ $Y2=1.875
cc_619 N_CON_c_924_n N_A_784_115#_c_1102_n 0.0115992f $X=3.97 $Y=1.59 $X2=4.31
+ $Y2=1.875
cc_620 N_CON_c_933_n N_A_784_115#_c_1102_n 0.0215575f $X=5.995 $Y=1.22 $X2=4.31
+ $Y2=1.875
cc_621 N_CON_c_936_n N_A_784_115#_c_1102_n 0.00193898f $X=4.115 $Y=1.22 $X2=4.31
+ $Y2=1.875
cc_622 N_CON_c_921_n N_A_784_115#_c_1103_n 0.00382203f $X=3.97 $Y=1.22 $X2=4.06
+ $Y2=0.74
cc_623 N_CON_c_933_n N_A_784_115#_c_1103_n 0.0047062f $X=5.995 $Y=1.22 $X2=4.06
+ $Y2=0.74
cc_624 N_CON_c_936_n N_A_784_115#_c_1103_n 0.00520903f $X=4.115 $Y=1.22 $X2=4.06
+ $Y2=0.74
cc_625 N_CON_M1020_g N_S_c_1244_n 0.00857064f $X=6.535 $Y=0.835 $X2=5.8 $Y2=0.74
cc_626 N_CON_c_922_n N_S_c_1244_n 0.0216008f $X=6.41 $Y=2.48 $X2=5.8 $Y2=0.74
cc_627 N_CON_c_925_n N_S_c_1244_n 0.0121035f $X=6.41 $Y=1.22 $X2=5.8 $Y2=0.74
cc_628 N_CON_c_933_n N_S_c_1244_n 0.021469f $X=5.995 $Y=1.22 $X2=5.8 $Y2=0.74
cc_629 CON N_S_c_1244_n 0.00260317f $X=6.14 $Y=1.22 $X2=5.8 $Y2=0.74
cc_630 N_CON_M1016_g N_S_c_1251_n 0.0214791f $X=6.535 $Y=4.195 $X2=5.8 $Y2=3.105
cc_631 N_CON_M1020_g N_S_c_1249_n 0.00130367f $X=6.535 $Y=0.835 $X2=5.925
+ $Y2=2.905
cc_632 N_CON_M1016_g N_S_c_1249_n 0.00437761f $X=6.535 $Y=4.195 $X2=5.925
+ $Y2=2.905
cc_633 N_CON_c_915_n N_S_c_1249_n 0.00305399f $X=6.41 $Y=2.48 $X2=5.925
+ $Y2=2.905
cc_634 N_CON_c_922_n N_S_c_1249_n 0.0278588f $X=6.41 $Y=2.48 $X2=5.925 $Y2=2.905
cc_635 N_CON_M1020_g N_S_c_1250_n 8.65886e-19 $X=6.535 $Y=0.835 $X2=5.925
+ $Y2=1.96
cc_636 N_CON_c_922_n N_S_c_1250_n 0.00863446f $X=6.41 $Y=2.48 $X2=5.925 $Y2=1.96
cc_637 N_CON_c_933_n N_S_c_1250_n 0.00384217f $X=5.995 $Y=1.22 $X2=5.925
+ $Y2=1.96
cc_638 CON N_S_c_1250_n 5.03075e-19 $X=6.14 $Y=1.22 $X2=5.925 $Y2=1.96
cc_639 N_CON_M1016_g N_S_c_1256_n 0.00293837f $X=6.535 $Y=4.195 $X2=5.925
+ $Y2=2.99
cc_640 N_CON_M1016_g S 0.0029718f $X=6.535 $Y=4.195 $X2=5.8 $Y2=3.105
cc_641 N_CON_M1020_g N_CO_c_1296_n 0.0791316f $X=6.535 $Y=0.835 $X2=6.75
+ $Y2=0.74
cc_642 N_CON_c_922_n N_CO_c_1296_n 0.0950906f $X=6.41 $Y=2.48 $X2=6.75 $Y2=0.74
cc_643 N_CON_c_925_n N_CO_c_1296_n 0.0122992f $X=6.41 $Y=1.22 $X2=6.75 $Y2=0.74
cc_644 CON N_CO_c_1296_n 0.00209642f $X=6.14 $Y=1.22 $X2=6.75 $Y2=0.74
cc_645 N_CON_M1016_g CO 0.00944261f $X=6.535 $Y=4.195 $X2=6.75 $Y2=2.7
cc_646 N_CON_c_915_n CO 0.00612215f $X=6.41 $Y=2.48 $X2=6.75 $Y2=2.7
cc_647 N_CON_c_922_n CO 0.0017516f $X=6.41 $Y=2.48 $X2=6.75 $Y2=2.7
cc_648 N_CON_c_931_n N_A_27_115#_c_1316_n 0.00463163f $X=1.695 $Y=1.22 $X2=1.035
+ $Y2=1.175
cc_649 N_CON_c_916_n N_A_27_115#_c_1318_n 2.23682e-19 $X=1.55 $Y=0.74 $X2=1.12
+ $Y2=0.74
cc_650 N_CON_c_927_n A_368_115# 0.0100396f $X=3.825 $Y=1.22 $X2=1.84 $Y2=0.575
cc_651 N_CON_c_927_n N_A_526_115#_M1019_d 0.00430935f $X=3.825 $Y=1.22 $X2=2.63
+ $Y2=0.575
cc_652 N_CON_c_927_n N_A_526_115#_M1012_d 0.00420198f $X=3.825 $Y=1.22 $X2=3.49
+ $Y2=0.575
cc_653 N_CON_c_921_n N_A_526_115#_c_1338_n 0.00639913f $X=3.97 $Y=1.22 $X2=3.545
+ $Y2=1.175
cc_654 N_CON_c_924_n N_A_526_115#_c_1338_n 0.00170558f $X=3.97 $Y=1.59 $X2=3.545
+ $Y2=1.175
cc_655 N_CON_c_927_n N_A_526_115#_c_1338_n 0.0589959f $X=3.825 $Y=1.22 $X2=3.545
+ $Y2=1.175
cc_656 N_CON_c_936_n N_A_526_115#_c_1338_n 0.00103977f $X=4.115 $Y=1.22
+ $X2=3.545 $Y2=1.175
cc_657 N_CON_c_927_n N_A_526_115#_c_1340_n 0.0167438f $X=3.825 $Y=1.22 $X2=2.855
+ $Y2=1.175
cc_658 N_CON_c_933_n A_870_115# 0.0102308f $X=5.995 $Y=1.22 $X2=4.35 $Y2=0.575
cc_659 N_CON_c_933_n A_952_115# 0.0121403f $X=5.995 $Y=1.22 $X2=4.76 $Y2=0.575
cc_660 N_A_784_115#_c_1118_n A_870_565# 0.0106531f $X=5.33 $Y=3.075 $X2=4.35
+ $Y2=2.825
cc_661 N_A_784_115#_c_1118_n A_952_565# 0.00986639f $X=5.33 $Y=3.075 $X2=4.76
+ $Y2=2.825
cc_662 N_A_784_115#_M1015_g N_S_c_1244_n 0.028079f $X=5.585 $Y=0.835 $X2=5.8
+ $Y2=0.74
cc_663 N_A_784_115#_M1011_g N_S_c_1251_n 0.0271619f $X=5.585 $Y=4.195 $X2=5.8
+ $Y2=3.105
cc_664 N_A_784_115#_c_1118_n N_S_c_1251_n 0.00473093f $X=5.33 $Y=3.075 $X2=5.8
+ $Y2=3.105
cc_665 N_A_784_115#_M1015_g N_S_c_1249_n 0.00949101f $X=5.585 $Y=0.835 $X2=5.925
+ $Y2=2.905
cc_666 N_A_784_115#_M1011_g N_S_c_1249_n 0.00506137f $X=5.585 $Y=4.195 $X2=5.925
+ $Y2=2.905
cc_667 N_A_784_115#_c_1098_n N_S_c_1249_n 0.00346737f $X=5.585 $Y=2.495
+ $X2=5.925 $Y2=2.905
cc_668 N_A_784_115#_c_1121_n N_S_c_1249_n 0.0113616f $X=5.415 $Y=2.99 $X2=5.925
+ $Y2=2.905
cc_669 N_A_784_115#_c_1106_n N_S_c_1249_n 0.0246408f $X=5.415 $Y=2.495 $X2=5.925
+ $Y2=2.905
cc_670 N_A_784_115#_M1015_g N_S_c_1250_n 0.00698062f $X=5.585 $Y=0.835 $X2=5.925
+ $Y2=1.96
cc_671 N_A_784_115#_M1011_g N_S_c_1256_n 0.00358675f $X=5.585 $Y=4.195 $X2=5.925
+ $Y2=2.99
cc_672 N_A_784_115#_c_1118_n N_S_c_1256_n 0.00477774f $X=5.33 $Y=3.075 $X2=5.925
+ $Y2=2.99
cc_673 N_A_784_115#_c_1121_n N_S_c_1256_n 0.00558264f $X=5.415 $Y=2.99 $X2=5.925
+ $Y2=2.99
cc_674 N_A_784_115#_M1011_g S 0.0118598f $X=5.585 $Y=4.195 $X2=5.8 $Y2=3.105
cc_675 N_A_784_115#_c_1098_n S 0.00105962f $X=5.585 $Y=2.495 $X2=5.8 $Y2=3.105
cc_676 N_A_784_115#_c_1118_n S 0.00549343f $X=5.33 $Y=3.075 $X2=5.8 $Y2=3.105
cc_677 N_A_784_115#_c_1106_n S 0.00428732f $X=5.415 $Y=2.495 $X2=5.8 $Y2=3.105
cc_678 N_A_784_115#_c_1103_n N_A_526_115#_c_1341_n 2.24479e-19 $X=4.06 $Y=0.74
+ $X2=3.63 $Y2=0.74
cc_679 N_S_c_1249_n N_CO_c_1296_n 0.0051304f $X=5.925 $Y=2.905 $X2=6.75 $Y2=0.74
cc_680 N_S_c_1256_n N_CO_c_1296_n 0.00509957f $X=5.925 $Y=2.99 $X2=6.75 $Y2=0.74
cc_681 N_S_c_1249_n CO 0.00370359f $X=5.925 $Y=2.905 $X2=6.75 $Y2=2.7
