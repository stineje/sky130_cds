* File: sky130_osu_sc_12T_hs__oai22_l.spice
* Created: Fri Nov 12 15:12:26 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__oai22_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__oai22_l  GND VDD A0 A1 B0 B1 Y
* 
* Y	Y
* B1	B1
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_A0_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1001 N_A_27_115#_M1001_d N_A1_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_115#_M1001_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_A_27_115#_M1007_d N_B1_M1007_g N_Y_M1002_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_A0_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A1_M1006_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.2205 AS=0.1323 PD=1.61 PS=1.47 NRD=5.4569 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 A_282_521# N_B0_M1005_g N_Y_M1006_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.2205 PD=1.47 PS=1.61 NRD=7.8012 NRS=5.4569 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_B1_M1004_g A_282_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=4.87485 P=8.85
pX9_noxref noxref_11 A0 A0 PROBETYPE=1
pX10_noxref noxref_12 A1 A1 PROBETYPE=1
pX11_noxref noxref_13 B0 B0 PROBETYPE=1
pX12_noxref noxref_14 Y Y PROBETYPE=1
pX13_noxref noxref_15 B1 B1 PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__oai22_l.pxi.spice"
*
.ends
*
*
