* File: sky130_osu_sc_18T_ls__xnor2_l.pex.spice
* Created: Thu Oct 29 17:38:56 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%GND 1 2 23 27 29 39 43 49 51
r69 49 51 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r70 43 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r71 37 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.825
r72 30 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r73 25 44 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r74 25 27 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r75 23 37 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r76 23 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r77 23 43 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r78 23 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.17
+ $X2=2.38 $Y2=0.17
r79 23 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r80 23 29 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r81 23 30 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r82 2 39 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.575 $X2=2.44 $Y2=0.825
r83 1 27 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%VDD 1 2 19 23 27 35 41 44 49 50
c40 23 0 1.59951e-19 $X=0.69 $Y=3.455
r41 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=6.49
+ $X2=2.38 $Y2=6.49
r42 44 49 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=2.38 $Y2=6.507
r43 44 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r44 41 53 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r45 41 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r46 35 38 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.44 $Y=3.455
+ $X2=2.44 $Y2=5.835
r47 33 50 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=6.355
+ $X2=2.44 $Y2=6.507
r48 33 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.44 $Y=6.355
+ $X2=2.44 $Y2=5.835
r49 30 32 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r50 28 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r51 28 30 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r52 27 50 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=6.507
+ $X2=2.44 $Y2=6.507
r53 27 32 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=6.507
+ $X2=1.7 $Y2=6.507
r54 23 26 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r55 21 42 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r56 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r57 19 50 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r58 19 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r59 19 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r60 19 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r61 2 38 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.3
+ $Y=3.085 $X2=2.44 $Y2=5.835
r62 2 35 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.3
+ $Y=3.085 $X2=2.44 $Y2=3.455
r63 1 26 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r64 1 23 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%A 3 5 8 9 13 16 18 19 20 24 27 28 31 33
+ 36 37 39 40 45
r114 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.85 $X2=0.845 $Y2=1.85
r115 39 43 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=0.845 $Y=1.725
+ $X2=0.845 $Y2=1.85
r116 39 40 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.725
+ $X2=0.845 $Y2=1.65
r117 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=1.48
+ $X2=2.145 $Y2=1.48
r118 31 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.845 $Y=1.48
+ $X2=0.845 $Y2=1.85
r119 31 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.845 $Y=1.48
+ $X2=0.845 $Y2=1.48
r120 28 33 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.99 $Y=1.48
+ $X2=0.845 $Y2=1.48
r121 27 36 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2 $Y=1.48
+ $X2=2.145 $Y2=1.48
r122 27 28 0.972511 $w=1.7e-07 $l=1.01e-06 $layer=MET1_cond $X=2 $Y=1.48
+ $X2=0.99 $Y2=1.48
r123 25 45 73.8383 $w=2.35e-07 $l=3.6e-07 $layer=POLY_cond $X=2.225 $Y=2.405
+ $X2=1.865 $Y2=2.405
r124 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=2.39 $X2=2.225 $Y2=2.39
r125 22 37 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.145 $Y=2.305
+ $X2=2.145 $Y2=1.48
r126 22 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.305
+ $X2=2.145 $Y2=2.39
r127 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.45 $Y=2.86 $X2=0.45
+ $Y2=3.01
r128 14 45 13.2911 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.865 $Y=2.555
+ $X2=1.865 $Y2=2.405
r129 14 16 1040.91 $w=1.5e-07 $l=2.03e-06 $layer=POLY_cond $X=1.865 $Y=2.555
+ $X2=1.865 $Y2=4.585
r130 13 40 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=1.65
r131 10 18 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=1.725
+ $X2=0.45 $Y2=1.725
r132 9 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=1.725
+ $X2=0.845 $Y2=1.725
r133 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=1.725
+ $X2=0.55 $Y2=1.725
r134 8 20 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=3.01
r135 3 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.45 $Y2=1.725
r136 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.475 $Y2=1.075
r137 1 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=1.8
+ $X2=0.45 $Y2=1.725
r138 1 19 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.425 $Y=1.8
+ $X2=0.425 $Y2=2.86
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%A_27_115# 1 2 9 11 13 16 20 24 28 31 32
+ 34
c78 31 0 1.07013e-19 $X=1.765 $Y=1.85
r79 32 39 15.9603 $w=3.02e-07 $l=1e-07 $layer=POLY_cond $X=1.765 $Y=1.85
+ $X2=1.865 $Y2=1.85
r80 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.85 $X2=1.765 $Y2=1.85
r81 29 31 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.765 $Y=2.305
+ $X2=1.765 $Y2=1.85
r82 28 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=2.39
+ $X2=0.845 $Y2=2.555
r83 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.39 $X2=0.845 $Y2=2.39
r84 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.39
+ $X2=0.26 $Y2=2.39
r85 25 27 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=2.39
+ $X2=0.845 $Y2=2.39
r86 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=2.39
+ $X2=1.765 $Y2=2.305
r87 24 27 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.68 $Y=2.39
+ $X2=0.845 $Y2=2.39
r88 20 22 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r89 18 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.475
+ $X2=0.26 $Y2=2.39
r90 18 20 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.26 $Y=2.475
+ $X2=0.26 $Y2=3.455
r91 14 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.305
+ $X2=0.26 $Y2=2.39
r92 14 16 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.26 $Y=2.305
+ $X2=0.26 $Y2=0.825
r93 11 39 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.685
+ $X2=1.865 $Y2=1.85
r94 11 13 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.865 $Y=1.685
+ $X2=1.865 $Y2=1.075
r95 9 37 1040.91 $w=1.5e-07 $l=2.03e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.555
r96 2 22 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r97 2 20 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r98 1 16 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%A_238_89# 1 2 9 13 15 18 22 26 30
r60 26 28 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.87 $Y=3.455
+ $X2=2.87 $Y2=5.835
r61 24 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.85 $X2=2.87
+ $Y2=2.765
r62 24 26 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.87 $Y=2.85
+ $X2=2.87 $Y2=3.455
r63 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.68 $X2=2.87
+ $Y2=2.765
r64 20 22 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=2.87 $Y=2.68
+ $X2=2.87 $Y2=0.825
r65 18 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.765
+ $X2=1.325 $Y2=2.93
r66 18 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.765
+ $X2=1.325 $Y2=2.6
r67 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.765 $X2=1.325 $Y2=2.765
r68 15 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=2.765
+ $X2=2.87 $Y2=2.765
r69 15 17 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=2.765
+ $X2=1.325 $Y2=2.765
r70 13 33 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.265 $Y=4.585
+ $X2=1.265 $Y2=2.93
r71 9 32 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=1.265 $Y=1.075
+ $X2=1.265 $Y2=2.6
r72 2 28 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.73
+ $Y=3.085 $X2=2.87 $Y2=5.835
r73 2 26 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.73
+ $Y=3.085 $X2=2.87 $Y2=3.455
r74 1 22 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.73
+ $Y=0.575 $X2=2.87 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 17 19 21 27
c56 27 0 1.07013e-19 $X=2.655 $Y=1.832
r57 26 27 21.9891 $w=2.74e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=1.832
+ $X2=2.655 $Y2=1.832
r58 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.85 $X2=2.53 $Y2=1.85
r59 19 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.85
+ $X2=2.53 $Y2=1.85
r60 14 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=3.01
+ $X2=2.655 $Y2=2.935
r61 14 16 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.655 $Y=3.01
+ $X2=2.655 $Y2=4.585
r62 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=2.86
+ $X2=2.655 $Y2=2.935
r63 12 27 16.847 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=2.655 $Y=2.015
+ $X2=2.655 $Y2=1.832
r64 12 13 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=2.655 $Y=2.015
+ $X2=2.655 $Y2=2.86
r65 9 27 16.847 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.832
r66 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.075
r67 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=2.935
+ $X2=2.655 $Y2=2.935
r68 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=2.935 $X2=2.3
+ $Y2=2.935
r69 4 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=3.01
+ $X2=2.3 $Y2=2.935
r70 4 6 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.225 $Y=3.01
+ $X2=2.225 $Y2=4.585
r71 1 26 53.6533 $w=2.74e-07 $l=3.85402e-07 $layer=POLY_cond $X=2.225 $Y=1.65
+ $X2=2.53 $Y2=1.832
r72 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.225 $Y=1.65
+ $X2=2.225 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%Y 1 2 9 11 13 19 23 26 27 30
c56 23 0 1.59951e-19 $X=1.42 $Y=2.135
r57 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=3.33
+ $X2=1.425 $Y2=3.33
r58 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=1.85
+ $X2=1.425 $Y2=1.85
r59 21 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=3.215
+ $X2=1.425 $Y2=3.33
r60 21 23 1.03991 $w=1.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.425 $Y=3.215
+ $X2=1.425 $Y2=2.135
r61 20 26 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.965
+ $X2=1.425 $Y2=1.85
r62 20 23 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.425 $Y=1.965
+ $X2=1.425 $Y2=2.135
r63 19 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.425 $Y=1.415
+ $X2=1.425 $Y2=1.85
r64 18 19 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.537 $Y=1.245
+ $X2=1.537 $Y2=1.415
r65 13 15 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.565 $Y=3.455
+ $X2=1.565 $Y2=5.835
r66 11 31 3.84112 $w=3.85e-07 $l=1.28238e-07 $layer=LI1_cond $X=1.565 $Y=3.445
+ $X2=1.537 $Y2=3.33
r67 11 13 0.338954 $w=3.38e-07 $l=1e-08 $layer=LI1_cond $X=1.565 $Y=3.445
+ $X2=1.565 $Y2=3.455
r68 9 18 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.565 $Y=0.825
+ $X2=1.565 $Y2=1.245
r69 2 15 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.565 $Y2=5.835
r70 2 13 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.565 $Y2=3.455
r71 1 9 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.825
.ends

