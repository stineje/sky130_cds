* File: sky130_osu_sc_15T_ls__addh_l.spice
* Created: Fri Nov 12 14:53:15 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__addh_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__addh_l  GND VDD CON B A S CO
* 
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1007 N_GND_M1007_d N_CON_M1007_g N_S_M1007_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0970254 AS=0.1378 PD=0.891429 PS=1.57 NRD=14.412 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1008 A_208_115# N_B_M1008_g N_GND_M1007_d N_GND_M1007_b NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.138075 PD=0.95 PS=1.26857 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_A_208_565#_M1009_d N_A_M1009_g A_208_115# N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_GND_M1000_d N_A_208_565#_M1000_g N_CO_M1000_s N_GND_M1007_b NSHORT
+ L=0.15 W=0.61 AD=0.10928 AS=0.16165 PD=0.976 PS=1.75 NRD=11.796 NRS=0 M=1
+ R=4.06667 SA=75000.2 SB=75001.5 A=0.0915 P=1.52 MULT=1
MM1010 N_A_570_115#_M1010_d N_A_208_565#_M1010_g N_GND_M1000_d N_GND_M1007_b
+ NSHORT L=0.15 W=0.74 AD=0.1036 AS=0.13257 PD=1.02 PS=1.184 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_CON_M1001_d N_B_M1001_g N_A_570_115#_M1010_d N_GND_M1007_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1003 N_A_570_115#_M1003_d N_A_M1003_g N_CON_M1001_d N_GND_M1007_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VDD_M1004_d N_CON_M1004_g N_S_M1004_s N_VDD_M1004_b PHIGHVT L=0.15
+ W=1.26 AD=0.241371 AS=0.3339 PD=1.80883 PS=3.05 NRD=9.5742 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 N_A_208_565#_M1002_d N_B_M1002_g N_VDD_M1004_d N_VDD_M1004_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.383129 PD=2.28 PS=2.87117 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.5 SB=75000.9 A=0.3 P=4.3 MULT=1
MM1013 N_VDD_M1013_d N_A_M1013_g N_A_208_565#_M1002_d N_VDD_M1004_b PHIGHVT
+ L=0.15 W=2 AD=0.383129 AS=0.28 PD=2.87117 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.9 SB=75000.5 A=0.3 P=4.3 MULT=1
MM1011 N_CO_M1011_d N_A_208_565#_M1011_g N_VDD_M1013_d N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.241371 PD=3.05 PS=1.80883 NRD=0 NRS=9.5742 M=1
+ R=8.4 SA=75001.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1012 N_VDD_M1012_d N_A_208_565#_M1012_g N_CON_M1012_s N_VDD_M1004_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1005 A_668_565# N_B_M1005_g N_VDD_M1012_d N_VDD_M1004_b PHIGHVT L=0.15 W=2
+ AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1006 N_CON_M1006_d N_A_M1006_g A_668_565# N_VDD_M1004_b PHIGHVT L=0.15 W=2
+ AD=0.56 AS=0.21 PD=4.56 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX14_noxref N_GND_M1007_b N_VDD_M1004_b NWDIODE A=12.4785 P=14.36
pX15_noxref noxref_12 S S PROBETYPE=1
pX16_noxref noxref_13 CO CO PROBETYPE=1
pX17_noxref noxref_14 B B PROBETYPE=1
pX18_noxref noxref_15 CON CON PROBETYPE=1
pX19_noxref noxref_16 A A PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__addh_l.pxi.spice"
*
.ends
*
*
