* File: sky130_osu_sc_18T_ms__and2_l.pex.spice
* Created: Thu Oct 29 17:27:44 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__AND2_L%GND 1 12 14 21 26 29
r33 26 29 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r34 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r35 12 19 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r36 12 14 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r37 12 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r38 12 14 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r39 1 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_L%VDD 1 2 13 17 23 32 33 35 38
r25 38 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r26 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r27 32 42 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r28 32 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r29 29 42 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r30 29 31 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r31 23 26 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=4.475
+ $X2=1.12 $Y2=5.835
r32 21 33 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r33 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r34 17 20 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=4.475
+ $X2=0.26 $Y2=5.835
r35 15 31 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r36 15 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r37 13 42 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r38 13 31 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r39 2 26 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=5.835
r40 2 23 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=4.475
r41 1 20 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=5.835
r42 1 17 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_L%A 3 7 12 15 18
r28 16 18 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.765
+ $X2=0.475 $Y2=2.765
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.765 $X2=0.27 $Y2=2.765
r30 11 15 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=2.765
r31 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r32 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=2.765
r33 5 7 1105.01 $w=1.5e-07 $l=2.155e-06 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=5.085
r34 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=2.765
r35 1 3 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_L%B 3 7 12 15 16
r39 16 18 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.59
r40 16 17 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.26
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.425 $X2=0.95 $Y2=2.425
r42 11 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.425
r43 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.96
r44 7 18 1279.35 $w=1.5e-07 $l=2.495e-06 $layer=POLY_cond $X=0.905 $Y=5.085
+ $X2=0.905 $Y2=2.59
r45 3 17 674.287 $w=1.5e-07 $l=1.315e-06 $layer=POLY_cond $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_L%A_27_115# 1 2 9 13 15 17 18 21 23 24 29
+ 35 38 39 40
r68 39 40 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=4.225
+ $X2=0.65 $Y2=4.395
r69 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r70 33 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=0.61 $Y2=1.935
r71 33 35 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=1.43 $Y2=1.935
r72 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=4.475
+ $X2=0.69 $Y2=5.835
r73 29 40 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=4.475 $X2=0.69
+ $Y2=4.395
r74 25 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=2.02 $X2=0.61
+ $Y2=1.935
r75 25 39 143.856 $w=1.68e-07 $l=2.205e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=4.225
r76 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.61 $Y2=1.935
r77 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.345 $Y2=1.935
r78 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.345 $Y2=1.935
r79 19 21 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r80 17 18 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.81
+ $X2=1.352 $Y2=2.96
r81 15 36 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.412 $Y2=1.935
r82 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1 $X2=1.37
+ $Y2=2.81
r83 13 18 1089.63 $w=1.5e-07 $l=2.125e-06 $layer=POLY_cond $X=1.335 $Y=5.085
+ $X2=1.335 $Y2=2.96
r84 7 36 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.412 $Y2=1.935
r85 7 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=0.945
r86 2 31 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=5.835
r87 2 29 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=4.475
r88 1 21 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_L%Y 1 2 10 13 17 18 21
r33 28 30 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=4.475
+ $X2=1.55 $Y2=5.835
r34 18 28 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=4.475
r35 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r36 14 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r37 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r38 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r39 8 10 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r40 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r41 7 10 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r42 2 30 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=4.085 $X2=1.55 $Y2=5.835
r43 2 28 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=4.085 $X2=1.55 $Y2=4.475
r44 1 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

