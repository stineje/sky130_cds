magic
tech sky130A
magscale 1 2
timestamp 1612372607
<< nwell >>
rect -9 529 1456 1119
<< nmoslvt >>
rect 85 115 115 243
rect 171 115 201 243
rect 243 115 273 243
rect 363 115 393 243
rect 435 115 465 243
rect 521 115 551 243
rect 593 115 623 243
rect 713 115 743 243
rect 785 115 815 243
rect 871 115 901 243
rect 1061 115 1091 243
rect 1251 115 1281 225
rect 1337 115 1367 225
<< pmos >>
rect 85 565 115 965
rect 171 565 201 965
rect 243 565 273 965
rect 363 565 393 965
rect 435 565 465 965
rect 521 565 551 965
rect 593 565 623 965
rect 713 565 743 965
rect 785 565 815 965
rect 871 565 901 965
rect 1061 565 1091 965
rect 1251 713 1281 965
rect 1337 713 1367 965
<< ndiff >>
rect 32 215 85 243
rect 32 131 40 215
rect 74 131 85 215
rect 32 115 85 131
rect 115 215 171 243
rect 115 131 126 215
rect 160 131 171 215
rect 115 115 171 131
rect 201 115 243 243
rect 273 215 363 243
rect 273 131 284 215
rect 352 131 363 215
rect 273 115 363 131
rect 393 115 435 243
rect 465 165 521 243
rect 465 131 476 165
rect 510 131 521 165
rect 465 115 521 131
rect 551 115 593 243
rect 623 215 713 243
rect 623 131 634 215
rect 702 131 713 215
rect 623 115 713 131
rect 743 115 785 243
rect 815 215 871 243
rect 815 131 826 215
rect 860 131 871 215
rect 815 115 871 131
rect 901 215 954 243
rect 901 131 912 215
rect 946 131 954 215
rect 901 115 954 131
rect 1008 215 1061 243
rect 1008 131 1016 215
rect 1050 131 1061 215
rect 1008 115 1061 131
rect 1091 215 1144 243
rect 1091 131 1102 215
rect 1136 131 1144 215
rect 1091 115 1144 131
rect 1198 165 1251 225
rect 1198 131 1206 165
rect 1240 131 1251 165
rect 1198 115 1251 131
rect 1281 165 1337 225
rect 1281 131 1292 165
rect 1326 131 1337 165
rect 1281 115 1337 131
rect 1367 165 1420 225
rect 1367 131 1378 165
rect 1412 131 1420 165
rect 1367 115 1420 131
<< pdiff >>
rect 32 949 85 965
rect 32 605 40 949
rect 74 605 85 949
rect 32 565 85 605
rect 115 949 171 965
rect 115 673 126 949
rect 160 673 171 949
rect 115 565 171 673
rect 201 565 243 965
rect 273 949 363 965
rect 273 605 284 949
rect 352 605 363 949
rect 273 565 363 605
rect 393 565 435 965
rect 465 949 521 965
rect 465 673 476 949
rect 510 673 521 949
rect 465 565 521 673
rect 551 565 593 965
rect 623 949 713 965
rect 623 673 634 949
rect 702 673 713 949
rect 623 565 713 673
rect 743 565 785 965
rect 815 949 871 965
rect 815 605 826 949
rect 860 605 871 949
rect 815 565 871 605
rect 901 949 954 965
rect 901 605 912 949
rect 946 605 954 949
rect 901 565 954 605
rect 1008 949 1061 965
rect 1008 673 1016 949
rect 1050 673 1061 949
rect 1008 565 1061 673
rect 1091 949 1144 965
rect 1091 605 1102 949
rect 1136 605 1144 949
rect 1198 949 1251 965
rect 1198 877 1206 949
rect 1240 877 1251 949
rect 1198 713 1251 877
rect 1281 949 1337 965
rect 1281 877 1292 949
rect 1326 877 1337 949
rect 1281 713 1337 877
rect 1367 949 1420 965
rect 1367 877 1378 949
rect 1412 877 1420 949
rect 1367 713 1420 877
rect 1091 565 1144 605
<< ndiffc >>
rect 40 131 74 215
rect 126 131 160 215
rect 284 131 352 215
rect 476 131 510 165
rect 634 131 702 215
rect 826 131 860 215
rect 912 131 946 215
rect 1016 131 1050 215
rect 1102 131 1136 215
rect 1206 131 1240 165
rect 1292 131 1326 165
rect 1378 131 1412 165
<< pdiffc >>
rect 40 605 74 949
rect 126 673 160 949
rect 284 605 352 949
rect 476 673 510 949
rect 634 673 702 949
rect 826 605 860 949
rect 912 605 946 949
rect 1016 673 1050 949
rect 1102 605 1136 949
rect 1206 877 1240 949
rect 1292 877 1326 949
rect 1378 877 1412 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
rect 979 27 1003 61
rect 1037 27 1061 61
rect 1115 27 1139 61
rect 1173 27 1197 61
rect 1251 27 1275 61
rect 1309 27 1333 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
rect 571 1049 595 1083
rect 629 1049 653 1083
rect 707 1049 731 1083
rect 765 1049 789 1083
rect 843 1049 867 1083
rect 901 1049 925 1083
rect 979 1049 1003 1083
rect 1037 1049 1061 1083
rect 1115 1049 1139 1083
rect 1173 1049 1197 1083
rect 1251 1049 1275 1083
rect 1309 1049 1333 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
rect 1003 27 1037 61
rect 1139 27 1173 61
rect 1275 27 1309 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
rect 595 1049 629 1083
rect 731 1049 765 1083
rect 867 1049 901 1083
rect 1003 1049 1037 1083
rect 1139 1049 1173 1083
rect 1275 1049 1309 1083
<< poly >>
rect 85 965 115 991
rect 171 965 201 991
rect 243 965 273 991
rect 363 965 393 991
rect 435 965 465 991
rect 521 965 551 991
rect 593 965 623 991
rect 713 965 743 991
rect 785 965 815 991
rect 871 965 901 991
rect 1061 965 1091 991
rect 1251 965 1281 991
rect 1337 965 1367 991
rect 85 534 115 565
rect 75 518 129 534
rect 75 484 85 518
rect 119 484 129 518
rect 75 468 129 484
rect 75 322 105 468
rect 171 425 201 565
rect 243 534 273 565
rect 243 518 297 534
rect 243 484 253 518
rect 287 484 297 518
rect 243 468 297 484
rect 171 409 225 425
rect 363 423 393 565
rect 435 528 465 565
rect 521 528 551 565
rect 435 518 551 528
rect 435 484 467 518
rect 501 484 551 518
rect 435 474 551 484
rect 593 423 623 565
rect 713 534 743 565
rect 689 518 743 534
rect 689 484 699 518
rect 733 484 743 518
rect 689 468 743 484
rect 171 375 181 409
rect 215 375 225 409
rect 171 359 225 375
rect 267 393 719 423
rect 75 292 115 322
rect 85 243 115 292
rect 171 243 201 359
rect 267 315 297 393
rect 689 351 719 393
rect 785 419 815 565
rect 871 534 901 565
rect 871 518 942 534
rect 871 504 898 518
rect 882 484 898 504
rect 932 484 942 518
rect 882 468 942 484
rect 785 403 839 419
rect 785 369 795 403
rect 829 369 839 403
rect 785 353 839 369
rect 243 285 297 315
rect 339 335 393 351
rect 339 301 349 335
rect 383 301 393 335
rect 339 285 393 301
rect 243 243 273 285
rect 363 243 393 285
rect 435 335 551 345
rect 435 301 467 335
rect 501 301 551 335
rect 435 291 551 301
rect 435 243 465 291
rect 521 243 551 291
rect 593 335 647 351
rect 593 301 603 335
rect 637 301 647 335
rect 593 285 647 301
rect 689 335 743 351
rect 689 301 699 335
rect 733 301 743 335
rect 689 285 743 301
rect 593 243 623 285
rect 713 243 743 285
rect 785 243 815 353
rect 882 315 912 468
rect 1061 351 1091 565
rect 1251 549 1281 713
rect 1241 519 1281 549
rect 1241 419 1271 519
rect 1337 460 1367 713
rect 1216 403 1271 419
rect 1216 369 1226 403
rect 1260 369 1271 403
rect 1313 444 1367 460
rect 1313 410 1323 444
rect 1357 410 1367 444
rect 1313 394 1367 410
rect 1216 353 1271 369
rect 871 285 912 315
rect 1008 335 1091 351
rect 1008 301 1018 335
rect 1052 301 1091 335
rect 1008 285 1091 301
rect 871 243 901 285
rect 1061 243 1091 285
rect 1241 308 1271 353
rect 1241 278 1281 308
rect 1251 225 1281 278
rect 1337 225 1367 394
rect 85 89 115 115
rect 171 89 201 115
rect 243 89 273 115
rect 363 89 393 115
rect 435 89 465 115
rect 521 89 551 115
rect 593 89 623 115
rect 713 89 743 115
rect 785 89 815 115
rect 871 89 901 115
rect 1061 89 1091 115
rect 1251 89 1281 115
rect 1337 89 1367 115
<< polycont >>
rect 85 484 119 518
rect 253 484 287 518
rect 467 484 501 518
rect 699 484 733 518
rect 181 375 215 409
rect 898 484 932 518
rect 795 369 829 403
rect 349 301 383 335
rect 467 301 501 335
rect 603 301 637 335
rect 699 301 733 335
rect 1226 369 1260 403
rect 1323 410 1357 444
rect 1018 301 1052 335
<< locali >>
rect 0 1089 1452 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 595 1089
rect 629 1049 731 1089
rect 765 1049 867 1089
rect 901 1049 1003 1089
rect 1037 1049 1139 1089
rect 1173 1049 1275 1089
rect 1309 1049 1452 1089
rect 40 949 74 965
rect 17 605 40 617
rect 126 949 160 1049
rect 126 657 160 673
rect 284 949 352 965
rect 17 583 74 605
rect 476 949 510 1049
rect 476 657 510 673
rect 634 949 702 965
rect 352 605 355 623
rect 284 602 355 605
rect 634 602 702 673
rect 17 335 51 583
rect 108 568 355 602
rect 535 568 702 602
rect 826 949 860 1049
rect 826 589 860 605
rect 912 949 946 965
rect 1016 949 1050 1049
rect 1016 657 1050 673
rect 1102 949 1136 965
rect 912 602 946 605
rect 912 568 1000 602
rect 108 534 142 568
rect 85 518 142 534
rect 119 484 142 518
rect 85 468 142 484
rect 17 301 40 335
rect 17 280 74 301
rect 108 318 142 468
rect 253 518 287 534
rect 253 483 287 484
rect 467 518 501 534
rect 287 449 383 483
rect 181 409 215 425
rect 181 359 215 375
rect 349 335 383 449
rect 467 335 501 484
rect 108 284 315 318
rect 349 285 383 301
rect 467 285 501 301
rect 535 335 569 568
rect 699 518 733 534
rect 699 483 733 484
rect 40 215 74 280
rect 281 231 315 284
rect 535 251 569 301
rect 603 449 699 483
rect 898 518 932 534
rect 898 483 932 484
rect 603 335 637 449
rect 966 403 1000 568
rect 779 369 795 403
rect 829 369 845 403
rect 912 369 1000 403
rect 1102 403 1136 605
rect 1206 949 1240 965
rect 1206 557 1240 877
rect 1292 949 1326 1049
rect 1292 861 1326 877
rect 1378 949 1412 965
rect 1378 631 1412 877
rect 1411 614 1412 631
rect 1411 597 1435 614
rect 1378 580 1435 597
rect 1206 518 1240 523
rect 1206 484 1357 518
rect 1323 444 1357 484
rect 1102 369 1226 403
rect 1260 369 1276 403
rect 912 335 946 369
rect 683 301 699 335
rect 733 301 946 335
rect 1002 301 1018 335
rect 1052 301 1068 335
rect 603 285 637 301
rect 40 115 74 131
rect 126 215 160 231
rect 281 215 352 231
rect 535 217 702 251
rect 281 197 284 215
rect 126 61 160 131
rect 634 215 702 217
rect 284 115 352 131
rect 476 165 510 181
rect 476 61 510 131
rect 634 115 702 131
rect 826 215 860 231
rect 826 61 860 131
rect 912 215 946 301
rect 912 115 946 131
rect 1016 215 1050 231
rect 1016 61 1050 131
rect 1102 215 1136 369
rect 1323 335 1357 410
rect 1102 115 1136 131
rect 1206 301 1357 335
rect 1206 165 1240 301
rect 1401 268 1435 580
rect 1378 234 1435 268
rect 1206 115 1240 131
rect 1292 165 1326 181
rect 1292 61 1326 131
rect 1378 165 1412 234
rect 1378 115 1412 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1003 61
rect 1037 21 1139 61
rect 1173 21 1275 61
rect 1309 21 1452 61
rect 0 0 1452 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 595 1083 629 1089
rect 595 1055 629 1083
rect 731 1083 765 1089
rect 731 1055 765 1083
rect 867 1083 901 1089
rect 867 1055 901 1083
rect 1003 1083 1037 1089
rect 1003 1055 1037 1083
rect 1139 1083 1173 1089
rect 1139 1055 1173 1083
rect 1275 1083 1309 1089
rect 1275 1055 1309 1083
rect 40 301 74 335
rect 253 449 287 483
rect 181 375 215 409
rect 449 301 467 335
rect 467 301 483 335
rect 535 301 569 335
rect 699 449 733 483
rect 898 449 932 483
rect 795 369 829 403
rect 1377 597 1411 631
rect 1206 523 1240 557
rect 1226 369 1260 403
rect 1018 301 1052 335
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
rect 1003 27 1037 55
rect 1003 21 1037 27
rect 1139 27 1173 55
rect 1139 21 1173 27
rect 1275 27 1309 55
rect 1275 21 1309 27
<< metal1 >>
rect 0 1089 1452 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 595 1089
rect 629 1055 731 1089
rect 765 1055 867 1089
rect 901 1055 1003 1089
rect 1037 1055 1139 1089
rect 1173 1055 1275 1089
rect 1309 1055 1452 1089
rect 0 1049 1452 1055
rect 1365 631 1423 637
rect 1343 597 1377 631
rect 1411 597 1423 631
rect 1365 591 1423 597
rect 1194 557 1252 563
rect 1172 523 1206 557
rect 1240 523 1252 557
rect 1194 517 1252 523
rect 241 483 299 489
rect 687 483 745 489
rect 886 483 944 489
rect 241 449 253 483
rect 287 449 699 483
rect 733 449 898 483
rect 932 449 944 483
rect 241 443 299 449
rect 687 443 745 449
rect 886 443 944 449
rect 169 409 227 415
rect 169 375 181 409
rect 215 375 249 409
rect 783 403 841 409
rect 1214 403 1272 409
rect 169 369 227 375
rect 783 369 795 403
rect 829 369 1226 403
rect 1260 369 1272 403
rect 783 363 841 369
rect 1214 363 1272 369
rect 28 335 86 341
rect 437 335 495 341
rect 28 301 40 335
rect 74 301 449 335
rect 483 301 495 335
rect 28 295 86 301
rect 437 295 495 301
rect 523 335 581 341
rect 1006 335 1064 341
rect 523 301 535 335
rect 569 301 1018 335
rect 1052 301 1064 335
rect 523 295 581 301
rect 1006 295 1064 301
rect 0 55 1452 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1003 55
rect 1037 21 1139 55
rect 1173 21 1275 55
rect 1309 21 1452 55
rect 0 0 1452 21
<< labels >>
rlabel viali 198 392 198 392 1 D
port 1 n
rlabel viali 1394 614 1394 614 1 Q
port 2 n
rlabel viali 1224 540 1224 540 1 QN
port 3 n
rlabel viali 915 466 915 466 1 CK
port 4 n
rlabel viali 68 49 68 49 1 gnd
rlabel viali 68 1063 68 1063 1 vdd
<< end >>
