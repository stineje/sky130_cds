* File: sky130_osu_sc_15T_ls__buf_2.pex.spice
* Created: Fri Nov 12 14:54:50 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__BUF_2%GND 1 2 21 23 30 32 40 44 47
r34 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r35 38 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.865
r36 33 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r37 32 38 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.305
r38 28 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r39 28 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.865
r40 23 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r41 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r42 21 32 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r43 21 33 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r44 21 23 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r45 2 40 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.865
r46 1 30 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_2%VDD 1 2 17 19 25 29 36 42 45
r26 42 45 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r27 36 39 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.205
+ $X2=1.55 $Y2=4.565
r28 34 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=5.245
+ $X2=1.55 $Y2=4.565
r29 32 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r30 30 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r31 30 32 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r32 29 34 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.465 $Y=5.397
+ $X2=1.55 $Y2=5.245
r33 29 32 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=5.397
+ $X2=1.02 $Y2=5.397
r34 25 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=3.885
+ $X2=0.69 $Y2=4.565
r35 23 40 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r36 23 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r37 19 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r38 19 21 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r39 17 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r40 17 21 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r41 2 39 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.565
r42 2 36 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.205
r43 1 28 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r44 1 25 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_2%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.07
+ $X2=0.635 $Y2=3.07
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2.22
+ $X2=0.635 $Y2=3.07
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.22 $X2=0.635 $Y2=2.22
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.22
+ $X2=0.585 $Y2=2.385
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.22
+ $X2=0.585 $Y2=2.055
r45 7 12 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.385
r46 3 11 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_2%A_27_115# 1 3 11 13 15 17 20 22 24 28 33
+ 37 41 45 47 50
r69 46 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.675
+ $X2=0.26 $Y2=1.675
r70 45 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.675
+ $X2=0.965 $Y2=1.675
r71 45 46 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.675
+ $X2=0.345 $Y2=1.675
r72 41 43 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r73 39 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.76 $X2=0.26
+ $Y2=1.675
r74 39 41 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=0.26 $Y=1.76
+ $X2=0.26 $Y2=3.205
r75 35 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.59 $X2=0.26
+ $Y2=1.675
r76 35 37 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.865
r77 32 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.675 $X2=0.965 $Y2=1.675
r78 32 33 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=1.18 $Y2=1.675
r79 30 32 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.965 $Y2=1.675
r80 27 28 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.675
+ $X2=1.335 $Y2=2.675
r81 25 27 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.675
+ $X2=1.18 $Y2=2.675
r82 22 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.75
+ $X2=1.335 $Y2=2.675
r83 22 24 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.335 $Y=2.75
+ $X2=1.335 $Y2=3.825
r84 18 33 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.18 $Y2=1.675
r85 18 20 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.945
r86 17 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.6 $X2=1.18
+ $Y2=2.675
r87 16 33 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.84
+ $X2=1.18 $Y2=1.675
r88 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.84
+ $X2=1.18 $Y2=2.6
r89 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=2.675
r90 13 15 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=3.825
r91 9 30 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.905 $Y2=1.675
r92 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.905 $Y2=0.945
r93 3 43 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r94 3 41 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r95 1 37 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_2%Y 1 3 10 16 26 29 32
r39 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.585
+ $X2=1.12 $Y2=2.7
r40 24 26 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.585
+ $X2=1.12 $Y2=2.01
r41 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=1.22
r42 23 26 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=2.01
r43 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=3.205
+ $X2=1.12 $Y2=4.565
r44 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.7 $X2=1.12
+ $Y2=2.7
r45 16 19 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.12 $Y=2.7
+ $X2=1.12 $Y2=3.205
r46 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.22
+ $X2=1.12 $Y2=1.22
r47 10 13 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.12 $Y=0.865
+ $X2=1.12 $Y2=1.22
r48 3 21 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r49 3 19 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.205
r50 1 10 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
.ends

