* File: sky130_osu_sc_15T_hs__inv_l.pxi.spice
* Created: Fri Nov 12 14:31:24 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__INV_L%GND N_GND_M1001_s N_GND_M1001_b N_GND_c_2_p
+ N_GND_c_3_p GND PM_SKY130_OSU_SC_15T_HS__INV_L%GND
x_PM_SKY130_OSU_SC_15T_HS__INV_L%VDD N_VDD_M1000_s N_VDD_M1000_b N_VDD_c_16_p
+ N_VDD_c_17_p VDD PM_SKY130_OSU_SC_15T_HS__INV_L%VDD
x_PM_SKY130_OSU_SC_15T_HS__INV_L%A N_A_M1001_g N_A_M1000_g N_A_c_29_n N_A_c_30_n
+ N_A_c_31_n N_A_c_32_n A PM_SKY130_OSU_SC_15T_HS__INV_L%A
x_PM_SKY130_OSU_SC_15T_HS__INV_L%Y N_Y_M1001_d N_Y_M1000_d N_Y_c_59_n N_Y_c_61_n
+ Y N_Y_c_63_n N_Y_c_64_n PM_SKY130_OSU_SC_15T_HS__INV_L%Y
cc_1 N_GND_M1001_b N_A_M1001_g 0.0934528f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_A_M1001_g 0.00502587f $X=0.26 $Y=0.74 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_A_M1001_g 0.00468827f $X=0.34 $Y=0.19 $X2=0.475 $Y2=0.85
cc_4 N_GND_M1001_b N_A_M1000_g 0.0337175f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.195
cc_5 N_GND_M1001_b N_A_c_29_n 0.0393936f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.045
cc_6 N_GND_M1001_b N_A_c_30_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.07
cc_7 N_GND_M1001_b N_A_c_31_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.045
cc_8 N_GND_M1001_b N_A_c_32_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.045
cc_9 N_GND_M1001_b N_Y_c_59_n 0.0166829f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.74
cc_10 N_GND_c_3_p N_Y_c_59_n 0.00476261f $X=0.34 $Y=0.19 $X2=0.69 $Y2=0.74
cc_11 N_GND_M1001_b N_Y_c_61_n 0.00237997f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.7
cc_12 N_GND_M1001_b Y 0.0587019f $X=-0.045 $Y=0 $X2=0.755 $Y2=1.945
cc_13 N_GND_M1001_b N_Y_c_63_n 0.0126319f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.22
cc_14 N_GND_M1001_b N_Y_c_64_n 0.00507896f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.7
cc_15 N_VDD_M1000_b N_A_M1000_g 0.0871966f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=4.195
cc_16 N_VDD_c_16_p N_A_M1000_g 0.00751602f $X=0.26 $Y=4.565 $X2=0.475 $Y2=4.195
cc_17 N_VDD_c_17_p N_A_M1000_g 0.00496961f $X=0.34 $Y=5.36 $X2=0.475 $Y2=4.195
cc_18 VDD N_A_M1000_g 0.00429146f $X=0.34 $Y=5.31 $X2=0.475 $Y2=4.195
cc_19 N_VDD_M1000_b N_A_c_30_n 0.0153337f $X=-0.045 $Y=2.645 $X2=0.32 $Y2=3.07
cc_20 N_VDD_M1000_b A 0.0221642f $X=-0.045 $Y=2.645 $X2=0.32 $Y2=3.07
cc_21 N_VDD_M1000_b N_Y_c_61_n 0.0415234f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.7
cc_22 N_VDD_c_17_p N_Y_c_61_n 0.00477009f $X=0.34 $Y=5.36 $X2=0.69 $Y2=2.7
cc_23 VDD N_Y_c_61_n 0.00435496f $X=0.34 $Y=5.31 $X2=0.69 $Y2=2.7
cc_24 N_VDD_M1000_b N_Y_c_64_n 0.00914195f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.7
cc_25 N_A_M1001_g N_Y_c_59_n 0.00971844f $X=0.475 $Y=0.85 $X2=0.69 $Y2=0.74
cc_26 N_A_c_29_n N_Y_c_59_n 6.24081e-19 $X=0.535 $Y=2.045 $X2=0.69 $Y2=0.74
cc_27 N_A_c_32_n N_Y_c_59_n 0.00124107f $X=0.535 $Y=2.045 $X2=0.69 $Y2=0.74
cc_28 N_A_M1000_g N_Y_c_61_n 0.0434722f $X=0.475 $Y=4.195 $X2=0.69 $Y2=2.7
cc_29 N_A_c_29_n N_Y_c_61_n 8.13098e-19 $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.7
cc_30 N_A_c_30_n N_Y_c_61_n 0.0305887f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.7
cc_31 N_A_c_32_n N_Y_c_61_n 0.00202105f $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.7
cc_32 A N_Y_c_61_n 0.0149533f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.7
cc_33 N_A_M1001_g Y 0.0127139f $X=0.475 $Y=0.85 $X2=0.755 $Y2=1.945
cc_34 N_A_M1000_g Y 0.00874077f $X=0.475 $Y=4.195 $X2=0.755 $Y2=1.945
cc_35 N_A_c_29_n Y 0.00719822f $X=0.535 $Y=2.045 $X2=0.755 $Y2=1.945
cc_36 N_A_c_30_n Y 0.0183799f $X=0.32 $Y=3.07 $X2=0.755 $Y2=1.945
cc_37 N_A_c_32_n Y 0.0178517f $X=0.535 $Y=2.045 $X2=0.755 $Y2=1.945
cc_38 N_A_M1001_g N_Y_c_63_n 0.0119993f $X=0.475 $Y=0.85 $X2=0.69 $Y2=1.22
cc_39 N_A_c_29_n N_Y_c_63_n 0.0011424f $X=0.535 $Y=2.045 $X2=0.69 $Y2=1.22
cc_40 N_A_M1000_g N_Y_c_64_n 0.00478745f $X=0.475 $Y=4.195 $X2=0.69 $Y2=2.7
cc_41 N_A_c_29_n N_Y_c_64_n 0.00126139f $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.7
cc_42 N_A_c_30_n N_Y_c_64_n 0.00640429f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.7
cc_43 N_A_c_32_n N_Y_c_64_n 0.00194461f $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.7
cc_44 A N_Y_c_64_n 0.00827053f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.7
