* File: sky130_osu_sc_18T_ms__or2_8.pex.spice
* Created: Thu Oct 29 17:31:22 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__OR2_8%GND 1 2 3 4 5 6 47 51 53 60 62 69 71 78
+ 80 87 91 100 105 107
r135 105 107 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r136 89 100 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.475 $Y2=0.152
r137 89 91 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.56 $Y2=0.825
r138 85 87 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.825
r139 81 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r140 76 95 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r141 76 78 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.825
r142 72 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r143 71 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r144 67 94 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r145 67 69 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r146 63 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r147 62 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r148 58 93 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r149 58 60 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r150 53 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r151 49 51 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r152 47 49 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r153 47 54 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r154 47 100 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.475 $Y2=0.152
r155 47 96 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=3.785 $Y2=0.152
r156 47 107 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.17
+ $X2=4.42 $Y2=0.17
r157 47 105 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r158 47 85 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.7 $Y2=0.305
r159 47 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.615 $Y2=0.152
r160 47 96 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.785 $Y2=0.152
r161 47 80 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r162 47 81 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r163 47 71 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r164 47 72 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r165 47 62 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r166 47 63 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r167 47 53 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r168 47 54 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r169 6 91 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.575 $X2=4.56 $Y2=0.825
r170 5 87 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.825
r171 4 78 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r172 3 69 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r173 2 60 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r174 1 51 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__OR2_8%VDD 1 2 3 4 5 37 41 45 51 55 61 65 71 77
+ 81 88 90 95
r81 99 102 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r82 95 104 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=6.49
+ $X2=4.42 $Y2=6.49
r83 90 95 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=4.42 $Y2=6.507
r84 90 99 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r85 88 104 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.475 $Y=6.507
+ $X2=4.42 $Y2=6.507
r86 85 104 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=6.507
+ $X2=4.42 $Y2=6.507
r87 85 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=6.507
+ $X2=3.7 $Y2=6.507
r88 81 102 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r89 81 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r90 77 80 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.56 $Y=3.455
+ $X2=4.56 $Y2=5.835
r91 75 88 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.56 $Y=6.355
+ $X2=4.475 $Y2=6.507
r92 75 80 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.56 $Y=6.355
+ $X2=4.56 $Y2=5.835
r93 71 74 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.7 $Y=3.455
+ $X2=3.7 $Y2=5.835
r94 69 87 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.7 $Y=6.355 $X2=3.7
+ $Y2=6.507
r95 69 74 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.7 $Y=6.355 $X2=3.7
+ $Y2=5.835
r96 66 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=6.507
+ $X2=2.84 $Y2=6.507
r97 66 68 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=6.507
+ $X2=3.06 $Y2=6.507
r98 65 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=6.507
+ $X2=3.7 $Y2=6.507
r99 65 68 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=6.507
+ $X2=3.06 $Y2=6.507
r100 61 64 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r101 59 84 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.84 $Y2=6.507
r102 59 64 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.84 $Y2=5.835
r103 56 83 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=1.98 $Y2=6.507
r104 56 58 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=2.38 $Y2=6.507
r105 55 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.84 $Y2=6.507
r106 55 58 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.38 $Y2=6.507
r107 51 54 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r108 49 83 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=6.507
r109 49 54 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r110 46 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r111 46 48 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r112 45 83 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.98 $Y2=6.507
r113 45 48 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r114 41 44 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=5.835
r115 39 82 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r116 39 44 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r117 37 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r118 37 102 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r119 37 99 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r120 37 87 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r121 37 68 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r122 37 58 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r123 37 48 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r124 5 80 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.42
+ $Y=3.085 $X2=4.56 $Y2=5.835
r125 5 77 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.42
+ $Y=3.085 $X2=4.56 $Y2=3.455
r126 4 74 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=5.835
r127 4 71 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=3.455
r128 3 64 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r129 3 61 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r130 2 54 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r131 2 51 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r132 1 44 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r133 1 41 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__OR2_8%B 3 7 10 15 18
r28 16 18 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.675
+ $X2=0.475 $Y2=2.675
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.675 $X2=0.27 $Y2=2.675
r30 12 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.96
+ $X2=0.27 $Y2=2.675
r31 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.96
+ $X2=0.27 $Y2=2.96
r32 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.84
+ $X2=0.475 $Y2=2.675
r33 5 7 894.777 $w=1.5e-07 $l=1.745e-06 $layer=POLY_cond $X=0.475 $Y=2.84
+ $X2=0.475 $Y2=4.585
r34 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.51
+ $X2=0.475 $Y2=2.675
r35 1 3 735.819 $w=1.5e-07 $l=1.435e-06 $layer=POLY_cond $X=0.475 $Y=2.51
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__OR2_8%A 3 7 10 15 16
c44 7 0 1.37149e-19 $X=0.905 $Y=4.585
r45 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=2.55
r46 16 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=2.22
r47 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.385 $X2=0.95 $Y2=2.385
r48 12 15 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.95 $Y2=2.385
r49 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=3.33
+ $X2=0.95 $Y2=3.33
r50 7 18 1043.48 $w=1.5e-07 $l=2.035e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.55
r51 3 17 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.22
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__OR2_8%A_27_617# 1 2 9 11 13 15 16 20 22 24 25
+ 26 27 31 33 35 36 38 42 44 46 47 49 53 56 57 59 60 62 66 68 70 71 73 77 79 81
+ 82 84 88 90 92 93 94 95 96 97 98 99 100 101 102 103 104 107 111 112 114 117
+ 121 124
c243 66 0 1.33323e-19 $X=3.485 $Y=1.075
c244 53 0 1.33323e-19 $X=3.055 $Y=1.075
c245 42 0 1.33323e-19 $X=2.625 $Y=1.075
c246 31 0 1.33323e-19 $X=2.195 $Y=1.075
c247 20 0 1.33323e-19 $X=1.765 $Y=1.075
r248 125 126 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.935
+ $X2=1.37 $Y2=1.935
r249 122 126 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.43 $Y=1.935
+ $X2=1.37 $Y2=1.935
r250 121 122 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r251 119 124 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.935
+ $X2=0.65 $Y2=1.935
r252 119 121 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.935
+ $X2=1.43 $Y2=1.935
r253 115 124 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.65 $Y2=1.935
r254 115 117 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=0.825
r255 113 124 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.65 $Y2=1.935
r256 113 114 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r257 111 114 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.63
+ $X2=0.61 $Y2=3.545
r258 111 112 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.63
+ $X2=0.345 $Y2=3.63
r259 107 109 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.26 $Y=3.795
+ $X2=0.26 $Y2=5.835
r260 105 112 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.715
+ $X2=0.345 $Y2=3.63
r261 105 107 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=3.715
+ $X2=0.26 $Y2=3.795
r262 90 92 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=4.345 $Y=2.96
+ $X2=4.345 $Y2=4.585
r263 86 88 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.345 $Y=1.77
+ $X2=4.345 $Y2=1.075
r264 85 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=2.885
+ $X2=3.915 $Y2=2.885
r265 84 90 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=2.885
+ $X2=4.345 $Y2=2.96
r266 84 85 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=2.885
+ $X2=3.99 $Y2=2.885
r267 83 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.845
+ $X2=3.915 $Y2=1.845
r268 82 86 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=1.845
+ $X2=4.345 $Y2=1.77
r269 82 83 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.845
+ $X2=3.99 $Y2=1.845
r270 79 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=2.96
+ $X2=3.915 $Y2=2.885
r271 79 81 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=3.915 $Y=2.96
+ $X2=3.915 $Y2=4.585
r272 75 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=1.77
+ $X2=3.915 $Y2=1.845
r273 75 77 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.915 $Y=1.77
+ $X2=3.915 $Y2=1.075
r274 74 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.885
+ $X2=3.485 $Y2=2.885
r275 73 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.885
+ $X2=3.915 $Y2=2.885
r276 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.885
+ $X2=3.56 $Y2=2.885
r277 72 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.845
+ $X2=3.485 $Y2=1.845
r278 71 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.845
+ $X2=3.915 $Y2=1.845
r279 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.845
+ $X2=3.56 $Y2=1.845
r280 68 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.96
+ $X2=3.485 $Y2=2.885
r281 68 70 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=3.485 $Y=2.96
+ $X2=3.485 $Y2=4.585
r282 64 101 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.845
r283 64 66 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.075
r284 63 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.885
+ $X2=3.055 $Y2=2.885
r285 62 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.885
+ $X2=3.485 $Y2=2.885
r286 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.885
+ $X2=3.13 $Y2=2.885
r287 61 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.845
+ $X2=3.055 $Y2=1.845
r288 60 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.485 $Y2=1.845
r289 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.13 $Y2=1.845
r290 57 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.96
+ $X2=3.055 $Y2=2.885
r291 57 59 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=3.055 $Y=2.96
+ $X2=3.055 $Y2=4.585
r292 56 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.81
+ $X2=3.055 $Y2=2.885
r293 55 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.92
+ $X2=3.055 $Y2=1.845
r294 55 56 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.055 $Y=1.92
+ $X2=3.055 $Y2=2.81
r295 51 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.845
r296 51 53 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.075
r297 50 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.885
+ $X2=2.625 $Y2=2.885
r298 49 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.885
+ $X2=3.055 $Y2=2.885
r299 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.885
+ $X2=2.7 $Y2=2.885
r300 48 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.845
+ $X2=2.625 $Y2=1.845
r301 47 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=3.055 $Y2=1.845
r302 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=2.7 $Y2=1.845
r303 44 98 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.96
+ $X2=2.625 $Y2=2.885
r304 44 46 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.625 $Y=2.96
+ $X2=2.625 $Y2=4.585
r305 40 97 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.845
r306 40 42 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.075
r307 39 96 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.885
+ $X2=2.195 $Y2=2.885
r308 38 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.625 $Y2=2.885
r309 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.27 $Y2=2.885
r310 37 95 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.195 $Y2=1.845
r311 36 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.625 $Y2=1.845
r312 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.27 $Y2=1.845
r313 33 96 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=2.885
r314 33 35 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=4.585
r315 29 95 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.845
r316 29 31 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r317 28 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.885
+ $X2=1.765 $Y2=2.885
r318 27 96 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=2.195 $Y2=2.885
r319 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=1.84 $Y2=2.885
r320 25 95 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.845
r321 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r322 22 94 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=2.885
r323 22 24 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r324 18 26 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.84 $Y2=1.845
r325 18 122 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.43 $Y2=1.935
r326 18 20 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r327 17 93 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.885
+ $X2=1.352 $Y2=2.885
r328 16 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.885
r329 16 17 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.445 $Y2=2.885
r330 15 93 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.81
+ $X2=1.352 $Y2=2.885
r331 14 126 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=1.935
r332 14 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=2.81
r333 11 93 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.352 $Y2=2.885
r334 11 13 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r335 7 125 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.935
r336 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r337 2 109 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=0.135 $Y=3.085 $X2=0.26 $Y2=5.835
r338 2 107 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=0.135 $Y=3.085 $X2=0.26 $Y2=3.795
r339 1 117 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__OR2_8%Y 1 2 3 4 5 6 7 8 25 26 28 30 32 35 36 37
+ 38 39 40 41 42 43 46 47 53 59 65 67 71 73 85 97 109
c160 53 0 1.37149e-19 $X=1.55 $Y=2.59
c161 46 0 1.33323e-19 $X=4.13 $Y=1.595
c162 40 0 1.33323e-19 $X=3.27 $Y=1.595
c163 37 0 2.66647e-19 $X=2.555 $Y=1.48
c164 25 0 1.33323e-19 $X=1.55 $Y=1.595
r165 116 118 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.13 $Y=3.455
+ $X2=4.13 $Y2=5.835
r166 104 106 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.27 $Y=3.455
+ $X2=3.27 $Y2=5.835
r167 92 94 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r168 80 82 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r169 71 116 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.13 $Y=2.59
+ $X2=4.13 $Y2=3.455
r170 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=2.59
+ $X2=4.13 $Y2=2.59
r171 68 109 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.13 $Y=1.48
+ $X2=4.13 $Y2=0.825
r172 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=1.48
+ $X2=4.13 $Y2=1.48
r173 65 104 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.27 $Y=2.59
+ $X2=3.27 $Y2=3.455
r174 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.59
+ $X2=3.27 $Y2=2.59
r175 62 97 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.27 $Y=1.48
+ $X2=3.27 $Y2=0.825
r176 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.48
+ $X2=3.27 $Y2=1.48
r177 59 92 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.41 $Y=2.59
+ $X2=2.41 $Y2=3.455
r178 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.59
+ $X2=2.41 $Y2=2.59
r179 56 85 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.41 $Y=1.48
+ $X2=2.41 $Y2=0.825
r180 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.48
+ $X2=2.41 $Y2=1.48
r181 53 80 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r182 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r183 50 73 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r184 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r185 47 70 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=2.475
+ $X2=4.13 $Y2=2.59
r186 46 67 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.595
+ $X2=4.13 $Y2=1.48
r187 46 47 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=4.13 $Y=1.595
+ $X2=4.13 $Y2=2.475
r188 43 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=2.59
+ $X2=3.27 $Y2=2.59
r189 42 70 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=2.59
+ $X2=4.13 $Y2=2.59
r190 42 43 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=2.59
+ $X2=3.415 $Y2=2.59
r191 41 64 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.475
+ $X2=3.27 $Y2=2.59
r192 40 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.595
+ $X2=3.27 $Y2=1.48
r193 40 41 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=3.27 $Y=1.595
+ $X2=3.27 $Y2=2.475
r194 39 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.59
+ $X2=2.41 $Y2=2.59
r195 38 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.59
+ $X2=3.27 $Y2=2.59
r196 38 39 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.59
+ $X2=2.555 $Y2=2.59
r197 37 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.48
+ $X2=2.41 $Y2=1.48
r198 36 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.48
+ $X2=3.27 $Y2=1.48
r199 36 37 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.48
+ $X2=2.555 $Y2=1.48
r200 35 58 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.475
+ $X2=2.41 $Y2=2.59
r201 34 55 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=1.48
r202 34 35 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=2.475
r203 33 52 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.59
+ $X2=1.55 $Y2=2.59
r204 32 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.59
+ $X2=2.41 $Y2=2.59
r205 32 33 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.59
+ $X2=1.695 $Y2=2.59
r206 31 49 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.48
+ $X2=1.55 $Y2=1.48
r207 30 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=2.41 $Y2=1.48
r208 30 31 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=1.695 $Y2=1.48
r209 26 52 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r210 26 28 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r211 25 49 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r212 25 28 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r213 8 118 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.99
+ $Y=3.085 $X2=4.13 $Y2=5.835
r214 8 116 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.99
+ $Y=3.085 $X2=4.13 $Y2=3.455
r215 7 106 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=5.835
r216 7 104 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=3.455
r217 6 94 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r218 6 92 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r219 5 82 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r220 5 80 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r221 4 109 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.825
r222 3 97 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.825
r223 2 85 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r224 1 73 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

