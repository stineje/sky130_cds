magic
tech sky130A
magscale 1 2
timestamp 1606864594
<< checkpaint >>
rect -1210 -1243 3248 2575
<< nwell >>
rect -10 581 2090 1341
<< nmos >>
rect 80 115 110 315
rect 272 115 302 263
rect 370 115 400 315
rect 442 115 472 315
rect 632 115 662 315
rect 704 115 734 315
rect 824 115 854 315
rect 896 115 926 315
rect 982 115 1012 315
rect 1054 115 1084 315
rect 1174 115 1204 315
rect 1246 115 1276 315
rect 1332 115 1362 315
rect 1522 115 1552 315
rect 1594 115 1624 315
rect 1692 115 1722 263
rect 1884 115 1914 263
rect 1970 115 2000 263
<< pmoshvt >>
rect 80 617 110 1217
rect 270 617 300 1217
rect 356 617 386 1217
rect 442 617 472 1217
rect 632 617 662 1217
rect 704 617 734 1217
rect 824 617 854 1217
rect 896 617 926 1217
rect 982 617 1012 1217
rect 1054 617 1084 1217
rect 1174 617 1204 1217
rect 1246 617 1276 1217
rect 1332 617 1362 1217
rect 1522 617 1552 1217
rect 1608 617 1638 1217
rect 1694 617 1724 1217
rect 1884 817 1914 1217
rect 1970 817 2000 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 163 315
rect 110 131 121 267
rect 155 131 163 267
rect 317 267 370 315
rect 317 263 325 267
rect 110 115 163 131
rect 219 199 272 263
rect 219 131 227 199
rect 261 131 272 199
rect 219 115 272 131
rect 302 131 325 263
rect 359 131 370 267
rect 302 115 370 131
rect 400 115 442 315
rect 472 267 525 315
rect 472 131 483 267
rect 517 131 525 267
rect 472 115 525 131
rect 579 267 632 315
rect 579 131 587 267
rect 621 131 632 267
rect 579 115 632 131
rect 662 115 704 315
rect 734 267 824 315
rect 734 131 745 267
rect 813 131 824 267
rect 734 115 824 131
rect 854 115 896 315
rect 926 199 982 315
rect 926 131 937 199
rect 971 131 982 199
rect 926 115 982 131
rect 1012 115 1054 315
rect 1084 267 1174 315
rect 1084 131 1095 267
rect 1163 131 1174 267
rect 1084 115 1174 131
rect 1204 115 1246 315
rect 1276 267 1332 315
rect 1276 131 1287 267
rect 1321 131 1332 267
rect 1276 115 1332 131
rect 1362 267 1415 315
rect 1362 131 1373 267
rect 1407 131 1415 267
rect 1362 115 1415 131
rect 1469 267 1522 315
rect 1469 131 1477 267
rect 1511 131 1522 267
rect 1469 115 1522 131
rect 1552 115 1594 315
rect 1624 267 1677 315
rect 1624 131 1635 267
rect 1669 263 1677 267
rect 1669 131 1692 263
rect 1624 115 1692 131
rect 1722 199 1775 263
rect 1722 131 1733 199
rect 1767 131 1775 199
rect 1722 115 1775 131
rect 1831 199 1884 263
rect 1831 131 1839 199
rect 1873 131 1884 199
rect 1831 115 1884 131
rect 1914 199 1970 263
rect 1914 131 1925 199
rect 1959 131 1970 199
rect 1914 115 1970 131
rect 2000 199 2053 263
rect 2000 131 2011 199
rect 2045 131 2053 199
rect 2000 115 2053 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 163 1217
rect 110 657 121 1201
rect 155 657 163 1201
rect 110 617 163 657
rect 217 1201 270 1217
rect 217 725 225 1201
rect 259 725 270 1201
rect 217 617 270 725
rect 300 1201 356 1217
rect 300 725 311 1201
rect 345 725 356 1201
rect 300 617 356 725
rect 386 1201 442 1217
rect 386 793 397 1201
rect 431 793 442 1201
rect 386 617 442 793
rect 472 1201 525 1217
rect 472 725 483 1201
rect 517 725 525 1201
rect 472 617 525 725
rect 579 1201 632 1217
rect 579 725 587 1201
rect 621 725 632 1201
rect 579 617 632 725
rect 662 617 704 1217
rect 734 1201 824 1217
rect 734 657 745 1201
rect 813 657 824 1201
rect 734 617 824 657
rect 854 617 896 1217
rect 926 1201 982 1217
rect 926 725 937 1201
rect 971 725 982 1201
rect 926 617 982 725
rect 1012 617 1054 1217
rect 1084 1201 1174 1217
rect 1084 725 1095 1201
rect 1163 725 1174 1201
rect 1084 617 1174 725
rect 1204 617 1246 1217
rect 1276 1201 1332 1217
rect 1276 657 1287 1201
rect 1321 657 1332 1201
rect 1276 617 1332 657
rect 1362 1201 1415 1217
rect 1362 657 1373 1201
rect 1407 657 1415 1201
rect 1362 617 1415 657
rect 1469 1201 1522 1217
rect 1469 725 1477 1201
rect 1511 725 1522 1201
rect 1469 617 1522 725
rect 1552 1201 1608 1217
rect 1552 793 1563 1201
rect 1597 793 1608 1201
rect 1552 617 1608 793
rect 1638 1201 1694 1217
rect 1638 725 1649 1201
rect 1683 725 1694 1201
rect 1638 617 1694 725
rect 1724 1201 1777 1217
rect 1724 725 1735 1201
rect 1769 725 1777 1201
rect 1831 1201 1884 1217
rect 1831 861 1839 1201
rect 1873 861 1884 1201
rect 1831 817 1884 861
rect 1914 1201 1970 1217
rect 1914 861 1925 1201
rect 1959 861 1970 1201
rect 1914 817 1970 861
rect 2000 1201 2053 1217
rect 2000 861 2011 1201
rect 2045 861 2053 1201
rect 2000 817 2053 861
rect 1724 617 1777 725
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 227 131 261 199
rect 325 131 359 267
rect 483 131 517 267
rect 587 131 621 267
rect 745 131 813 267
rect 937 131 971 199
rect 1095 131 1163 267
rect 1287 131 1321 267
rect 1373 131 1407 267
rect 1477 131 1511 267
rect 1635 131 1669 267
rect 1733 131 1767 199
rect 1839 131 1873 199
rect 1925 131 1959 199
rect 2011 131 2045 199
<< pdiffc >>
rect 35 793 69 1201
rect 121 657 155 1201
rect 225 725 259 1201
rect 311 725 345 1201
rect 397 793 431 1201
rect 483 725 517 1201
rect 587 725 621 1201
rect 745 657 813 1201
rect 937 725 971 1201
rect 1095 725 1163 1201
rect 1287 657 1321 1201
rect 1373 657 1407 1201
rect 1477 725 1511 1201
rect 1563 793 1597 1201
rect 1649 725 1683 1201
rect 1735 725 1769 1201
rect 1839 861 1873 1201
rect 1925 861 1959 1201
rect 2011 861 2045 1201
<< psubdiff >>
rect 26 27 50 61
rect 84 27 108 61
rect 162 27 186 61
rect 220 27 244 61
rect 298 27 322 61
rect 356 27 380 61
rect 434 27 458 61
rect 492 27 516 61
rect 570 27 594 61
rect 628 27 652 61
rect 706 27 730 61
rect 764 27 788 61
rect 842 27 866 61
rect 900 27 924 61
rect 978 27 1002 61
rect 1036 27 1060 61
rect 1114 27 1138 61
rect 1172 27 1196 61
rect 1250 27 1274 61
rect 1308 27 1332 61
rect 1386 27 1410 61
rect 1444 27 1468 61
rect 1522 27 1546 61
rect 1580 27 1604 61
rect 1658 27 1682 61
rect 1716 27 1740 61
rect 1794 27 1818 61
rect 1852 27 1876 61
rect 1930 27 1954 61
rect 1988 27 2012 61
<< nsubdiff >>
rect 26 1271 50 1305
rect 84 1271 108 1305
rect 162 1271 186 1305
rect 220 1271 244 1305
rect 298 1271 322 1305
rect 356 1271 380 1305
rect 434 1271 458 1305
rect 492 1271 516 1305
rect 570 1271 594 1305
rect 628 1271 652 1305
rect 706 1271 730 1305
rect 764 1271 788 1305
rect 842 1271 866 1305
rect 900 1271 924 1305
rect 978 1271 1002 1305
rect 1036 1271 1060 1305
rect 1114 1271 1138 1305
rect 1172 1271 1196 1305
rect 1250 1271 1274 1305
rect 1308 1271 1332 1305
rect 1386 1271 1410 1305
rect 1444 1271 1468 1305
rect 1522 1271 1546 1305
rect 1580 1271 1604 1305
rect 1658 1271 1682 1305
rect 1716 1271 1740 1305
rect 1794 1271 1818 1305
rect 1852 1271 1876 1305
rect 1930 1271 1954 1305
rect 1988 1271 2012 1305
<< psubdiffcont >>
rect 50 27 84 61
rect 186 27 220 61
rect 322 27 356 61
rect 458 27 492 61
rect 594 27 628 61
rect 730 27 764 61
rect 866 27 900 61
rect 1002 27 1036 61
rect 1138 27 1172 61
rect 1274 27 1308 61
rect 1410 27 1444 61
rect 1546 27 1580 61
rect 1682 27 1716 61
rect 1818 27 1852 61
rect 1954 27 1988 61
<< nsubdiffcont >>
rect 50 1271 84 1305
rect 186 1271 220 1305
rect 322 1271 356 1305
rect 458 1271 492 1305
rect 594 1271 628 1305
rect 730 1271 764 1305
rect 866 1271 900 1305
rect 1002 1271 1036 1305
rect 1138 1271 1172 1305
rect 1274 1271 1308 1305
rect 1410 1271 1444 1305
rect 1546 1271 1580 1305
rect 1682 1271 1716 1305
rect 1818 1271 1852 1305
rect 1954 1271 1988 1305
<< poly >>
rect 80 1217 110 1243
rect 270 1217 300 1243
rect 356 1217 386 1243
rect 442 1217 472 1243
rect 632 1217 662 1243
rect 704 1217 734 1243
rect 824 1217 854 1243
rect 896 1217 926 1243
rect 982 1217 1012 1243
rect 1054 1217 1084 1243
rect 1174 1217 1204 1243
rect 1246 1217 1276 1243
rect 1332 1217 1362 1243
rect 1522 1217 1552 1243
rect 1608 1217 1638 1243
rect 1694 1217 1724 1243
rect 1884 1217 1914 1243
rect 1970 1217 2000 1243
rect 80 494 110 617
rect 270 579 300 617
rect 243 549 300 579
rect 79 478 133 494
rect 79 444 89 478
rect 123 444 133 478
rect 79 428 133 444
rect 79 427 110 428
rect 80 315 110 427
rect 243 351 273 549
rect 356 507 386 617
rect 442 586 472 617
rect 432 570 486 586
rect 432 536 442 570
rect 476 536 486 570
rect 432 520 486 536
rect 315 491 386 507
rect 315 457 325 491
rect 359 457 386 491
rect 315 441 386 457
rect 356 385 386 441
rect 356 355 400 385
rect 219 335 273 351
rect 219 301 229 335
rect 263 317 273 335
rect 263 301 302 317
rect 370 315 400 355
rect 442 315 472 520
rect 632 477 662 617
rect 704 586 734 617
rect 704 570 758 586
rect 704 536 714 570
rect 748 536 758 570
rect 704 520 758 536
rect 632 461 686 477
rect 824 475 854 617
rect 896 580 926 617
rect 982 580 1012 617
rect 896 570 1012 580
rect 896 536 928 570
rect 962 536 1012 570
rect 896 526 1012 536
rect 1054 475 1084 617
rect 1174 586 1204 617
rect 1150 570 1204 586
rect 1150 536 1160 570
rect 1194 536 1204 570
rect 1150 520 1204 536
rect 632 427 642 461
rect 676 427 686 461
rect 632 411 686 427
rect 728 445 1180 475
rect 632 315 662 411
rect 728 367 758 445
rect 1150 403 1180 445
rect 1246 471 1276 617
rect 1332 586 1362 617
rect 1332 570 1403 586
rect 1522 580 1552 617
rect 1332 556 1359 570
rect 1343 536 1359 556
rect 1393 536 1403 570
rect 1343 520 1403 536
rect 1486 570 1552 580
rect 1486 536 1502 570
rect 1536 536 1552 570
rect 1486 526 1552 536
rect 1246 455 1300 471
rect 1246 421 1256 455
rect 1290 421 1300 455
rect 1246 405 1300 421
rect 704 337 758 367
rect 800 387 854 403
rect 800 353 810 387
rect 844 353 854 387
rect 800 337 854 353
rect 704 315 734 337
rect 824 315 854 337
rect 896 387 1012 397
rect 896 353 928 387
rect 962 353 1012 387
rect 896 343 1012 353
rect 896 315 926 343
rect 982 315 1012 343
rect 1054 387 1108 403
rect 1054 353 1064 387
rect 1098 353 1108 387
rect 1054 337 1108 353
rect 1150 387 1204 403
rect 1150 353 1160 387
rect 1194 353 1204 387
rect 1150 337 1204 353
rect 1054 315 1084 337
rect 1174 315 1204 337
rect 1246 315 1276 405
rect 1343 367 1373 520
rect 1332 337 1373 367
rect 1486 370 1516 526
rect 1608 484 1638 617
rect 1694 579 1724 617
rect 1884 601 1914 817
rect 1694 549 1775 579
rect 1576 468 1638 484
rect 1576 434 1588 468
rect 1622 434 1638 468
rect 1576 418 1638 434
rect 1486 338 1552 370
rect 1332 315 1362 337
rect 1522 315 1552 338
rect 1594 315 1624 418
rect 1745 351 1775 549
rect 1874 571 1914 601
rect 1874 471 1904 571
rect 1970 512 2000 817
rect 1849 455 1904 471
rect 1849 421 1859 455
rect 1893 421 1904 455
rect 1946 496 2000 512
rect 1946 462 1956 496
rect 1990 462 2000 496
rect 1946 446 2000 462
rect 1849 405 1904 421
rect 1874 360 1904 405
rect 1745 335 1799 351
rect 1745 315 1755 335
rect 219 285 302 301
rect 272 263 302 285
rect 1692 301 1755 315
rect 1789 301 1799 335
rect 1874 330 1914 360
rect 1692 285 1799 301
rect 1692 263 1722 285
rect 1884 263 1914 330
rect 1970 263 2000 446
rect 80 89 110 115
rect 272 89 302 115
rect 370 89 400 115
rect 442 89 472 115
rect 632 89 662 115
rect 704 89 734 115
rect 824 89 854 115
rect 896 89 926 115
rect 982 89 1012 115
rect 1054 89 1084 115
rect 1174 89 1204 115
rect 1246 89 1276 115
rect 1332 89 1362 115
rect 1522 89 1552 115
rect 1594 89 1624 115
rect 1692 89 1722 115
rect 1884 89 1914 115
rect 1970 89 2000 115
<< polycont >>
rect 89 444 123 478
rect 442 536 476 570
rect 325 457 359 491
rect 229 301 263 335
rect 714 536 748 570
rect 928 536 962 570
rect 1160 536 1194 570
rect 642 427 676 461
rect 1359 536 1393 570
rect 1502 536 1536 570
rect 1256 421 1290 455
rect 810 353 844 387
rect 928 353 962 387
rect 1064 353 1098 387
rect 1160 353 1194 387
rect 1588 434 1622 468
rect 1859 421 1893 455
rect 1956 462 1990 496
rect 1755 301 1789 335
<< locali >>
rect 0 1311 2090 1332
rect 0 1271 50 1311
rect 84 1271 186 1311
rect 220 1271 322 1311
rect 356 1271 458 1311
rect 492 1271 594 1311
rect 628 1271 730 1311
rect 764 1271 866 1311
rect 900 1271 1002 1311
rect 1036 1271 1138 1311
rect 1172 1271 1274 1311
rect 1308 1271 1410 1311
rect 1444 1271 1546 1311
rect 1580 1271 1682 1311
rect 1716 1271 1818 1311
rect 1852 1271 1954 1311
rect 1988 1271 2090 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 47 494 81 649
rect 121 565 155 657
rect 225 1201 259 1217
rect 121 531 191 565
rect 47 478 123 494
rect 47 444 89 478
rect 89 428 123 444
rect 157 335 191 531
rect 225 421 259 725
rect 311 1201 345 1217
rect 397 1201 431 1271
rect 397 777 431 793
rect 483 1201 517 1217
rect 345 725 483 743
rect 311 709 517 725
rect 587 1201 621 1271
rect 587 709 621 725
rect 745 1201 813 1217
rect 937 1201 971 1271
rect 937 709 971 725
rect 1095 1201 1163 1217
rect 813 657 816 675
rect 745 654 816 657
rect 1095 654 1163 725
rect 442 620 816 654
rect 996 620 1163 654
rect 1287 1201 1321 1271
rect 1287 641 1321 657
rect 1373 1201 1407 1217
rect 1477 1201 1511 1217
rect 1563 1201 1597 1271
rect 1563 777 1597 793
rect 1649 1201 1683 1217
rect 1511 725 1649 743
rect 1477 709 1683 725
rect 1735 1201 1769 1217
rect 1373 654 1407 657
rect 1373 620 1461 654
rect 325 491 359 575
rect 442 570 476 620
rect 309 457 325 491
rect 359 457 375 491
rect 225 387 359 421
rect 121 301 229 335
rect 263 301 279 335
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 301
rect 325 267 359 353
rect 442 370 476 536
rect 714 570 748 586
rect 714 535 748 536
rect 928 570 962 586
rect 748 501 844 535
rect 642 461 676 477
rect 642 411 676 427
rect 810 387 844 501
rect 928 387 962 536
rect 442 336 776 370
rect 810 337 844 353
rect 928 337 962 353
rect 996 387 1030 620
rect 1160 570 1194 586
rect 1160 535 1194 536
rect 742 283 776 336
rect 996 303 1030 353
rect 1064 501 1160 535
rect 1359 570 1393 586
rect 1359 535 1393 536
rect 1064 387 1098 501
rect 1427 455 1461 620
rect 1240 421 1256 455
rect 1290 421 1306 455
rect 1373 421 1461 455
rect 1502 570 1536 586
rect 1373 387 1407 421
rect 1144 353 1160 387
rect 1194 353 1407 387
rect 1502 387 1536 536
rect 1570 484 1604 575
rect 1570 468 1638 484
rect 1570 434 1588 468
rect 1622 434 1638 468
rect 1735 455 1769 725
rect 1839 1201 1873 1217
rect 1839 609 1873 861
rect 1925 1201 1959 1271
rect 1925 845 1959 861
rect 2011 1201 2045 1217
rect 2011 683 2045 861
rect 2044 666 2045 683
rect 2044 649 2068 666
rect 2011 632 2068 649
rect 1839 570 1873 575
rect 1839 536 1990 570
rect 1956 496 1990 536
rect 1672 421 1859 455
rect 1893 421 1909 455
rect 1672 399 1706 421
rect 1635 365 1706 399
rect 1956 387 1990 462
rect 1064 337 1098 353
rect 121 115 155 131
rect 227 199 261 215
rect 227 61 261 131
rect 325 115 359 131
rect 483 267 517 283
rect 483 61 517 131
rect 587 267 621 283
rect 742 267 813 283
rect 996 269 1163 303
rect 742 249 745 267
rect 587 61 621 131
rect 1095 267 1163 269
rect 745 115 813 131
rect 937 199 971 215
rect 937 61 971 131
rect 1095 115 1163 131
rect 1287 267 1321 283
rect 1287 61 1321 131
rect 1373 267 1407 353
rect 1373 115 1407 131
rect 1477 267 1511 283
rect 1477 61 1511 131
rect 1635 267 1669 365
rect 1839 353 1990 387
rect 1739 301 1755 335
rect 1789 301 1805 335
rect 1635 115 1669 131
rect 1733 199 1767 215
rect 1733 61 1767 131
rect 1839 199 1873 353
rect 2034 320 2068 632
rect 2011 286 2068 320
rect 1839 115 1873 131
rect 1925 199 1959 215
rect 1925 61 1959 131
rect 2011 199 2045 286
rect 2011 115 2045 131
rect 0 21 50 61
rect 84 21 186 61
rect 220 21 322 61
rect 356 21 458 61
rect 492 21 594 61
rect 628 21 730 61
rect 764 21 866 61
rect 900 21 1002 61
rect 1036 21 1138 61
rect 1172 21 1274 61
rect 1308 21 1410 61
rect 1444 21 1546 61
rect 1580 21 1682 61
rect 1716 21 1818 61
rect 1852 21 1954 61
rect 1988 21 2090 61
rect 0 0 2090 21
<< viali >>
rect 50 1305 84 1311
rect 50 1277 84 1305
rect 186 1305 220 1311
rect 186 1277 220 1305
rect 322 1305 356 1311
rect 322 1277 356 1305
rect 458 1305 492 1311
rect 458 1277 492 1305
rect 594 1305 628 1311
rect 594 1277 628 1305
rect 730 1305 764 1311
rect 730 1277 764 1305
rect 866 1305 900 1311
rect 866 1277 900 1305
rect 1002 1305 1036 1311
rect 1002 1277 1036 1305
rect 1138 1305 1172 1311
rect 1138 1277 1172 1305
rect 1274 1305 1308 1311
rect 1274 1277 1308 1305
rect 1410 1305 1444 1311
rect 1410 1277 1444 1305
rect 1546 1305 1580 1311
rect 1546 1277 1580 1305
rect 1682 1305 1716 1311
rect 1682 1277 1716 1305
rect 1818 1305 1852 1311
rect 1818 1277 1852 1305
rect 1954 1305 1988 1311
rect 1954 1277 1988 1305
rect 47 649 81 683
rect 325 575 359 609
rect 325 353 359 387
rect 229 301 263 313
rect 229 279 263 301
rect 714 501 748 535
rect 642 427 676 461
rect 910 353 928 387
rect 928 353 944 387
rect 996 353 1030 387
rect 1160 501 1194 535
rect 1359 501 1393 535
rect 1256 421 1290 455
rect 1570 575 1604 609
rect 2010 649 2044 683
rect 1839 575 1873 609
rect 1859 421 1893 455
rect 1502 353 1536 387
rect 1755 301 1789 313
rect 1755 279 1789 301
rect 50 27 84 55
rect 50 21 84 27
rect 186 27 220 55
rect 186 21 220 27
rect 322 27 356 55
rect 322 21 356 27
rect 458 27 492 55
rect 458 21 492 27
rect 594 27 628 55
rect 594 21 628 27
rect 730 27 764 55
rect 730 21 764 27
rect 866 27 900 55
rect 866 21 900 27
rect 1002 27 1036 55
rect 1002 21 1036 27
rect 1138 27 1172 55
rect 1138 21 1172 27
rect 1274 27 1308 55
rect 1274 21 1308 27
rect 1410 27 1444 55
rect 1410 21 1444 27
rect 1546 27 1580 55
rect 1546 21 1580 27
rect 1682 27 1716 55
rect 1682 21 1716 27
rect 1818 27 1852 55
rect 1818 21 1852 27
rect 1954 27 1988 55
rect 1954 21 1988 27
<< metal1 >>
rect 0 1311 2090 1332
rect 0 1277 50 1311
rect 84 1277 186 1311
rect 220 1277 322 1311
rect 356 1277 458 1311
rect 492 1277 594 1311
rect 628 1277 730 1311
rect 764 1277 866 1311
rect 900 1277 1002 1311
rect 1036 1277 1138 1311
rect 1172 1277 1274 1311
rect 1308 1277 1410 1311
rect 1444 1277 1546 1311
rect 1580 1277 1682 1311
rect 1716 1277 1818 1311
rect 1852 1277 1954 1311
rect 1988 1277 2090 1311
rect 0 1271 2090 1277
rect 35 683 93 689
rect 1998 683 2056 689
rect 35 649 47 683
rect 81 649 127 683
rect 1976 649 2010 683
rect 2044 649 2056 683
rect 35 643 93 649
rect 1998 643 2056 649
rect 313 609 371 615
rect 1558 609 1616 615
rect 1827 609 1885 615
rect 313 575 325 609
rect 359 575 1570 609
rect 1604 575 1616 609
rect 1804 575 1839 609
rect 1873 575 1885 609
rect 313 569 371 575
rect 1558 569 1616 575
rect 1827 569 1885 575
rect 702 535 760 541
rect 1148 535 1206 541
rect 1347 535 1405 541
rect 702 501 714 535
rect 748 501 1160 535
rect 1194 501 1359 535
rect 1393 501 1405 535
rect 702 495 760 501
rect 1148 495 1206 501
rect 1347 495 1405 501
rect 630 461 688 467
rect 630 427 642 461
rect 676 427 710 461
rect 1244 455 1302 461
rect 1847 455 1905 461
rect 630 421 688 427
rect 1244 421 1256 455
rect 1290 421 1859 455
rect 1893 421 1905 455
rect 1244 415 1302 421
rect 1847 415 1905 421
rect 313 387 371 393
rect 898 387 956 393
rect 313 353 325 387
rect 359 353 910 387
rect 944 353 956 387
rect 313 347 371 353
rect 898 347 956 353
rect 984 387 1042 393
rect 1490 387 1548 393
rect 984 353 996 387
rect 1030 353 1502 387
rect 1536 353 1548 387
rect 984 347 1042 353
rect 1490 347 1548 353
rect 217 313 275 319
rect 1743 313 1801 319
rect 217 279 229 313
rect 263 279 1755 313
rect 1789 279 1801 313
rect 217 273 275 279
rect 1743 273 1801 279
rect 0 55 2090 61
rect 0 21 50 55
rect 84 21 186 55
rect 220 21 322 55
rect 356 21 458 55
rect 492 21 594 55
rect 628 21 730 55
rect 764 21 866 55
rect 900 21 1002 55
rect 1036 21 1138 55
rect 1172 21 1274 55
rect 1308 21 1410 55
rect 1444 21 1546 55
rect 1580 21 1682 55
rect 1716 21 1818 55
rect 1852 21 1954 55
rect 1988 21 2090 55
rect 0 0 2090 21
<< labels >>
rlabel metal1 659 444 659 444 1 D
port 1 n
rlabel metal1 1376 518 1376 518 1 CK
port 2 n
rlabel metal1 1857 592 1857 592 1 QN
port 3 n
rlabel metal1 2027 666 2027 666 1 Q
port 4 n
rlabel metal1 1587 592 1587 592 1 SN
port 5 n
rlabel metal1 65 666 65 666 1 RN
port 6 n
rlabel viali 67 48 67 48 1 gnd
rlabel viali 67 1284 67 1284 1 vdd
<< end >>
