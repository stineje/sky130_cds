* File: sky130_osu_sc_15T_ls__tnbufi_1.pex.spice
* Created: Fri Nov 12 15:00:28 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__TNBUFI_1%GND 1 17 19 26 35 38
r34 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r35 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r36 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r37 24 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.865
r38 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r39 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r40 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r41 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r42 1 26 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TNBUFI_1%VDD 1 13 15 21 27 31 34
r19 31 34 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r20 27 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r21 25 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r22 25 27 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397 $X2=1.02
+ $Y2=5.397
r23 21 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=3.545
+ $X2=0.69 $Y2=4.565
r24 19 29 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r25 19 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r26 15 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r27 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r28 13 27 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r29 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r30 1 24 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r31 1 21 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.545
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TNBUFI_1%A_27_115# 1 3 11 16 20 24 28 30 33
r44 29 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.915
+ $X2=0.26 $Y2=1.915
r45 28 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=1.915
+ $X2=0.69 $Y2=1.915
r46 28 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.915
+ $X2=0.345 $Y2=1.915
r47 24 26 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r48 22 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2 $X2=0.26
+ $Y2=1.915
r49 22 24 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=0.26 $Y=2 $X2=0.26
+ $Y2=3.205
r50 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.83 $X2=0.26
+ $Y2=1.915
r51 18 20 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=0.26 $Y=1.83
+ $X2=0.26 $Y2=0.865
r52 14 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.915 $X2=0.69 $Y2=1.915
r53 14 16 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=1.915
+ $X2=0.905 $Y2=1.915
r54 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.75
+ $X2=0.905 $Y2=1.915
r55 9 11 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.905 $Y=1.75
+ $X2=0.905 $Y2=0.945
r56 3 26 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r57 3 24 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r58 1 20 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TNBUFI_1%OE 3 5 6 8 11 14 19 25
r42 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.7 $X2=0.69
+ $Y2=2.7
r43 19 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.69 $Y=2.505
+ $X2=0.69 $Y2=2.7
r44 17 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.505 $X2=0.69 $Y2=2.505
r45 12 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.475 $Y2=1.465
r46 6 17 49.2914 $w=4.58e-07 $l=4.23124e-07 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.587 $Y2=2.505
r47 6 11 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=3.825
r48 6 8 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=3.825
r49 3 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.475 $Y2=1.465
r50 3 5 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.475 $Y2=0.945
r51 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=1.54 $X2=0.27
+ $Y2=1.465
r52 1 6 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.54 $X2=0.27
+ $Y2=2.6
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TNBUFI_1%A 3 7 10 15 20 23
r47 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.83
+ $X2=1.325 $Y2=1.83
r48 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=3.07
+ $X2=1.14 $Y2=3.07
r49 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.915
+ $X2=1.14 $Y2=1.83
r50 13 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=1.915
+ $X2=1.14 $Y2=3.07
r51 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.83 $X2=1.325 $Y2=1.83
r52 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.83
+ $X2=1.325 $Y2=1.995
r53 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.83
+ $X2=1.325 $Y2=1.665
r54 7 12 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=1.265 $Y=3.825
+ $X2=1.265 $Y2=1.995
r55 3 11 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.265 $Y=0.945
+ $X2=1.265 $Y2=1.665
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TNBUFI_1%Y 1 3 10 16 26 29 32
r32 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.215
+ $X2=1.48 $Y2=2.33
r33 24 26 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.215
+ $X2=1.48 $Y2=1.56
r34 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.335
+ $X2=1.48 $Y2=1.22
r35 23 26 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.335
+ $X2=1.48 $Y2=1.56
r36 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.48 $Y=3.205
+ $X2=1.48 $Y2=4.565
r37 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.33
+ $X2=1.48 $Y2=2.33
r38 16 19 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.48 $Y=2.33
+ $X2=1.48 $Y2=3.205
r39 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.22
+ $X2=1.48 $Y2=1.22
r40 10 13 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.48 $Y=0.865
+ $X2=1.48 $Y2=1.22
r41 3 21 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.48 $Y2=4.565
r42 3 19 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.48 $Y2=3.205
r43 1 10 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.865
.ends

