* File: sky130_osu_sc_18T_hs__addf_l.pxi.spice
* Created: Thu Oct 29 17:05:28 2020
* 
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%GND N_GND_M1012_d N_GND_M1027_d N_GND_M1024_d
+ N_GND_M1006_d N_GND_M1021_s N_GND_M1012_b N_GND_c_28_p N_GND_c_3_p N_GND_c_4_p
+ N_GND_c_34_p N_GND_c_72_p N_GND_c_39_p N_GND_c_25_p N_GND_c_135_p
+ N_GND_c_106_p N_GND_c_29_p GND N_GND_c_5_p PM_SKY130_OSU_SC_18T_HS__ADDF_L%GND
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%VDD N_VDD_M1010_d N_VDD_M1026_d N_VDD_M1022_d
+ N_VDD_M1002_d N_VDD_M1008_s N_VDD_M1010_b N_VDD_c_181_p N_VDD_c_185_p
+ N_VDD_c_186_p N_VDD_c_193_p N_VDD_c_212_p N_VDD_c_196_p N_VDD_c_197_p
+ N_VDD_c_244_p N_VDD_c_233_p N_VDD_c_182_p VDD N_VDD_c_183_p N_VDD_c_235_p
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%VDD
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%A N_A_M1012_g N_A_M1010_g N_A_c_288_n
+ N_A_M1027_g N_A_c_332_n N_A_M1026_g N_A_c_292_n N_A_c_294_n N_A_c_295_n
+ N_A_c_296_n N_A_c_297_n N_A_M1020_g N_A_c_339_n N_A_M1019_g N_A_M1006_g
+ N_A_M1002_g N_A_c_298_n N_A_c_299_n N_A_c_300_n N_A_c_301_n N_A_c_303_n
+ N_A_c_304_n N_A_c_305_n A N_A_c_306_n N_A_c_307_n N_A_c_309_n N_A_c_310_n
+ N_A_c_312_n N_A_c_313_n N_A_c_317_n N_A_c_318_n N_A_c_322_n N_A_c_324_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%A
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%B N_B_M1003_g N_B_M1000_g N_B_M1025_g
+ N_B_M1023_g N_B_M1024_g N_B_M1022_g N_B_M1017_g N_B_M1016_g N_B_c_508_n
+ N_B_c_509_n N_B_c_510_n N_B_c_511_n N_B_c_512_n N_B_c_513_n B N_B_c_514_n
+ N_B_c_515_n N_B_c_516_n N_B_c_517_n N_B_c_518_n N_B_c_519_n N_B_c_520_n
+ N_B_c_521_n N_B_c_522_n N_B_c_523_n N_B_c_527_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%B
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%CI N_CI_M1005_g N_CI_M1004_g N_CI_M1014_g
+ N_CI_M1011_g N_CI_M1009_g N_CI_M1007_g N_CI_c_736_n N_CI_c_737_n N_CI_c_738_n
+ N_CI_c_739_n N_CI_c_740_n N_CI_c_741_n CI N_CI_c_743_n N_CI_c_744_n
+ N_CI_c_745_n N_CI_c_746_n N_CI_c_747_n N_CI_c_748_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%CI
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%CON N_CON_M1005_d N_CON_M1004_d N_CON_c_906_n
+ N_CON_M1015_g N_CON_M1013_g N_CON_M1021_g N_CON_M1008_g N_CON_c_945_n
+ N_CON_c_913_n N_CON_c_914_n N_CON_c_915_n N_CON_c_916_n N_CON_c_917_n
+ N_CON_c_918_n N_CON_c_919_n N_CON_c_923_n N_CON_c_925_n N_CON_c_928_n
+ N_CON_c_929_n CON N_CON_c_932_n N_CON_c_936_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%CON
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_784_115# N_A_784_115#_M1015_d
+ N_A_784_115#_M1013_d N_A_784_115#_M1018_g N_A_784_115#_M1001_g
+ N_A_784_115#_c_1096_n N_A_784_115#_c_1097_n N_A_784_115#_c_1098_n
+ N_A_784_115#_c_1099_n N_A_784_115#_c_1113_n N_A_784_115#_c_1114_n
+ N_A_784_115#_c_1117_n N_A_784_115#_c_1102_n N_A_784_115#_c_1120_n
+ N_A_784_115#_c_1103_n N_A_784_115#_c_1105_n N_A_784_115#_c_1106_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_784_115#
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_27_617# N_A_27_617#_M1010_s
+ N_A_27_617#_M1000_d N_A_27_617#_c_1219_n N_A_27_617#_c_1222_n
+ N_A_27_617#_c_1224_n PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_27_617#
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_526_617# N_A_526_617#_M1019_d
+ N_A_526_617#_M1011_d N_A_526_617#_c_1232_n N_A_526_617#_c_1235_n
+ N_A_526_617#_c_1237_n PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_526_617#
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%S N_S_M1018_d N_S_M1001_d N_S_c_1246_n
+ N_S_c_1251_n N_S_c_1252_n N_S_c_1254_n S N_S_c_1256_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%S
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%CO N_CO_M1021_d N_CO_M1008_d CO N_CO_c_1300_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%CO
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_27_115# N_A_27_115#_M1012_s
+ N_A_27_115#_M1003_d N_A_27_115#_c_1316_n N_A_27_115#_c_1319_n
+ N_A_27_115#_c_1330_n N_A_27_115#_c_1321_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_526_115# N_A_526_115#_M1020_d
+ N_A_526_115#_M1014_d N_A_526_115#_c_1338_n N_A_526_115#_c_1343_n
+ N_A_526_115#_c_1345_n N_A_526_115#_c_1346_n
+ PM_SKY130_OSU_SC_18T_HS__ADDF_L%A_526_115#
cc_1 N_GND_M1012_b N_A_M1010_g 0.0637211f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_2 N_GND_M1012_b N_A_c_288_n 0.0173144f $X=-0.045 $Y=0 $X2=2.125 $Y2=1.685
cc_3 N_GND_c_3_p N_A_c_288_n 0.0063578f $X=2.255 $Y=0.152 $X2=2.125 $Y2=1.685
cc_4 N_GND_c_4_p N_A_c_288_n 0.0043948f $X=2.34 $Y=0.825 $X2=2.125 $Y2=1.685
cc_5 N_GND_c_5_p N_A_c_288_n 0.00478641f $X=6.46 $Y=0.17 $X2=2.125 $Y2=1.685
cc_6 N_GND_M1012_b N_A_c_292_n 0.00936689f $X=-0.045 $Y=0 $X2=2.36 $Y2=1.76
cc_7 N_GND_c_4_p N_A_c_292_n 0.00243181f $X=2.34 $Y=0.825 $X2=2.36 $Y2=1.76
cc_8 N_GND_M1012_b N_A_c_294_n 0.0080793f $X=-0.045 $Y=0 $X2=2.2 $Y2=1.76
cc_9 N_GND_M1012_b N_A_c_295_n 0.00539004f $X=-0.045 $Y=0 $X2=2.36 $Y2=2.885
cc_10 N_GND_M1012_b N_A_c_296_n 0.00610054f $X=-0.045 $Y=0 $X2=2.2 $Y2=2.885
cc_11 N_GND_M1012_b N_A_c_297_n 0.0425162f $X=-0.045 $Y=0 $X2=2.435 $Y2=2.81
cc_12 N_GND_M1012_b N_A_c_298_n 0.0092911f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.885
cc_13 N_GND_M1012_b N_A_c_299_n 0.0401101f $X=-0.045 $Y=0 $X2=5.13 $Y2=2.775
cc_14 N_GND_M1012_b N_A_c_300_n 0.011447f $X=-0.045 $Y=0 $X2=5.13 $Y2=2.925
cc_15 N_GND_M1012_b N_A_c_301_n 0.0156806f $X=-0.045 $Y=0 $X2=2.35 $Y2=1.85
cc_16 N_GND_c_4_p N_A_c_301_n 3.93842e-19 $X=2.34 $Y=0.825 $X2=2.35 $Y2=1.85
cc_17 N_GND_M1012_b N_A_c_303_n 0.0035587f $X=-0.045 $Y=0 $X2=0.63 $Y2=1.85
cc_18 N_GND_M1012_b N_A_c_304_n 0.0206251f $X=-0.045 $Y=0 $X2=5.01 $Y2=1.85
cc_19 N_GND_M1012_b N_A_c_305_n 0.00106394f $X=-0.045 $Y=0 $X2=2.64 $Y2=1.85
cc_20 N_GND_M1012_b N_A_c_306_n 0.0100886f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.85
cc_21 N_GND_M1012_b N_A_c_307_n 0.0025848f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.85
cc_22 N_GND_c_4_p N_A_c_307_n 0.00283727f $X=2.34 $Y=0.825 $X2=2.495 $Y2=1.85
cc_23 N_GND_M1012_b N_A_c_309_n 0.00221228f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.85
cc_24 N_GND_M1012_b N_A_c_310_n 0.00467055f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.85
cc_25 N_GND_c_25_p N_A_c_310_n 0.00285667f $X=5.31 $Y=0.825 $X2=5.155 $Y2=1.85
cc_26 N_GND_M1012_b N_A_c_312_n 0.032623f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.85
cc_27 N_GND_M1012_b N_A_c_313_n 0.0266765f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.685
cc_28 N_GND_c_28_p N_A_c_313_n 0.00457513f $X=0.69 $Y=0.825 $X2=0.485 $Y2=1.685
cc_29 N_GND_c_29_p N_A_c_313_n 0.00640094f $X=0.605 $Y=0.152 $X2=0.485 $Y2=1.685
cc_30 N_GND_c_5_p N_A_c_313_n 0.0048006f $X=6.46 $Y=0.17 $X2=0.485 $Y2=1.685
cc_31 N_GND_M1012_b N_A_c_317_n 0.0211914f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.76
cc_32 N_GND_M1012_b N_A_c_318_n 0.0181429f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.685
cc_33 N_GND_c_4_p N_A_c_318_n 0.00434147f $X=2.34 $Y=0.825 $X2=2.495 $Y2=1.685
cc_34 N_GND_c_34_p N_A_c_318_n 0.0063578f $X=3.115 $Y=0.152 $X2=2.495 $Y2=1.685
cc_35 N_GND_c_5_p N_A_c_318_n 0.00478641f $X=6.46 $Y=0.17 $X2=2.495 $Y2=1.685
cc_36 N_GND_M1012_b N_A_c_322_n 0.0286791f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.85
cc_37 N_GND_c_25_p N_A_c_322_n 0.00140903f $X=5.31 $Y=0.825 $X2=5.155 $Y2=1.85
cc_38 N_GND_M1012_b N_A_c_324_n 0.0189719f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.685
cc_39 N_GND_c_39_p N_A_c_324_n 0.0063578f $X=5.225 $Y=0.152 $X2=5.155 $Y2=1.685
cc_40 N_GND_c_25_p N_A_c_324_n 0.00474705f $X=5.31 $Y=0.825 $X2=5.155 $Y2=1.685
cc_41 N_GND_c_5_p N_A_c_324_n 0.00478641f $X=6.46 $Y=0.17 $X2=5.155 $Y2=1.685
cc_42 N_GND_M1012_b N_B_M1003_g 0.0614047f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.075
cc_43 N_GND_c_28_p N_B_M1003_g 0.00431874f $X=0.69 $Y=0.825 $X2=0.905 $Y2=1.075
cc_44 N_GND_c_3_p N_B_M1003_g 0.0063578f $X=2.255 $Y=0.152 $X2=0.905 $Y2=1.075
cc_45 N_GND_c_5_p N_B_M1003_g 0.00478641f $X=6.46 $Y=0.17 $X2=0.905 $Y2=1.075
cc_46 N_GND_M1012_b N_B_M1025_g 0.0477186f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.075
cc_47 N_GND_c_3_p N_B_M1025_g 0.0063578f $X=2.255 $Y=0.152 $X2=1.765 $Y2=1.075
cc_48 N_GND_c_5_p N_B_M1025_g 0.00478641f $X=6.46 $Y=0.17 $X2=1.765 $Y2=1.075
cc_49 N_GND_M1012_b N_B_M1023_g 0.0177314f $X=-0.045 $Y=0 $X2=1.765 $Y2=4.585
cc_50 N_GND_M1012_b N_B_M1022_g 0.0445732f $X=-0.045 $Y=0 $X2=2.985 $Y2=4.585
cc_51 N_GND_M1012_b N_B_M1017_g 0.050864f $X=-0.045 $Y=0 $X2=4.275 $Y2=1.075
cc_52 N_GND_c_39_p N_B_M1017_g 0.00486945f $X=5.225 $Y=0.152 $X2=4.275 $Y2=1.075
cc_53 N_GND_c_5_p N_B_M1017_g 0.00478641f $X=6.46 $Y=0.17 $X2=4.275 $Y2=1.075
cc_54 N_GND_M1012_b N_B_M1016_g 0.00794292f $X=-0.045 $Y=0 $X2=4.275 $Y2=4.585
cc_55 N_GND_M1012_b N_B_c_508_n 0.00747922f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.76
cc_56 N_GND_M1012_b N_B_c_509_n 0.020418f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.76
cc_57 N_GND_M1012_b N_B_c_510_n 0.00462048f $X=-0.045 $Y=0 $X2=2.015 $Y2=2.43
cc_58 N_GND_M1012_b N_B_c_511_n 0.0408357f $X=-0.045 $Y=0 $X2=2.015 $Y2=2.43
cc_59 N_GND_M1012_b N_B_c_512_n 0.0254763f $X=-0.045 $Y=0 $X2=2.16 $Y2=2.59
cc_60 N_GND_M1012_b N_B_c_513_n 0.0127164f $X=-0.045 $Y=0 $X2=0.63 $Y2=2.59
cc_61 N_GND_M1012_b N_B_c_514_n 0.011565f $X=-0.045 $Y=0 $X2=2.83 $Y2=2.59
cc_62 N_GND_M1012_b N_B_c_515_n 0.00467059f $X=-0.045 $Y=0 $X2=2.45 $Y2=2.59
cc_63 N_GND_M1012_b N_B_c_516_n 0.00762182f $X=-0.045 $Y=0 $X2=4.06 $Y2=2.592
cc_64 N_GND_M1012_b N_B_c_517_n 0.0195197f $X=-0.045 $Y=0 $X2=3.67 $Y2=2.592
cc_65 N_GND_M1012_b N_B_c_518_n 0.00291156f $X=-0.045 $Y=0 $X2=0.485 $Y2=2.59
cc_66 N_GND_M1012_b N_B_c_519_n 0.00586424f $X=-0.045 $Y=0 $X2=2.305 $Y2=2.59
cc_67 N_GND_M1012_b N_B_c_520_n 0.00316881f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.59
cc_68 N_GND_M1012_b N_B_c_521_n 0.00792941f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.85
cc_69 N_GND_M1012_b N_B_c_522_n 0.0259978f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.85
cc_70 N_GND_M1012_b N_B_c_523_n 0.0186037f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.685
cc_71 N_GND_c_34_p N_B_c_523_n 0.0063578f $X=3.115 $Y=0.152 $X2=2.975 $Y2=1.685
cc_72 N_GND_c_72_p N_B_c_523_n 0.00431874f $X=3.2 $Y=0.825 $X2=2.975 $Y2=1.685
cc_73 N_GND_c_5_p N_B_c_523_n 0.00478641f $X=6.46 $Y=0.17 $X2=2.975 $Y2=1.685
cc_74 N_GND_M1012_b N_B_c_527_n 0.0239449f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.59
cc_75 N_GND_M1012_b N_CI_M1005_g 0.0366615f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.075
cc_76 N_GND_c_3_p N_CI_M1005_g 0.0063578f $X=2.255 $Y=0.152 $X2=1.335 $Y2=1.075
cc_77 N_GND_c_5_p N_CI_M1005_g 0.00478641f $X=6.46 $Y=0.17 $X2=1.335 $Y2=1.075
cc_78 N_GND_M1012_b N_CI_M1004_g 0.0255405f $X=-0.045 $Y=0 $X2=1.335 $Y2=4.585
cc_79 N_GND_M1012_b N_CI_M1014_g 0.0516904f $X=-0.045 $Y=0 $X2=3.415 $Y2=1.075
cc_80 N_GND_c_72_p N_CI_M1014_g 0.00431874f $X=3.2 $Y=0.825 $X2=3.415 $Y2=1.075
cc_81 N_GND_c_39_p N_CI_M1014_g 0.0063578f $X=5.225 $Y=0.152 $X2=3.415 $Y2=1.075
cc_82 N_GND_c_5_p N_CI_M1014_g 0.00478641f $X=6.46 $Y=0.17 $X2=3.415 $Y2=1.075
cc_83 N_GND_M1012_b N_CI_M1011_g 0.00805841f $X=-0.045 $Y=0 $X2=3.415 $Y2=4.585
cc_84 N_GND_M1012_b N_CI_M1009_g 0.0444321f $X=-0.045 $Y=0 $X2=4.685 $Y2=1.075
cc_85 N_GND_c_39_p N_CI_M1009_g 0.0063578f $X=5.225 $Y=0.152 $X2=4.685 $Y2=1.075
cc_86 N_GND_c_5_p N_CI_M1009_g 0.00478641f $X=6.46 $Y=0.17 $X2=4.685 $Y2=1.075
cc_87 N_GND_M1012_b N_CI_M1007_g 0.0180089f $X=-0.045 $Y=0 $X2=4.685 $Y2=4.585
cc_88 N_GND_M1012_b N_CI_c_736_n 0.00272047f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.59
cc_89 N_GND_M1012_b N_CI_c_737_n 0.0265765f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.59
cc_90 N_GND_M1012_b N_CI_c_738_n 0.015493f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.22
cc_91 N_GND_M1012_b N_CI_c_739_n 0.00162047f $X=-0.045 $Y=0 $X2=1.47 $Y2=2.22
cc_92 N_GND_M1012_b N_CI_c_740_n 0.0152192f $X=-0.045 $Y=0 $X2=4.6 $Y2=2.22
cc_93 N_GND_M1012_b N_CI_c_741_n 0.00269437f $X=-0.045 $Y=0 $X2=3.56 $Y2=2.22
cc_94 N_GND_M1012_b CI 0.0130618f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.22
cc_95 N_GND_M1012_b N_CI_c_743_n 4.344e-19 $X=-0.045 $Y=0 $X2=1.325 $Y2=2.22
cc_96 N_GND_M1012_b N_CI_c_744_n 0.00355008f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.22
cc_97 N_GND_M1012_b N_CI_c_745_n 0.00618156f $X=-0.045 $Y=0 $X2=4.745 $Y2=2.22
cc_98 N_GND_M1012_b N_CI_c_746_n 0.00482822f $X=-0.045 $Y=0 $X2=4.745 $Y2=2.22
cc_99 N_GND_M1012_b N_CI_c_747_n 0.0263369f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.22
cc_100 N_GND_M1012_b N_CI_c_748_n 0.027099f $X=-0.045 $Y=0 $X2=4.745 $Y2=2.4
cc_101 N_GND_M1012_b N_CON_c_906_n 0.0180088f $X=-0.045 $Y=0 $X2=3.845 $Y2=1.685
cc_102 N_GND_c_39_p N_CON_c_906_n 0.0063578f $X=5.225 $Y=0.152 $X2=3.845
+ $Y2=1.685
cc_103 N_GND_c_5_p N_CON_c_906_n 0.00478641f $X=6.46 $Y=0.17 $X2=3.845 $Y2=1.685
cc_104 N_GND_M1012_b N_CON_M1013_g 0.0372583f $X=-0.045 $Y=0 $X2=3.845 $Y2=4.585
cc_105 N_GND_M1012_b N_CON_M1021_g 0.107867f $X=-0.045 $Y=0 $X2=6.535 $Y2=0.945
cc_106 N_GND_c_106_p N_CON_M1021_g 0.00887945f $X=6.32 $Y=0.825 $X2=6.535
+ $Y2=0.945
cc_107 N_GND_c_5_p N_CON_M1021_g 0.00481485f $X=6.46 $Y=0.17 $X2=6.535 $Y2=0.945
cc_108 N_GND_M1012_b N_CON_c_913_n 0.00911049f $X=-0.045 $Y=0 $X2=1.665
+ $Y2=3.025
cc_109 N_GND_M1012_b N_CON_c_914_n 0.0107538f $X=-0.045 $Y=0 $X2=6.41 $Y2=2.74
cc_110 N_GND_M1012_b N_CON_c_915_n 0.0356508f $X=-0.045 $Y=0 $X2=6.41 $Y2=2.74
cc_111 N_GND_M1012_b N_CON_c_916_n 0.00462698f $X=-0.045 $Y=0 $X2=1.665
+ $Y2=1.765
cc_112 N_GND_M1012_b N_CON_c_917_n 0.0252944f $X=-0.045 $Y=0 $X2=3.845 $Y2=1.85
cc_113 N_GND_M1012_b N_CON_c_918_n 0.00293622f $X=-0.045 $Y=0 $X2=3.97 $Y2=1.85
cc_114 N_GND_M1027_d N_CON_c_919_n 0.00601493f $X=2.2 $Y=0.575 $X2=3.825
+ $Y2=1.48
cc_115 N_GND_M1024_d N_CON_c_919_n 0.00243973f $X=3.06 $Y=0.575 $X2=3.825
+ $Y2=1.48
cc_116 N_GND_c_4_p N_CON_c_919_n 0.0130682f $X=2.34 $Y=0.825 $X2=3.825 $Y2=1.48
cc_117 N_GND_c_72_p N_CON_c_919_n 0.00105102f $X=3.2 $Y=0.825 $X2=3.825 $Y2=1.48
cc_118 N_GND_M1012_b N_CON_c_923_n 5.54826e-19 $X=-0.045 $Y=0 $X2=1.695 $Y2=1.48
cc_119 N_GND_c_4_p N_CON_c_923_n 5.67165e-19 $X=2.34 $Y=0.825 $X2=1.695 $Y2=1.48
cc_120 N_GND_M1006_d N_CON_c_925_n 0.00891659f $X=5.17 $Y=0.575 $X2=5.995
+ $Y2=1.48
cc_121 N_GND_M1012_b N_CON_c_925_n 0.0146888f $X=-0.045 $Y=0 $X2=5.995 $Y2=1.48
cc_122 N_GND_c_25_p N_CON_c_925_n 0.0133019f $X=5.31 $Y=0.825 $X2=5.995 $Y2=1.48
cc_123 N_GND_M1012_b N_CON_c_928_n 4.50048e-19 $X=-0.045 $Y=0 $X2=4.115 $Y2=1.48
cc_124 N_GND_M1012_b N_CON_c_929_n 0.00107881f $X=-0.045 $Y=0 $X2=3.97 $Y2=1.48
cc_125 N_GND_M1012_b CON 0.0206838f $X=-0.045 $Y=0 $X2=6.14 $Y2=1.48
cc_126 N_GND_c_106_p CON 0.00133737f $X=6.32 $Y=0.825 $X2=6.14 $Y2=1.48
cc_127 N_GND_M1012_b N_CON_c_932_n 0.00417041f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_128 N_GND_c_3_p N_CON_c_932_n 0.00779312f $X=2.255 $Y=0.152 $X2=1.55
+ $Y2=0.825
cc_129 N_GND_c_4_p N_CON_c_932_n 4.05842e-19 $X=2.34 $Y=0.825 $X2=1.55 $Y2=0.825
cc_130 N_GND_c_5_p N_CON_c_932_n 0.00478039f $X=6.46 $Y=0.17 $X2=1.55 $Y2=0.825
cc_131 N_GND_M1012_b N_CON_c_936_n 0.0126281f $X=-0.045 $Y=0 $X2=6.41 $Y2=1.48
cc_132 N_GND_c_106_p N_CON_c_936_n 0.00804004f $X=6.32 $Y=0.825 $X2=6.41
+ $Y2=1.48
cc_133 N_GND_M1012_b N_A_784_115#_M1018_g 0.0885152f $X=-0.045 $Y=0 $X2=5.585
+ $Y2=0.945
cc_134 N_GND_c_25_p N_A_784_115#_M1018_g 0.0114373f $X=5.31 $Y=0.825 $X2=5.585
+ $Y2=0.945
cc_135 N_GND_c_135_p N_A_784_115#_M1018_g 0.00644441f $X=6.235 $Y=0.152
+ $X2=5.585 $Y2=0.945
cc_136 N_GND_c_106_p N_A_784_115#_M1018_g 0.00495414f $X=6.32 $Y=0.825 $X2=5.585
+ $Y2=0.945
cc_137 N_GND_c_5_p N_A_784_115#_M1018_g 0.00481485f $X=6.46 $Y=0.17 $X2=5.585
+ $Y2=0.945
cc_138 N_GND_M1012_b N_A_784_115#_c_1096_n 0.00887593f $X=-0.045 $Y=0 $X2=3.845
+ $Y2=3.03
cc_139 N_GND_M1012_b N_A_784_115#_c_1097_n 0.00593307f $X=-0.045 $Y=0 $X2=4.225
+ $Y2=2.22
cc_140 N_GND_M1012_b N_A_784_115#_c_1098_n 9.19767e-19 $X=-0.045 $Y=0 $X2=3.93
+ $Y2=2.22
cc_141 N_GND_M1012_b N_A_784_115#_c_1099_n 0.00156608f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=0.905
cc_142 N_GND_c_39_p N_A_784_115#_c_1099_n 0.00756162f $X=5.225 $Y=0.152 $X2=4.06
+ $Y2=0.905
cc_143 N_GND_c_5_p N_A_784_115#_c_1099_n 0.00467629f $X=6.46 $Y=0.17 $X2=4.06
+ $Y2=0.905
cc_144 N_GND_M1012_b N_A_784_115#_c_1102_n 0.00483243f $X=-0.045 $Y=0 $X2=4.31
+ $Y2=2.135
cc_145 N_GND_c_39_p N_A_784_115#_c_1103_n 0.0029768f $X=5.225 $Y=0.152 $X2=4.31
+ $Y2=0.99
cc_146 N_GND_c_5_p N_A_784_115#_c_1103_n 0.00530192f $X=6.46 $Y=0.17 $X2=4.31
+ $Y2=0.99
cc_147 N_GND_M1012_b N_A_784_115#_c_1105_n 0.00798748f $X=-0.045 $Y=0 $X2=5.415
+ $Y2=2.755
cc_148 N_GND_M1012_b N_A_784_115#_c_1106_n 0.0268831f $X=-0.045 $Y=0 $X2=5.585
+ $Y2=2.755
cc_149 N_GND_M1012_b N_S_c_1246_n 0.0215204f $X=-0.045 $Y=0 $X2=5.8 $Y2=0.825
cc_150 N_GND_c_25_p N_S_c_1246_n 0.0212016f $X=5.31 $Y=0.825 $X2=5.8 $Y2=0.825
cc_151 N_GND_c_135_p N_S_c_1246_n 0.00736239f $X=6.235 $Y=0.152 $X2=5.8
+ $Y2=0.825
cc_152 N_GND_c_106_p N_S_c_1246_n 0.0213592f $X=6.32 $Y=0.825 $X2=5.8 $Y2=0.825
cc_153 N_GND_c_5_p N_S_c_1246_n 0.00476261f $X=6.46 $Y=0.17 $X2=5.8 $Y2=0.825
cc_154 N_GND_M1012_b N_S_c_1251_n 0.0135159f $X=-0.045 $Y=0 $X2=5.925 $Y2=3.165
cc_155 N_GND_M1012_b N_S_c_1252_n 0.0121999f $X=-0.045 $Y=0 $X2=5.925 $Y2=2.22
cc_156 N_GND_M1012_b CO 0.00667411f $X=-0.045 $Y=0 $X2=6.75 $Y2=2.96
cc_157 N_GND_M1012_b N_CO_c_1300_n 0.080877f $X=-0.045 $Y=0 $X2=6.75 $Y2=0.825
cc_158 N_GND_c_5_p N_CO_c_1300_n 0.00476261f $X=6.46 $Y=0.17 $X2=6.75 $Y2=0.825
cc_159 N_GND_M1012_b N_A_27_115#_c_1316_n 0.00156053f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_160 N_GND_c_29_p N_A_27_115#_c_1316_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_161 N_GND_c_5_p N_A_27_115#_c_1316_n 0.00476261f $X=6.46 $Y=0.17 $X2=0.26
+ $Y2=0.825
cc_162 N_GND_M1012_d N_A_27_115#_c_1319_n 0.00427893f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.345
cc_163 N_GND_c_28_p N_A_27_115#_c_1319_n 0.0126786f $X=0.69 $Y=0.825 $X2=1.035
+ $Y2=1.345
cc_164 N_GND_M1012_b N_A_27_115#_c_1321_n 0.00158615f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.825
cc_165 N_GND_c_28_p N_A_27_115#_c_1321_n 2.23682e-19 $X=0.69 $Y=0.825 $X2=1.12
+ $Y2=0.825
cc_166 N_GND_c_3_p N_A_27_115#_c_1321_n 0.00775613f $X=2.255 $Y=0.152 $X2=1.12
+ $Y2=0.825
cc_167 N_GND_c_5_p N_A_27_115#_c_1321_n 0.00478039f $X=6.46 $Y=0.17 $X2=1.12
+ $Y2=0.825
cc_168 N_GND_M1012_b N_A_526_115#_c_1338_n 0.00158615f $X=-0.045 $Y=0 $X2=2.77
+ $Y2=0.825
cc_169 N_GND_c_4_p N_A_526_115#_c_1338_n 2.23682e-19 $X=2.34 $Y=0.825 $X2=2.77
+ $Y2=0.825
cc_170 N_GND_c_34_p N_A_526_115#_c_1338_n 0.00797044f $X=3.115 $Y=0.152 $X2=2.77
+ $Y2=0.825
cc_171 N_GND_c_72_p N_A_526_115#_c_1338_n 2.23682e-19 $X=3.2 $Y=0.825 $X2=2.77
+ $Y2=0.825
cc_172 N_GND_c_5_p N_A_526_115#_c_1338_n 0.00478039f $X=6.46 $Y=0.17 $X2=2.77
+ $Y2=0.825
cc_173 N_GND_M1024_d N_A_526_115#_c_1343_n 0.00465706f $X=3.06 $Y=0.575
+ $X2=3.545 $Y2=1.345
cc_174 N_GND_c_72_p N_A_526_115#_c_1343_n 0.0116202f $X=3.2 $Y=0.825 $X2=3.545
+ $Y2=1.345
cc_175 N_GND_c_4_p N_A_526_115#_c_1345_n 4.77496e-19 $X=2.34 $Y=0.825 $X2=2.855
+ $Y2=1.345
cc_176 N_GND_M1012_b N_A_526_115#_c_1346_n 0.00158615f $X=-0.045 $Y=0 $X2=3.63
+ $Y2=0.825
cc_177 N_GND_c_72_p N_A_526_115#_c_1346_n 2.23682e-19 $X=3.2 $Y=0.825 $X2=3.63
+ $Y2=0.825
cc_178 N_GND_c_39_p N_A_526_115#_c_1346_n 0.00775613f $X=5.225 $Y=0.152 $X2=3.63
+ $Y2=0.825
cc_179 N_GND_c_5_p N_A_526_115#_c_1346_n 0.00478039f $X=6.46 $Y=0.17 $X2=3.63
+ $Y2=0.825
cc_180 N_VDD_M1010_b N_A_M1010_g 0.0292364f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_181 N_VDD_c_181_p N_A_M1010_g 0.00354579f $X=0.69 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_182 N_VDD_c_182_p N_A_M1010_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_183 N_VDD_c_183_p N_A_M1010_g 0.00468827f $X=6.46 $Y=6.49 $X2=0.475 $Y2=4.585
cc_184 N_VDD_M1010_b N_A_c_332_n 0.0164334f $X=-0.045 $Y=2.905 $X2=2.125
+ $Y2=2.96
cc_185 N_VDD_c_185_p N_A_c_332_n 0.00606474f $X=2.255 $Y=6.507 $X2=2.125
+ $Y2=2.96
cc_186 N_VDD_c_186_p N_A_c_332_n 0.00354579f $X=2.34 $Y=3.795 $X2=2.125 $Y2=2.96
cc_187 N_VDD_c_183_p N_A_c_332_n 0.00468827f $X=6.46 $Y=6.49 $X2=2.125 $Y2=2.96
cc_188 N_VDD_M1010_b N_A_c_295_n 0.00298392f $X=-0.045 $Y=2.905 $X2=2.36
+ $Y2=2.885
cc_189 N_VDD_c_186_p N_A_c_295_n 0.00280084f $X=2.34 $Y=3.795 $X2=2.36 $Y2=2.885
cc_190 N_VDD_M1010_b N_A_c_296_n 0.00180595f $X=-0.045 $Y=2.905 $X2=2.2
+ $Y2=2.885
cc_191 N_VDD_M1010_b N_A_c_339_n 0.0171656f $X=-0.045 $Y=2.905 $X2=2.555
+ $Y2=2.96
cc_192 N_VDD_c_186_p N_A_c_339_n 0.00354579f $X=2.34 $Y=3.795 $X2=2.555 $Y2=2.96
cc_193 N_VDD_c_193_p N_A_c_339_n 0.00606474f $X=3.115 $Y=6.507 $X2=2.555
+ $Y2=2.96
cc_194 N_VDD_c_183_p N_A_c_339_n 0.00468827f $X=6.46 $Y=6.49 $X2=2.555 $Y2=2.96
cc_195 N_VDD_M1010_b N_A_M1002_g 0.0203606f $X=-0.045 $Y=2.905 $X2=5.095
+ $Y2=4.585
cc_196 N_VDD_c_196_p N_A_M1002_g 0.0061469f $X=5.225 $Y=6.507 $X2=5.095
+ $Y2=4.585
cc_197 N_VDD_c_197_p N_A_M1002_g 0.0039779f $X=5.31 $Y=4.135 $X2=5.095 $Y2=4.585
cc_198 N_VDD_c_183_p N_A_M1002_g 0.00471609f $X=6.46 $Y=6.49 $X2=5.095 $Y2=4.585
cc_199 N_VDD_M1010_b N_A_c_298_n 0.00372423f $X=-0.045 $Y=2.905 $X2=2.555
+ $Y2=2.885
cc_200 N_VDD_M1010_b N_A_c_300_n 0.0032155f $X=-0.045 $Y=2.905 $X2=5.13
+ $Y2=2.925
cc_201 N_VDD_M1010_b N_B_M1000_g 0.0194747f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_202 N_VDD_c_181_p N_B_M1000_g 0.00354579f $X=0.69 $Y=4.135 $X2=0.905
+ $Y2=4.585
cc_203 N_VDD_c_185_p N_B_M1000_g 0.00606474f $X=2.255 $Y=6.507 $X2=0.905
+ $Y2=4.585
cc_204 N_VDD_c_183_p N_B_M1000_g 0.00468827f $X=6.46 $Y=6.49 $X2=0.905 $Y2=4.585
cc_205 N_VDD_M1010_b N_B_M1023_g 0.0193281f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=4.585
cc_206 N_VDD_c_185_p N_B_M1023_g 0.0061469f $X=2.255 $Y=6.507 $X2=1.765
+ $Y2=4.585
cc_207 N_VDD_c_186_p N_B_M1023_g 0.00460842f $X=2.34 $Y=3.795 $X2=1.765
+ $Y2=4.585
cc_208 N_VDD_c_183_p N_B_M1023_g 0.00471609f $X=6.46 $Y=6.49 $X2=1.765 $Y2=4.585
cc_209 N_VDD_M1010_b N_B_M1022_g 0.0212396f $X=-0.045 $Y=2.905 $X2=2.985
+ $Y2=4.585
cc_210 N_VDD_c_186_p N_B_M1022_g 4.9048e-19 $X=2.34 $Y=3.795 $X2=2.985 $Y2=4.585
cc_211 N_VDD_c_193_p N_B_M1022_g 0.0061469f $X=3.115 $Y=6.507 $X2=2.985
+ $Y2=4.585
cc_212 N_VDD_c_212_p N_B_M1022_g 0.00378444f $X=3.2 $Y=4.135 $X2=2.985 $Y2=4.585
cc_213 N_VDD_c_183_p N_B_M1022_g 0.00471609f $X=6.46 $Y=6.49 $X2=2.985 $Y2=4.585
cc_214 N_VDD_M1010_b N_B_M1016_g 0.0209183f $X=-0.045 $Y=2.905 $X2=4.275
+ $Y2=4.585
cc_215 N_VDD_c_196_p N_B_M1016_g 0.0061469f $X=5.225 $Y=6.507 $X2=4.275
+ $Y2=4.585
cc_216 N_VDD_c_183_p N_B_M1016_g 0.00471609f $X=6.46 $Y=6.49 $X2=4.275 $Y2=4.585
cc_217 N_VDD_M1010_b N_B_c_509_n 0.00479818f $X=-0.045 $Y=2.905 $X2=0.895
+ $Y2=2.76
cc_218 N_VDD_M1010_b N_CI_M1004_g 0.0211777f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=4.585
cc_219 N_VDD_c_181_p N_CI_M1004_g 4.9048e-19 $X=0.69 $Y=4.135 $X2=1.335
+ $Y2=4.585
cc_220 N_VDD_c_185_p N_CI_M1004_g 0.0061469f $X=2.255 $Y=6.507 $X2=1.335
+ $Y2=4.585
cc_221 N_VDD_c_183_p N_CI_M1004_g 0.00471609f $X=6.46 $Y=6.49 $X2=1.335
+ $Y2=4.585
cc_222 N_VDD_M1010_b N_CI_M1011_g 0.0211273f $X=-0.045 $Y=2.905 $X2=3.415
+ $Y2=4.585
cc_223 N_VDD_c_212_p N_CI_M1011_g 0.00378444f $X=3.2 $Y=4.135 $X2=3.415
+ $Y2=4.585
cc_224 N_VDD_c_196_p N_CI_M1011_g 0.0061469f $X=5.225 $Y=6.507 $X2=3.415
+ $Y2=4.585
cc_225 N_VDD_c_183_p N_CI_M1011_g 0.00471609f $X=6.46 $Y=6.49 $X2=3.415
+ $Y2=4.585
cc_226 N_VDD_M1010_b N_CI_M1007_g 0.0206974f $X=-0.045 $Y=2.905 $X2=4.685
+ $Y2=4.585
cc_227 N_VDD_c_196_p N_CI_M1007_g 0.0061469f $X=5.225 $Y=6.507 $X2=4.685
+ $Y2=4.585
cc_228 N_VDD_c_183_p N_CI_M1007_g 0.00471609f $X=6.46 $Y=6.49 $X2=4.685
+ $Y2=4.585
cc_229 N_VDD_M1010_b N_CON_M1013_g 0.01904f $X=-0.045 $Y=2.905 $X2=3.845
+ $Y2=4.585
cc_230 N_VDD_c_196_p N_CON_M1013_g 0.0061469f $X=5.225 $Y=6.507 $X2=3.845
+ $Y2=4.585
cc_231 N_VDD_c_183_p N_CON_M1013_g 0.00471609f $X=6.46 $Y=6.49 $X2=3.845
+ $Y2=4.585
cc_232 N_VDD_M1010_b N_CON_M1008_g 0.0955179f $X=-0.045 $Y=2.905 $X2=6.535
+ $Y2=5.085
cc_233 N_VDD_c_233_p N_CON_M1008_g 0.00809569f $X=6.32 $Y=4.46 $X2=6.535
+ $Y2=5.085
cc_234 N_VDD_c_183_p N_CON_M1008_g 0.00471609f $X=6.46 $Y=6.49 $X2=6.535
+ $Y2=5.085
cc_235 N_VDD_c_235_p N_CON_M1008_g 0.0061469f $X=6.46 $Y=6.44 $X2=6.535
+ $Y2=5.085
cc_236 N_VDD_M1010_b N_CON_c_945_n 0.00155118f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=3.795
cc_237 N_VDD_c_185_p N_CON_c_945_n 0.00737727f $X=2.255 $Y=6.507 $X2=1.55
+ $Y2=3.795
cc_238 N_VDD_c_183_p N_CON_c_945_n 0.00475776f $X=6.46 $Y=6.49 $X2=1.55
+ $Y2=3.795
cc_239 N_VDD_M1010_b N_CON_c_913_n 0.00397971f $X=-0.045 $Y=2.905 $X2=1.665
+ $Y2=3.025
cc_240 N_VDD_M1010_b N_CON_c_914_n 0.00545748f $X=-0.045 $Y=2.905 $X2=6.41
+ $Y2=2.74
cc_241 N_VDD_M1010_b N_CON_c_915_n 0.00643378f $X=-0.045 $Y=2.905 $X2=6.41
+ $Y2=2.74
cc_242 N_VDD_M1010_b N_A_784_115#_M1001_g 0.0840054f $X=-0.045 $Y=2.905
+ $X2=5.585 $Y2=5.085
cc_243 N_VDD_c_197_p N_A_784_115#_M1001_g 0.0224174f $X=5.31 $Y=4.135 $X2=5.585
+ $Y2=5.085
cc_244 N_VDD_c_244_p N_A_784_115#_M1001_g 0.0061469f $X=6.235 $Y=6.507 $X2=5.585
+ $Y2=5.085
cc_245 N_VDD_c_233_p N_A_784_115#_M1001_g 0.00701284f $X=6.32 $Y=4.46 $X2=5.585
+ $Y2=5.085
cc_246 N_VDD_c_183_p N_A_784_115#_M1001_g 0.00471609f $X=6.46 $Y=6.49 $X2=5.585
+ $Y2=5.085
cc_247 N_VDD_M1010_b N_A_784_115#_c_1096_n 0.00257504f $X=-0.045 $Y=2.905
+ $X2=3.845 $Y2=3.03
cc_248 N_VDD_M1010_b N_A_784_115#_c_1113_n 0.00427075f $X=-0.045 $Y=2.905
+ $X2=4.06 $Y2=3.42
cc_249 N_VDD_M1010_b N_A_784_115#_c_1114_n 0.00155118f $X=-0.045 $Y=2.905
+ $X2=4.06 $Y2=3.795
cc_250 N_VDD_c_196_p N_A_784_115#_c_1114_n 0.0075556f $X=5.225 $Y=6.507 $X2=4.06
+ $Y2=3.795
cc_251 N_VDD_c_183_p N_A_784_115#_c_1114_n 0.00475776f $X=6.46 $Y=6.49 $X2=4.06
+ $Y2=3.795
cc_252 N_VDD_M1002_d N_A_784_115#_c_1117_n 0.00913117f $X=5.17 $Y=3.085 $X2=5.33
+ $Y2=3.335
cc_253 N_VDD_M1010_b N_A_784_115#_c_1117_n 0.00388557f $X=-0.045 $Y=2.905
+ $X2=5.33 $Y2=3.335
cc_254 N_VDD_c_197_p N_A_784_115#_c_1117_n 0.00666443f $X=5.31 $Y=4.135 $X2=5.33
+ $Y2=3.335
cc_255 N_VDD_M1002_d N_A_784_115#_c_1120_n 0.00259083f $X=5.17 $Y=3.085
+ $X2=5.415 $Y2=3.25
cc_256 N_VDD_M1010_b N_A_784_115#_c_1120_n 0.00416996f $X=-0.045 $Y=2.905
+ $X2=5.415 $Y2=3.25
cc_257 N_VDD_M1010_b N_A_784_115#_c_1105_n 6.65464e-19 $X=-0.045 $Y=2.905
+ $X2=5.415 $Y2=2.755
cc_258 N_VDD_M1010_b N_A_784_115#_c_1106_n 0.00469272f $X=-0.045 $Y=2.905
+ $X2=5.585 $Y2=2.755
cc_259 N_VDD_M1010_b N_A_27_617#_c_1219_n 0.00156053f $X=-0.045 $Y=2.905
+ $X2=0.26 $Y2=3.795
cc_260 N_VDD_c_182_p N_A_27_617#_c_1219_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=3.795
cc_261 N_VDD_c_183_p N_A_27_617#_c_1219_n 0.00476261f $X=6.46 $Y=6.49 $X2=0.26
+ $Y2=3.795
cc_262 N_VDD_M1010_d N_A_27_617#_c_1222_n 0.00549367f $X=0.55 $Y=3.085 $X2=1.035
+ $Y2=3.46
cc_263 N_VDD_c_181_p N_A_27_617#_c_1222_n 0.00809661f $X=0.69 $Y=4.135 $X2=1.035
+ $Y2=3.46
cc_264 N_VDD_M1010_b N_A_27_617#_c_1224_n 0.00155118f $X=-0.045 $Y=2.905
+ $X2=1.12 $Y2=3.795
cc_265 N_VDD_c_185_p N_A_27_617#_c_1224_n 0.00734006f $X=2.255 $Y=6.507 $X2=1.12
+ $Y2=3.795
cc_266 N_VDD_c_183_p N_A_27_617#_c_1224_n 0.00475776f $X=6.46 $Y=6.49 $X2=1.12
+ $Y2=3.795
cc_267 N_VDD_M1010_b N_A_526_617#_c_1232_n 0.00155118f $X=-0.045 $Y=2.905
+ $X2=2.77 $Y2=3.795
cc_268 N_VDD_c_193_p N_A_526_617#_c_1232_n 0.0075556f $X=3.115 $Y=6.507 $X2=2.77
+ $Y2=3.795
cc_269 N_VDD_c_183_p N_A_526_617#_c_1232_n 0.00475776f $X=6.46 $Y=6.49 $X2=2.77
+ $Y2=3.795
cc_270 N_VDD_M1022_d N_A_526_617#_c_1235_n 0.00868143f $X=3.06 $Y=3.085
+ $X2=3.545 $Y2=3.455
cc_271 N_VDD_c_212_p N_A_526_617#_c_1235_n 0.00800981f $X=3.2 $Y=4.135 $X2=3.545
+ $Y2=3.455
cc_272 N_VDD_M1010_b N_A_526_617#_c_1237_n 0.00155118f $X=-0.045 $Y=2.905
+ $X2=3.63 $Y2=3.795
cc_273 N_VDD_c_196_p N_A_526_617#_c_1237_n 0.00734006f $X=5.225 $Y=6.507
+ $X2=3.63 $Y2=3.795
cc_274 N_VDD_c_183_p N_A_526_617#_c_1237_n 0.00475776f $X=6.46 $Y=6.49 $X2=3.63
+ $Y2=3.795
cc_275 N_VDD_M1010_b N_S_c_1251_n 0.00671597f $X=-0.045 $Y=2.905 $X2=5.925
+ $Y2=3.165
cc_276 N_VDD_M1010_b N_S_c_1254_n 0.0123513f $X=-0.045 $Y=2.905 $X2=5.925
+ $Y2=3.25
cc_277 N_VDD_M1010_b S 0.00760382f $X=-0.045 $Y=2.905 $X2=5.8 $Y2=3.365
cc_278 N_VDD_M1010_b N_S_c_1256_n 0.0225911f $X=-0.045 $Y=2.905 $X2=5.8
+ $Y2=3.365
cc_279 N_VDD_c_197_p N_S_c_1256_n 0.0549735f $X=5.31 $Y=4.135 $X2=5.8 $Y2=3.365
cc_280 N_VDD_c_244_p N_S_c_1256_n 0.00736239f $X=6.235 $Y=6.507 $X2=5.8
+ $Y2=3.365
cc_281 N_VDD_c_233_p N_S_c_1256_n 0.0807378f $X=6.32 $Y=4.46 $X2=5.8 $Y2=3.365
cc_282 N_VDD_c_183_p N_S_c_1256_n 0.00476261f $X=6.46 $Y=6.49 $X2=5.8 $Y2=3.365
cc_283 N_VDD_M1010_b CO 0.0109934f $X=-0.045 $Y=2.905 $X2=6.75 $Y2=2.96
cc_284 N_VDD_M1010_b N_CO_c_1300_n 0.056519f $X=-0.045 $Y=2.905 $X2=6.75
+ $Y2=0.825
cc_285 N_VDD_c_183_p N_CO_c_1300_n 0.00476261f $X=6.46 $Y=6.49 $X2=6.75
+ $Y2=0.825
cc_286 N_VDD_c_235_p N_CO_c_1300_n 0.00757793f $X=6.46 $Y=6.44 $X2=6.75
+ $Y2=0.825
cc_287 N_A_M1010_g N_B_M1003_g 0.0285181f $X=0.475 $Y=4.585 $X2=0.905 $Y2=1.075
cc_288 N_A_c_301_n N_B_M1003_g 0.00620979f $X=2.35 $Y=1.85 $X2=0.905 $Y2=1.075
cc_289 N_A_c_303_n N_B_M1003_g 8.6716e-19 $X=0.63 $Y=1.85 $X2=0.905 $Y2=1.075
cc_290 N_A_c_306_n N_B_M1003_g 0.00278747f $X=0.485 $Y=1.85 $X2=0.905 $Y2=1.075
cc_291 N_A_c_312_n N_B_M1003_g 0.0223074f $X=0.485 $Y=1.85 $X2=0.905 $Y2=1.075
cc_292 N_A_c_313_n N_B_M1003_g 0.03796f $X=0.485 $Y=1.685 $X2=0.905 $Y2=1.075
cc_293 N_A_M1010_g N_B_M1000_g 0.0531399f $X=0.475 $Y=4.585 $X2=0.905 $Y2=4.585
cc_294 N_A_c_288_n N_B_M1025_g 0.0874539f $X=2.125 $Y=1.685 $X2=1.765 $Y2=1.075
cc_295 N_A_c_301_n N_B_M1025_g 0.0037004f $X=2.35 $Y=1.85 $X2=1.765 $Y2=1.075
cc_296 N_A_c_305_n N_B_M1025_g 5.04344e-19 $X=2.64 $Y=1.85 $X2=1.765 $Y2=1.075
cc_297 N_A_c_307_n N_B_M1025_g 0.00113262f $X=2.495 $Y=1.85 $X2=1.765 $Y2=1.075
cc_298 N_A_c_317_n N_B_M1025_g 0.00810048f $X=2.495 $Y=1.76 $X2=1.765 $Y2=1.075
cc_299 N_A_c_296_n N_B_M1023_g 0.202045f $X=2.2 $Y=2.885 $X2=1.765 $Y2=4.585
cc_300 N_A_c_297_n N_B_M1023_g 0.00269561f $X=2.435 $Y=2.81 $X2=1.765 $Y2=4.585
cc_301 N_A_c_297_n N_B_M1022_g 0.0237419f $X=2.435 $Y=2.81 $X2=2.985 $Y2=4.585
cc_302 N_A_c_298_n N_B_M1022_g 0.0455598f $X=2.555 $Y=2.885 $X2=2.985 $Y2=4.585
cc_303 N_A_c_304_n N_B_M1017_g 0.00127853f $X=5.01 $Y=1.85 $X2=4.275 $Y2=1.075
cc_304 N_A_M1010_g N_B_c_508_n 4.31631e-19 $X=0.475 $Y=4.585 $X2=0.895 $Y2=2.76
cc_305 N_A_c_312_n N_B_c_508_n 8.97793e-19 $X=0.485 $Y=1.85 $X2=0.895 $Y2=2.76
cc_306 N_A_M1010_g N_B_c_509_n 0.0218907f $X=0.475 $Y=4.585 $X2=0.895 $Y2=2.76
cc_307 N_A_c_294_n N_B_c_510_n 4.19356e-19 $X=2.2 $Y=1.76 $X2=2.015 $Y2=2.43
cc_308 N_A_c_296_n N_B_c_510_n 9.92874e-19 $X=2.2 $Y=2.885 $X2=2.015 $Y2=2.43
cc_309 N_A_c_297_n N_B_c_510_n 0.00170298f $X=2.435 $Y=2.81 $X2=2.015 $Y2=2.43
cc_310 N_A_c_301_n N_B_c_510_n 0.00231345f $X=2.35 $Y=1.85 $X2=2.015 $Y2=2.43
cc_311 N_A_c_294_n N_B_c_511_n 0.00301833f $X=2.2 $Y=1.76 $X2=2.015 $Y2=2.43
cc_312 N_A_c_296_n N_B_c_511_n 0.00640881f $X=2.2 $Y=2.885 $X2=2.015 $Y2=2.43
cc_313 N_A_c_297_n N_B_c_511_n 0.022133f $X=2.435 $Y=2.81 $X2=2.015 $Y2=2.43
cc_314 N_A_c_301_n N_B_c_511_n 5.24163e-19 $X=2.35 $Y=1.85 $X2=2.015 $Y2=2.43
cc_315 N_A_c_296_n N_B_c_512_n 0.00100445f $X=2.2 $Y=2.885 $X2=2.16 $Y2=2.59
cc_316 N_A_M1010_g N_B_c_513_n 0.00322062f $X=0.475 $Y=4.585 $X2=0.63 $Y2=2.59
cc_317 N_A_c_303_n N_B_c_513_n 0.003172f $X=0.63 $Y=1.85 $X2=0.63 $Y2=2.59
cc_318 N_A_c_306_n N_B_c_513_n 9.8095e-19 $X=0.485 $Y=1.85 $X2=0.63 $Y2=2.59
cc_319 N_A_c_312_n N_B_c_513_n 7.14347e-19 $X=0.485 $Y=1.85 $X2=0.63 $Y2=2.59
cc_320 N_A_c_297_n N_B_c_514_n 0.00451179f $X=2.435 $Y=2.81 $X2=2.83 $Y2=2.59
cc_321 N_A_c_298_n N_B_c_514_n 0.00349205f $X=2.555 $Y=2.885 $X2=2.83 $Y2=2.59
cc_322 N_A_c_296_n N_B_c_515_n 0.00563612f $X=2.2 $Y=2.885 $X2=2.45 $Y2=2.59
cc_323 N_A_c_297_n N_B_c_515_n 0.0049099f $X=2.435 $Y=2.81 $X2=2.45 $Y2=2.59
cc_324 N_A_c_297_n N_B_c_517_n 3.06713e-19 $X=2.435 $Y=2.81 $X2=3.67 $Y2=2.592
cc_325 N_A_M1010_g N_B_c_518_n 0.0206591f $X=0.475 $Y=4.585 $X2=0.485 $Y2=2.59
cc_326 N_A_c_306_n N_B_c_518_n 0.00208589f $X=0.485 $Y=1.85 $X2=0.485 $Y2=2.59
cc_327 N_A_c_312_n N_B_c_518_n 3.21671e-19 $X=0.485 $Y=1.85 $X2=0.485 $Y2=2.59
cc_328 N_A_c_294_n N_B_c_519_n 0.00243929f $X=2.2 $Y=1.76 $X2=2.305 $Y2=2.59
cc_329 N_A_c_296_n N_B_c_519_n 0.00867832f $X=2.2 $Y=2.885 $X2=2.305 $Y2=2.59
cc_330 N_A_c_297_n N_B_c_519_n 0.00530786f $X=2.435 $Y=2.81 $X2=2.305 $Y2=2.59
cc_331 N_A_c_307_n N_B_c_519_n 9.1275e-19 $X=2.495 $Y=1.85 $X2=2.305 $Y2=2.59
cc_332 N_A_c_297_n N_B_c_521_n 0.00846275f $X=2.435 $Y=2.81 $X2=2.975 $Y2=1.85
cc_333 N_A_c_304_n N_B_c_521_n 0.0130411f $X=5.01 $Y=1.85 $X2=2.975 $Y2=1.85
cc_334 N_A_c_305_n N_B_c_521_n 0.00248328f $X=2.64 $Y=1.85 $X2=2.975 $Y2=1.85
cc_335 N_A_c_307_n N_B_c_521_n 0.00843011f $X=2.495 $Y=1.85 $X2=2.975 $Y2=1.85
cc_336 N_A_c_317_n N_B_c_521_n 0.00129442f $X=2.495 $Y=1.76 $X2=2.975 $Y2=1.85
cc_337 N_A_c_304_n N_B_c_522_n 0.00261058f $X=5.01 $Y=1.85 $X2=2.975 $Y2=1.85
cc_338 N_A_c_305_n N_B_c_522_n 8.85796e-19 $X=2.64 $Y=1.85 $X2=2.975 $Y2=1.85
cc_339 N_A_c_307_n N_B_c_522_n 7.65216e-19 $X=2.495 $Y=1.85 $X2=2.975 $Y2=1.85
cc_340 N_A_c_317_n N_B_c_522_n 0.0225603f $X=2.495 $Y=1.76 $X2=2.975 $Y2=1.85
cc_341 N_A_c_318_n N_B_c_523_n 0.0247128f $X=2.495 $Y=1.685 $X2=2.975 $Y2=1.685
cc_342 N_A_c_301_n N_CI_M1005_g 0.00986519f $X=2.35 $Y=1.85 $X2=1.335 $Y2=1.075
cc_343 N_A_c_304_n N_CI_M1014_g 0.00481368f $X=5.01 $Y=1.85 $X2=3.415 $Y2=1.075
cc_344 N_A_c_299_n N_CI_M1009_g 0.00809446f $X=5.13 $Y=2.775 $X2=4.685 $Y2=1.075
cc_345 N_A_c_304_n N_CI_M1009_g 0.00570385f $X=5.01 $Y=1.85 $X2=4.685 $Y2=1.075
cc_346 N_A_c_309_n N_CI_M1009_g 8.57008e-19 $X=5.155 $Y=1.85 $X2=4.685 $Y2=1.075
cc_347 N_A_c_310_n N_CI_M1009_g 0.00116181f $X=5.155 $Y=1.85 $X2=4.685 $Y2=1.075
cc_348 N_A_c_324_n N_CI_M1009_g 0.0805808f $X=5.155 $Y=1.685 $X2=4.685 $Y2=1.075
cc_349 N_A_c_299_n N_CI_M1007_g 0.00831744f $X=5.13 $Y=2.775 $X2=4.685 $Y2=4.585
cc_350 N_A_c_300_n N_CI_M1007_g 0.175024f $X=5.13 $Y=2.925 $X2=4.685 $Y2=4.585
cc_351 N_A_c_294_n N_CI_c_738_n 0.00109073f $X=2.2 $Y=1.76 $X2=3.27 $Y2=2.22
cc_352 N_A_c_297_n N_CI_c_738_n 0.00626944f $X=2.435 $Y=2.81 $X2=3.27 $Y2=2.22
cc_353 N_A_c_301_n N_CI_c_738_n 0.0733404f $X=2.35 $Y=1.85 $X2=3.27 $Y2=2.22
cc_354 N_A_c_304_n N_CI_c_738_n 0.0520212f $X=5.01 $Y=1.85 $X2=3.27 $Y2=2.22
cc_355 N_A_c_305_n N_CI_c_738_n 0.0266076f $X=2.64 $Y=1.85 $X2=3.27 $Y2=2.22
cc_356 N_A_c_307_n N_CI_c_738_n 0.00394572f $X=2.495 $Y=1.85 $X2=3.27 $Y2=2.22
cc_357 N_A_c_317_n N_CI_c_738_n 0.00232838f $X=2.495 $Y=1.76 $X2=3.27 $Y2=2.22
cc_358 N_A_c_301_n N_CI_c_739_n 0.0259569f $X=2.35 $Y=1.85 $X2=1.47 $Y2=2.22
cc_359 N_A_c_304_n N_CI_c_740_n 0.0858968f $X=5.01 $Y=1.85 $X2=4.6 $Y2=2.22
cc_360 N_A_c_304_n N_CI_c_741_n 0.0268181f $X=5.01 $Y=1.85 $X2=3.56 $Y2=2.22
cc_361 N_A_M1010_g CI 0.00555516f $X=0.475 $Y=4.585 $X2=1.325 $Y2=2.22
cc_362 N_A_c_301_n CI 0.0466623f $X=2.35 $Y=1.85 $X2=1.325 $Y2=2.22
cc_363 N_A_c_303_n CI 0.0210627f $X=0.63 $Y=1.85 $X2=1.325 $Y2=2.22
cc_364 N_A_c_306_n CI 0.00205922f $X=0.485 $Y=1.85 $X2=1.325 $Y2=2.22
cc_365 N_A_c_312_n CI 0.00108997f $X=0.485 $Y=1.85 $X2=1.325 $Y2=2.22
cc_366 N_A_c_301_n N_CI_c_743_n 0.00446594f $X=2.35 $Y=1.85 $X2=1.325 $Y2=2.22
cc_367 N_A_c_304_n N_CI_c_744_n 0.00257813f $X=5.01 $Y=1.85 $X2=3.415 $Y2=2.22
cc_368 N_A_c_299_n N_CI_c_745_n 0.00413683f $X=5.13 $Y=2.775 $X2=4.745 $Y2=2.22
cc_369 N_A_c_304_n N_CI_c_745_n 0.0268056f $X=5.01 $Y=1.85 $X2=4.745 $Y2=2.22
cc_370 N_A_c_299_n N_CI_c_746_n 0.00385032f $X=5.13 $Y=2.775 $X2=4.745 $Y2=2.22
cc_371 N_A_c_304_n N_CI_c_746_n 0.00203847f $X=5.01 $Y=1.85 $X2=4.745 $Y2=2.22
cc_372 N_A_c_301_n N_CI_c_747_n 0.00157267f $X=2.35 $Y=1.85 $X2=1.325 $Y2=2.22
cc_373 N_A_c_299_n N_CI_c_748_n 0.0209004f $X=5.13 $Y=2.775 $X2=4.745 $Y2=2.4
cc_374 N_A_c_304_n N_CI_c_748_n 2.31739e-19 $X=5.01 $Y=1.85 $X2=4.745 $Y2=2.4
cc_375 N_A_c_332_n N_CON_c_913_n 9.92167e-19 $X=2.125 $Y=2.96 $X2=1.665
+ $Y2=3.025
cc_376 N_A_c_296_n N_CON_c_913_n 0.00127956f $X=2.2 $Y=2.885 $X2=1.665 $Y2=3.025
cc_377 N_A_c_301_n N_CON_c_913_n 0.00898724f $X=2.35 $Y=1.85 $X2=1.665 $Y2=3.025
cc_378 N_A_c_305_n N_CON_c_913_n 8.75747e-19 $X=2.64 $Y=1.85 $X2=1.665 $Y2=3.025
cc_379 N_A_c_307_n N_CON_c_913_n 0.00126357f $X=2.495 $Y=1.85 $X2=1.665
+ $Y2=3.025
cc_380 N_A_c_317_n N_CON_c_913_n 0.00171426f $X=2.495 $Y=1.76 $X2=1.665
+ $Y2=3.025
cc_381 N_A_c_288_n N_CON_c_916_n 8.12393e-19 $X=2.125 $Y=1.685 $X2=1.665
+ $Y2=1.765
cc_382 N_A_c_301_n N_CON_c_916_n 0.0122304f $X=2.35 $Y=1.85 $X2=1.665 $Y2=1.765
cc_383 N_A_c_305_n N_CON_c_916_n 8.13159e-19 $X=2.64 $Y=1.85 $X2=1.665 $Y2=1.765
cc_384 N_A_c_307_n N_CON_c_916_n 0.00101586f $X=2.495 $Y=1.85 $X2=1.665
+ $Y2=1.765
cc_385 N_A_c_304_n N_CON_c_917_n 0.00283756f $X=5.01 $Y=1.85 $X2=3.845 $Y2=1.85
cc_386 N_A_c_304_n N_CON_c_918_n 0.0171992f $X=5.01 $Y=1.85 $X2=3.97 $Y2=1.85
cc_387 N_A_c_288_n N_CON_c_919_n 0.0105668f $X=2.125 $Y=1.685 $X2=3.825 $Y2=1.48
cc_388 N_A_c_292_n N_CON_c_919_n 0.00146289f $X=2.36 $Y=1.76 $X2=3.825 $Y2=1.48
cc_389 N_A_c_301_n N_CON_c_919_n 0.0546721f $X=2.35 $Y=1.85 $X2=3.825 $Y2=1.48
cc_390 N_A_c_304_n N_CON_c_919_n 0.0991618f $X=5.01 $Y=1.85 $X2=3.825 $Y2=1.48
cc_391 N_A_c_305_n N_CON_c_919_n 0.0265009f $X=2.64 $Y=1.85 $X2=3.825 $Y2=1.48
cc_392 N_A_c_307_n N_CON_c_919_n 0.00363336f $X=2.495 $Y=1.85 $X2=3.825 $Y2=1.48
cc_393 N_A_c_318_n N_CON_c_919_n 0.00989984f $X=2.495 $Y=1.685 $X2=3.825
+ $Y2=1.48
cc_394 N_A_c_288_n N_CON_c_923_n 2.65615e-19 $X=2.125 $Y=1.685 $X2=1.695
+ $Y2=1.48
cc_395 N_A_c_301_n N_CON_c_923_n 0.0250774f $X=2.35 $Y=1.85 $X2=1.695 $Y2=1.48
cc_396 N_A_c_304_n N_CON_c_925_n 0.0740962f $X=5.01 $Y=1.85 $X2=5.995 $Y2=1.48
cc_397 N_A_c_309_n N_CON_c_925_n 0.0265607f $X=5.155 $Y=1.85 $X2=5.995 $Y2=1.48
cc_398 N_A_c_310_n N_CON_c_925_n 0.00405354f $X=5.155 $Y=1.85 $X2=5.995 $Y2=1.48
cc_399 N_A_c_322_n N_CON_c_925_n 0.00213677f $X=5.155 $Y=1.85 $X2=5.995 $Y2=1.48
cc_400 N_A_c_324_n N_CON_c_925_n 0.010321f $X=5.155 $Y=1.685 $X2=5.995 $Y2=1.48
cc_401 N_A_c_304_n N_CON_c_928_n 0.0252799f $X=5.01 $Y=1.85 $X2=4.115 $Y2=1.48
cc_402 N_A_c_304_n N_CON_c_929_n 6.93264e-19 $X=5.01 $Y=1.85 $X2=3.97 $Y2=1.48
cc_403 N_A_c_299_n N_A_784_115#_M1018_g 0.0266804f $X=5.13 $Y=2.775 $X2=5.585
+ $Y2=0.945
cc_404 N_A_c_309_n N_A_784_115#_M1018_g 9.02444e-19 $X=5.155 $Y=1.85 $X2=5.585
+ $Y2=0.945
cc_405 N_A_c_310_n N_A_784_115#_M1018_g 0.00131152f $X=5.155 $Y=1.85 $X2=5.585
+ $Y2=0.945
cc_406 N_A_c_322_n N_A_784_115#_M1018_g 0.0195004f $X=5.155 $Y=1.85 $X2=5.585
+ $Y2=0.945
cc_407 N_A_c_324_n N_A_784_115#_M1018_g 0.0279443f $X=5.155 $Y=1.685 $X2=5.585
+ $Y2=0.945
cc_408 N_A_M1002_g N_A_784_115#_M1001_g 0.0660764f $X=5.095 $Y=4.585 $X2=5.585
+ $Y2=5.085
cc_409 N_A_c_304_n N_A_784_115#_c_1097_n 0.0018868f $X=5.01 $Y=1.85 $X2=4.225
+ $Y2=2.22
cc_410 N_A_c_304_n N_A_784_115#_c_1098_n 7.77654e-19 $X=5.01 $Y=1.85 $X2=3.93
+ $Y2=2.22
cc_411 N_A_M1002_g N_A_784_115#_c_1117_n 0.0193311f $X=5.095 $Y=4.585 $X2=5.33
+ $Y2=3.335
cc_412 N_A_c_300_n N_A_784_115#_c_1117_n 0.0016251f $X=5.13 $Y=2.925 $X2=5.33
+ $Y2=3.335
cc_413 N_A_c_304_n N_A_784_115#_c_1102_n 0.0140552f $X=5.01 $Y=1.85 $X2=4.31
+ $Y2=2.135
cc_414 N_A_c_309_n N_A_784_115#_c_1102_n 0.00192851f $X=5.155 $Y=1.85 $X2=4.31
+ $Y2=2.135
cc_415 N_A_c_310_n N_A_784_115#_c_1102_n 0.00296302f $X=5.155 $Y=1.85 $X2=4.31
+ $Y2=2.135
cc_416 N_A_M1002_g N_A_784_115#_c_1120_n 0.00698879f $X=5.095 $Y=4.585 $X2=5.415
+ $Y2=3.25
cc_417 N_A_c_299_n N_A_784_115#_c_1105_n 0.00675793f $X=5.13 $Y=2.775 $X2=5.415
+ $Y2=2.755
cc_418 N_A_c_299_n N_A_784_115#_c_1106_n 0.0199271f $X=5.13 $Y=2.775 $X2=5.585
+ $Y2=2.755
cc_419 N_A_M1010_g N_A_27_617#_c_1222_n 0.0179393f $X=0.475 $Y=4.585 $X2=1.035
+ $Y2=3.46
cc_420 N_A_c_309_n N_S_c_1246_n 0.00346849f $X=5.155 $Y=1.85 $X2=5.8 $Y2=0.825
cc_421 N_A_c_310_n N_S_c_1246_n 0.00615434f $X=5.155 $Y=1.85 $X2=5.8 $Y2=0.825
cc_422 N_A_M1002_g S 2.86673e-19 $X=5.095 $Y=4.585 $X2=5.8 $Y2=3.365
cc_423 N_A_c_301_n N_A_27_115#_c_1319_n 0.0221351f $X=2.35 $Y=1.85 $X2=1.035
+ $Y2=1.345
cc_424 N_A_c_303_n N_A_27_115#_c_1319_n 0.00620246f $X=0.63 $Y=1.85 $X2=1.035
+ $Y2=1.345
cc_425 N_A_c_306_n N_A_27_115#_c_1319_n 0.00707705f $X=0.485 $Y=1.85 $X2=1.035
+ $Y2=1.345
cc_426 N_A_c_312_n N_A_27_115#_c_1319_n 0.00133715f $X=0.485 $Y=1.85 $X2=1.035
+ $Y2=1.345
cc_427 N_A_c_313_n N_A_27_115#_c_1319_n 0.0150777f $X=0.485 $Y=1.685 $X2=1.035
+ $Y2=1.345
cc_428 N_A_c_306_n N_A_27_115#_c_1330_n 0.0011584f $X=0.485 $Y=1.85 $X2=0.345
+ $Y2=1.345
cc_429 N_A_c_318_n N_A_526_115#_c_1338_n 2.68807e-19 $X=2.495 $Y=1.685 $X2=2.77
+ $Y2=0.825
cc_430 N_A_c_304_n N_A_526_115#_c_1343_n 0.00487455f $X=5.01 $Y=1.85 $X2=3.545
+ $Y2=1.345
cc_431 N_A_c_304_n N_A_526_115#_c_1345_n 8.88228e-19 $X=5.01 $Y=1.85 $X2=2.855
+ $Y2=1.345
cc_432 N_A_c_318_n N_A_526_115#_c_1345_n 4.66174e-19 $X=2.495 $Y=1.685 $X2=2.855
+ $Y2=1.345
cc_433 N_B_M1003_g N_CI_M1005_g 0.0419673f $X=0.905 $Y=1.075 $X2=1.335 $Y2=1.075
cc_434 N_B_M1025_g N_CI_M1005_g 0.0413128f $X=1.765 $Y=1.075 $X2=1.335 $Y2=1.075
cc_435 N_B_M1003_g N_CI_M1004_g 0.0101134f $X=0.905 $Y=1.075 $X2=1.335 $Y2=4.585
cc_436 N_B_M1000_g N_CI_M1004_g 0.0376075f $X=0.905 $Y=4.585 $X2=1.335 $Y2=4.585
cc_437 N_B_c_508_n N_CI_M1004_g 0.00162835f $X=0.895 $Y=2.76 $X2=1.335 $Y2=4.585
cc_438 N_B_c_509_n N_CI_M1004_g 0.0188528f $X=0.895 $Y=2.76 $X2=1.335 $Y2=4.585
cc_439 N_B_c_511_n N_CI_M1004_g 0.0572759f $X=2.015 $Y=2.43 $X2=1.335 $Y2=4.585
cc_440 N_B_c_512_n N_CI_M1004_g 0.0102981f $X=2.16 $Y=2.59 $X2=1.335 $Y2=4.585
cc_441 N_B_M1022_g N_CI_M1014_g 0.0184719f $X=2.985 $Y=4.585 $X2=3.415 $Y2=1.075
cc_442 N_B_c_521_n N_CI_M1014_g 0.00290674f $X=2.975 $Y=1.85 $X2=3.415 $Y2=1.075
cc_443 N_B_c_522_n N_CI_M1014_g 0.0199829f $X=2.975 $Y=1.85 $X2=3.415 $Y2=1.075
cc_444 N_B_c_523_n N_CI_M1014_g 0.0378945f $X=2.975 $Y=1.685 $X2=3.415 $Y2=1.075
cc_445 N_B_M1022_g N_CI_M1011_g 0.0615923f $X=2.985 $Y=4.585 $X2=3.415 $Y2=4.585
cc_446 N_B_M1017_g N_CI_M1009_g 0.0981211f $X=4.275 $Y=1.075 $X2=4.685 $Y2=1.075
cc_447 N_B_M1016_g N_CI_M1007_g 0.174408f $X=4.275 $Y=4.585 $X2=4.685 $Y2=4.585
cc_448 N_B_M1022_g N_CI_c_736_n 6.79377e-19 $X=2.985 $Y=4.585 $X2=3.415 $Y2=2.59
cc_449 N_B_c_517_n N_CI_c_736_n 0.0188576f $X=3.67 $Y=2.592 $X2=3.415 $Y2=2.59
cc_450 N_B_c_521_n N_CI_c_736_n 0.0103583f $X=2.975 $Y=1.85 $X2=3.415 $Y2=2.59
cc_451 N_B_M1022_g N_CI_c_737_n 0.0204315f $X=2.985 $Y=4.585 $X2=3.415 $Y2=2.59
cc_452 N_B_c_517_n N_CI_c_737_n 0.0120043f $X=3.67 $Y=2.592 $X2=3.415 $Y2=2.59
cc_453 N_B_c_521_n N_CI_c_737_n 9.41528e-19 $X=2.975 $Y=1.85 $X2=3.415 $Y2=2.59
cc_454 N_B_M1025_g N_CI_c_738_n 0.00219877f $X=1.765 $Y=1.075 $X2=3.27 $Y2=2.22
cc_455 N_B_M1022_g N_CI_c_738_n 0.00107346f $X=2.985 $Y=4.585 $X2=3.27 $Y2=2.22
cc_456 N_B_c_510_n N_CI_c_738_n 0.00748189f $X=2.015 $Y=2.43 $X2=3.27 $Y2=2.22
cc_457 N_B_c_511_n N_CI_c_738_n 0.00482273f $X=2.015 $Y=2.43 $X2=3.27 $Y2=2.22
cc_458 N_B_c_512_n N_CI_c_738_n 0.055048f $X=2.16 $Y=2.59 $X2=3.27 $Y2=2.22
cc_459 N_B_c_514_n N_CI_c_738_n 0.0323265f $X=2.83 $Y=2.59 $X2=3.27 $Y2=2.22
cc_460 N_B_c_515_n N_CI_c_738_n 0.0269315f $X=2.45 $Y=2.59 $X2=3.27 $Y2=2.22
cc_461 N_B_c_517_n N_CI_c_738_n 0.0380655f $X=3.67 $Y=2.592 $X2=3.27 $Y2=2.22
cc_462 N_B_c_519_n N_CI_c_738_n 0.0023297f $X=2.305 $Y=2.59 $X2=3.27 $Y2=2.22
cc_463 N_B_c_521_n N_CI_c_738_n 0.0164089f $X=2.975 $Y=1.85 $X2=3.27 $Y2=2.22
cc_464 N_B_c_522_n N_CI_c_738_n 0.00159733f $X=2.975 $Y=1.85 $X2=3.27 $Y2=2.22
cc_465 N_B_M1003_g N_CI_c_739_n 8.6716e-19 $X=0.905 $Y=1.075 $X2=1.47 $Y2=2.22
cc_466 N_B_c_512_n N_CI_c_739_n 0.0259579f $X=2.16 $Y=2.59 $X2=1.47 $Y2=2.22
cc_467 N_B_M1017_g N_CI_c_740_n 0.00112864f $X=4.275 $Y=1.075 $X2=4.6 $Y2=2.22
cc_468 N_B_c_516_n N_CI_c_740_n 0.062156f $X=4.06 $Y=2.592 $X2=4.6 $Y2=2.22
cc_469 N_B_c_517_n N_CI_c_740_n 0.0092809f $X=3.67 $Y=2.592 $X2=4.6 $Y2=2.22
cc_470 N_B_c_520_n N_CI_c_740_n 0.00192504f $X=4.265 $Y=2.59 $X2=4.6 $Y2=2.22
cc_471 N_B_c_527_n N_CI_c_740_n 0.00116782f $X=4.265 $Y=2.59 $X2=4.6 $Y2=2.22
cc_472 N_B_M1022_g N_CI_c_741_n 8.88888e-19 $X=2.985 $Y=4.585 $X2=3.56 $Y2=2.22
cc_473 N_B_c_517_n N_CI_c_741_n 0.0247742f $X=3.67 $Y=2.592 $X2=3.56 $Y2=2.22
cc_474 N_B_c_521_n N_CI_c_741_n 0.00213923f $X=2.975 $Y=1.85 $X2=3.56 $Y2=2.22
cc_475 N_B_M1003_g CI 0.00562571f $X=0.905 $Y=1.075 $X2=1.325 $Y2=2.22
cc_476 N_B_c_508_n CI 2.90821e-19 $X=0.895 $Y=2.76 $X2=1.325 $Y2=2.22
cc_477 N_B_c_509_n CI 5.74814e-19 $X=0.895 $Y=2.76 $X2=1.325 $Y2=2.22
cc_478 N_B_c_512_n CI 0.0466415f $X=2.16 $Y=2.59 $X2=1.325 $Y2=2.22
cc_479 N_B_c_513_n CI 0.0211771f $X=0.63 $Y=2.59 $X2=1.325 $Y2=2.22
cc_480 N_B_c_518_n CI 0.00110643f $X=0.485 $Y=2.59 $X2=1.325 $Y2=2.22
cc_481 N_B_M1003_g N_CI_c_743_n 0.00277751f $X=0.905 $Y=1.075 $X2=1.325 $Y2=2.22
cc_482 N_B_M1025_g N_CI_c_743_n 4.162e-19 $X=1.765 $Y=1.075 $X2=1.325 $Y2=2.22
cc_483 N_B_c_512_n N_CI_c_743_n 0.00446594f $X=2.16 $Y=2.59 $X2=1.325 $Y2=2.22
cc_484 N_B_M1022_g N_CI_c_744_n 0.00154506f $X=2.985 $Y=4.585 $X2=3.415 $Y2=2.22
cc_485 N_B_c_517_n N_CI_c_744_n 8.40427e-19 $X=3.67 $Y=2.592 $X2=3.415 $Y2=2.22
cc_486 N_B_c_521_n N_CI_c_744_n 0.016155f $X=2.975 $Y=1.85 $X2=3.415 $Y2=2.22
cc_487 N_B_M1017_g N_CI_c_745_n 4.28504e-19 $X=4.275 $Y=1.075 $X2=4.745 $Y2=2.22
cc_488 N_B_M1017_g N_CI_c_746_n 0.00109484f $X=4.275 $Y=1.075 $X2=4.745 $Y2=2.22
cc_489 N_B_c_516_n N_CI_c_746_n 0.00164652f $X=4.06 $Y=2.592 $X2=4.745 $Y2=2.22
cc_490 N_B_c_520_n N_CI_c_746_n 0.00317294f $X=4.265 $Y=2.59 $X2=4.745 $Y2=2.22
cc_491 N_B_c_527_n N_CI_c_746_n 5.51285e-19 $X=4.265 $Y=2.59 $X2=4.745 $Y2=2.22
cc_492 N_B_M1003_g N_CI_c_747_n 0.0219985f $X=0.905 $Y=1.075 $X2=1.325 $Y2=2.22
cc_493 N_B_M1025_g N_CI_c_747_n 0.0193664f $X=1.765 $Y=1.075 $X2=1.325 $Y2=2.22
cc_494 N_B_c_512_n N_CI_c_747_n 0.00157267f $X=2.16 $Y=2.59 $X2=1.325 $Y2=2.22
cc_495 N_B_c_516_n N_CI_c_748_n 9.10645e-19 $X=4.06 $Y=2.592 $X2=4.745 $Y2=2.4
cc_496 N_B_c_520_n N_CI_c_748_n 0.00282159f $X=4.265 $Y=2.59 $X2=4.745 $Y2=2.4
cc_497 N_B_c_527_n N_CI_c_748_n 0.0208261f $X=4.265 $Y=2.59 $X2=4.745 $Y2=2.4
cc_498 N_B_M1017_g N_CON_c_906_n 0.0384031f $X=4.275 $Y=1.075 $X2=3.845
+ $Y2=1.685
cc_499 N_B_M1017_g N_CON_M1013_g 0.0179106f $X=4.275 $Y=1.075 $X2=3.845
+ $Y2=4.585
cc_500 N_B_M1016_g N_CON_M1013_g 0.04207f $X=4.275 $Y=4.585 $X2=3.845 $Y2=4.585
cc_501 N_B_c_520_n N_CON_M1013_g 4.28168e-19 $X=4.265 $Y=2.59 $X2=3.845
+ $Y2=4.585
cc_502 N_B_c_527_n N_CON_M1013_g 0.0211897f $X=4.265 $Y=2.59 $X2=3.845 $Y2=4.585
cc_503 N_B_M1025_g N_CON_c_913_n 0.0112485f $X=1.765 $Y=1.075 $X2=1.665
+ $Y2=3.025
cc_504 N_B_M1023_g N_CON_c_913_n 0.0204831f $X=1.765 $Y=4.585 $X2=1.665
+ $Y2=3.025
cc_505 N_B_c_508_n N_CON_c_913_n 0.00630121f $X=0.895 $Y=2.76 $X2=1.665
+ $Y2=3.025
cc_506 N_B_c_510_n N_CON_c_913_n 0.0257712f $X=2.015 $Y=2.43 $X2=1.665 $Y2=3.025
cc_507 N_B_c_511_n N_CON_c_913_n 0.00754141f $X=2.015 $Y=2.43 $X2=1.665
+ $Y2=3.025
cc_508 N_B_c_512_n N_CON_c_913_n 0.0208106f $X=2.16 $Y=2.59 $X2=1.665 $Y2=3.025
cc_509 N_B_c_515_n N_CON_c_913_n 0.00105333f $X=2.45 $Y=2.59 $X2=1.665 $Y2=3.025
cc_510 N_B_M1025_g N_CON_c_916_n 0.00525936f $X=1.765 $Y=1.075 $X2=1.665
+ $Y2=1.765
cc_511 N_B_M1017_g N_CON_c_917_n 0.0200025f $X=4.275 $Y=1.075 $X2=3.845 $Y2=1.85
cc_512 N_B_M1017_g N_CON_c_918_n 7.2637e-19 $X=4.275 $Y=1.075 $X2=3.97 $Y2=1.85
cc_513 N_B_c_521_n N_CON_c_918_n 0.0022487f $X=2.975 $Y=1.85 $X2=3.97 $Y2=1.85
cc_514 N_B_M1025_g N_CON_c_919_n 0.00888363f $X=1.765 $Y=1.075 $X2=3.825
+ $Y2=1.48
cc_515 N_B_c_521_n N_CON_c_919_n 0.00143374f $X=2.975 $Y=1.85 $X2=3.825 $Y2=1.48
cc_516 N_B_c_522_n N_CON_c_919_n 0.00159733f $X=2.975 $Y=1.85 $X2=3.825 $Y2=1.48
cc_517 N_B_c_523_n N_CON_c_919_n 0.00280657f $X=2.975 $Y=1.685 $X2=3.825
+ $Y2=1.48
cc_518 N_B_M1003_g N_CON_c_923_n 7.56281e-19 $X=0.905 $Y=1.075 $X2=1.695
+ $Y2=1.48
cc_519 N_B_M1025_g N_CON_c_923_n 0.0026062f $X=1.765 $Y=1.075 $X2=1.695 $Y2=1.48
cc_520 N_B_M1017_g N_CON_c_925_n 0.001558f $X=4.275 $Y=1.075 $X2=5.995 $Y2=1.48
cc_521 N_B_M1017_g N_CON_c_928_n 9.72315e-19 $X=4.275 $Y=1.075 $X2=4.115
+ $Y2=1.48
cc_522 N_B_M1017_g N_CON_c_929_n 0.0018911f $X=4.275 $Y=1.075 $X2=3.97 $Y2=1.48
cc_523 N_B_M1025_g N_CON_c_932_n 0.00500773f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_524 N_B_M1017_g N_A_784_115#_c_1096_n 0.00218215f $X=4.275 $Y=1.075 $X2=3.845
+ $Y2=3.03
cc_525 N_B_M1016_g N_A_784_115#_c_1096_n 0.00502446f $X=4.275 $Y=4.585 $X2=3.845
+ $Y2=3.03
cc_526 N_B_c_516_n N_A_784_115#_c_1096_n 0.0204781f $X=4.06 $Y=2.592 $X2=3.845
+ $Y2=3.03
cc_527 N_B_c_520_n N_A_784_115#_c_1096_n 0.0120274f $X=4.265 $Y=2.59 $X2=3.845
+ $Y2=3.03
cc_528 N_B_c_527_n N_A_784_115#_c_1096_n 0.003498f $X=4.265 $Y=2.59 $X2=3.845
+ $Y2=3.03
cc_529 N_B_M1017_g N_A_784_115#_c_1097_n 0.00690261f $X=4.275 $Y=1.075 $X2=4.225
+ $Y2=2.22
cc_530 N_B_c_516_n N_A_784_115#_c_1097_n 0.00247487f $X=4.06 $Y=2.592 $X2=4.225
+ $Y2=2.22
cc_531 N_B_c_520_n N_A_784_115#_c_1097_n 0.016625f $X=4.265 $Y=2.59 $X2=4.225
+ $Y2=2.22
cc_532 N_B_c_527_n N_A_784_115#_c_1097_n 0.00274037f $X=4.265 $Y=2.59 $X2=4.225
+ $Y2=2.22
cc_533 N_B_M1017_g N_A_784_115#_c_1099_n 3.31145e-19 $X=4.275 $Y=1.075 $X2=4.06
+ $Y2=0.905
cc_534 N_B_M1016_g N_A_784_115#_c_1113_n 0.00221174f $X=4.275 $Y=4.585 $X2=4.06
+ $Y2=3.42
cc_535 N_B_c_516_n N_A_784_115#_c_1113_n 0.00840219f $X=4.06 $Y=2.592 $X2=4.06
+ $Y2=3.42
cc_536 N_B_c_520_n N_A_784_115#_c_1113_n 0.0015127f $X=4.265 $Y=2.59 $X2=4.06
+ $Y2=3.42
cc_537 N_B_c_527_n N_A_784_115#_c_1113_n 3.44204e-19 $X=4.265 $Y=2.59 $X2=4.06
+ $Y2=3.42
cc_538 N_B_M1016_g N_A_784_115#_c_1117_n 0.0162839f $X=4.275 $Y=4.585 $X2=5.33
+ $Y2=3.335
cc_539 N_B_c_516_n N_A_784_115#_c_1117_n 0.00471773f $X=4.06 $Y=2.592 $X2=5.33
+ $Y2=3.335
cc_540 N_B_c_520_n N_A_784_115#_c_1117_n 0.00328494f $X=4.265 $Y=2.59 $X2=5.33
+ $Y2=3.335
cc_541 N_B_M1017_g N_A_784_115#_c_1102_n 0.0251036f $X=4.275 $Y=1.075 $X2=4.31
+ $Y2=2.135
cc_542 N_B_M1017_g N_A_784_115#_c_1103_n 0.00797271f $X=4.275 $Y=1.075 $X2=4.31
+ $Y2=0.99
cc_543 N_B_M1000_g N_A_27_617#_c_1222_n 0.0163254f $X=0.905 $Y=4.585 $X2=1.035
+ $Y2=3.46
cc_544 N_B_c_508_n N_A_27_617#_c_1222_n 0.0124135f $X=0.895 $Y=2.76 $X2=1.035
+ $Y2=3.46
cc_545 N_B_c_509_n N_A_27_617#_c_1222_n 0.00110112f $X=0.895 $Y=2.76 $X2=1.035
+ $Y2=3.46
cc_546 N_B_c_518_n N_A_27_617#_c_1222_n 0.00457576f $X=0.485 $Y=2.59 $X2=1.035
+ $Y2=3.46
cc_547 N_B_M1022_g N_A_526_617#_c_1235_n 0.0167311f $X=2.985 $Y=4.585 $X2=3.545
+ $Y2=3.455
cc_548 N_B_c_521_n N_A_526_617#_c_1235_n 0.00240309f $X=2.975 $Y=1.85 $X2=3.545
+ $Y2=3.455
cc_549 N_B_M1003_g N_A_27_115#_c_1319_n 0.0143352f $X=0.905 $Y=1.075 $X2=1.035
+ $Y2=1.345
cc_550 N_B_M1003_g N_A_27_115#_c_1321_n 2.68807e-19 $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_551 N_B_c_523_n N_A_526_115#_c_1338_n 2.68807e-19 $X=2.975 $Y=1.685 $X2=2.77
+ $Y2=0.825
cc_552 N_B_c_521_n N_A_526_115#_c_1343_n 0.00664394f $X=2.975 $Y=1.85 $X2=3.545
+ $Y2=1.345
cc_553 N_B_c_522_n N_A_526_115#_c_1343_n 0.00217805f $X=2.975 $Y=1.85 $X2=3.545
+ $Y2=1.345
cc_554 N_B_c_523_n N_A_526_115#_c_1343_n 0.0131914f $X=2.975 $Y=1.685 $X2=3.545
+ $Y2=1.345
cc_555 N_B_c_522_n N_A_526_115#_c_1345_n 4.88342e-19 $X=2.975 $Y=1.85 $X2=2.855
+ $Y2=1.345
cc_556 N_CI_M1014_g N_CON_c_906_n 0.0248153f $X=3.415 $Y=1.075 $X2=3.845
+ $Y2=1.685
cc_557 N_CI_M1014_g N_CON_M1013_g 0.0190239f $X=3.415 $Y=1.075 $X2=3.845
+ $Y2=4.585
cc_558 N_CI_M1011_g N_CON_M1013_g 0.0435751f $X=3.415 $Y=4.585 $X2=3.845
+ $Y2=4.585
cc_559 N_CI_c_736_n N_CON_M1013_g 4.41794e-19 $X=3.415 $Y=2.59 $X2=3.845
+ $Y2=4.585
cc_560 N_CI_c_737_n N_CON_M1013_g 0.0196718f $X=3.415 $Y=2.59 $X2=3.845
+ $Y2=4.585
cc_561 N_CI_c_740_n N_CON_M1013_g 9.30638e-19 $X=4.6 $Y=2.22 $X2=3.845 $Y2=4.585
cc_562 N_CI_c_741_n N_CON_M1013_g 4.44444e-19 $X=3.56 $Y=2.22 $X2=3.845
+ $Y2=4.585
cc_563 N_CI_c_744_n N_CON_M1013_g 9.22089e-19 $X=3.415 $Y=2.22 $X2=3.845
+ $Y2=4.585
cc_564 N_CI_M1005_g N_CON_c_913_n 0.00386404f $X=1.335 $Y=1.075 $X2=1.665
+ $Y2=3.025
cc_565 N_CI_M1004_g N_CON_c_913_n 0.0126133f $X=1.335 $Y=4.585 $X2=1.665
+ $Y2=3.025
cc_566 N_CI_c_738_n N_CON_c_913_n 0.0138278f $X=3.27 $Y=2.22 $X2=1.665 $Y2=3.025
cc_567 N_CI_c_739_n N_CON_c_913_n 0.00183606f $X=1.47 $Y=2.22 $X2=1.665
+ $Y2=3.025
cc_568 N_CI_c_743_n N_CON_c_913_n 0.0223962f $X=1.325 $Y=2.22 $X2=1.665
+ $Y2=3.025
cc_569 N_CI_c_747_n N_CON_c_913_n 0.00170665f $X=1.325 $Y=2.22 $X2=1.665
+ $Y2=3.025
cc_570 N_CI_M1005_g N_CON_c_916_n 0.00402444f $X=1.335 $Y=1.075 $X2=1.665
+ $Y2=1.765
cc_571 N_CI_c_738_n N_CON_c_916_n 7.55969e-19 $X=3.27 $Y=2.22 $X2=1.665
+ $Y2=1.765
cc_572 N_CI_M1014_g N_CON_c_917_n 0.02064f $X=3.415 $Y=1.075 $X2=3.845 $Y2=1.85
cc_573 N_CI_c_740_n N_CON_c_917_n 0.00158152f $X=4.6 $Y=2.22 $X2=3.845 $Y2=1.85
cc_574 N_CI_M1014_g N_CON_c_918_n 0.00127353f $X=3.415 $Y=1.075 $X2=3.97
+ $Y2=1.85
cc_575 N_CI_c_740_n N_CON_c_918_n 0.00187655f $X=4.6 $Y=2.22 $X2=3.97 $Y2=1.85
cc_576 N_CI_M1014_g N_CON_c_919_n 0.00314002f $X=3.415 $Y=1.075 $X2=3.825
+ $Y2=1.48
cc_577 N_CI_M1005_g N_CON_c_923_n 0.00532501f $X=1.335 $Y=1.075 $X2=1.695
+ $Y2=1.48
cc_578 N_CI_M1009_g N_CON_c_925_n 0.0107454f $X=4.685 $Y=1.075 $X2=5.995
+ $Y2=1.48
cc_579 N_CI_M1014_g N_CON_c_929_n 0.00211142f $X=3.415 $Y=1.075 $X2=3.97
+ $Y2=1.48
cc_580 N_CI_M1005_g N_CON_c_932_n 0.00480051f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_581 N_CI_M1014_g N_A_784_115#_c_1096_n 3.97727e-19 $X=3.415 $Y=1.075
+ $X2=3.845 $Y2=3.03
cc_582 N_CI_M1011_g N_A_784_115#_c_1096_n 0.00502446f $X=3.415 $Y=4.585
+ $X2=3.845 $Y2=3.03
cc_583 N_CI_c_736_n N_A_784_115#_c_1096_n 0.0114194f $X=3.415 $Y=2.59 $X2=3.845
+ $Y2=3.03
cc_584 N_CI_c_737_n N_A_784_115#_c_1096_n 0.00241496f $X=3.415 $Y=2.59 $X2=3.845
+ $Y2=3.03
cc_585 N_CI_c_741_n N_A_784_115#_c_1096_n 8.66056e-19 $X=3.56 $Y=2.22 $X2=3.845
+ $Y2=3.03
cc_586 N_CI_c_744_n N_A_784_115#_c_1096_n 0.0104334f $X=3.415 $Y=2.22 $X2=3.845
+ $Y2=3.03
cc_587 N_CI_M1009_g N_A_784_115#_c_1097_n 8.45664e-19 $X=4.685 $Y=1.075
+ $X2=4.225 $Y2=2.22
cc_588 N_CI_c_740_n N_A_784_115#_c_1097_n 0.0202332f $X=4.6 $Y=2.22 $X2=4.225
+ $Y2=2.22
cc_589 N_CI_c_746_n N_A_784_115#_c_1097_n 0.00742016f $X=4.745 $Y=2.22 $X2=4.225
+ $Y2=2.22
cc_590 N_CI_M1014_g N_A_784_115#_c_1098_n 5.06918e-19 $X=3.415 $Y=1.075 $X2=3.93
+ $Y2=2.22
cc_591 N_CI_c_740_n N_A_784_115#_c_1098_n 0.00872498f $X=4.6 $Y=2.22 $X2=3.93
+ $Y2=2.22
cc_592 N_CI_c_744_n N_A_784_115#_c_1098_n 0.00810858f $X=3.415 $Y=2.22 $X2=3.93
+ $Y2=2.22
cc_593 N_CI_M1011_g N_A_784_115#_c_1113_n 0.00150127f $X=3.415 $Y=4.585 $X2=4.06
+ $Y2=3.42
cc_594 N_CI_M1007_g N_A_784_115#_c_1117_n 0.0193185f $X=4.685 $Y=4.585 $X2=5.33
+ $Y2=3.335
cc_595 N_CI_c_748_n N_A_784_115#_c_1117_n 0.00136691f $X=4.745 $Y=2.4 $X2=5.33
+ $Y2=3.335
cc_596 N_CI_M1009_g N_A_784_115#_c_1102_n 0.0110662f $X=4.685 $Y=1.075 $X2=4.31
+ $Y2=2.135
cc_597 N_CI_c_745_n N_A_784_115#_c_1102_n 0.00139142f $X=4.745 $Y=2.22 $X2=4.31
+ $Y2=2.135
cc_598 N_CI_M1011_g N_A_526_617#_c_1235_n 0.0191262f $X=3.415 $Y=4.585 $X2=3.545
+ $Y2=3.455
cc_599 N_CI_c_737_n N_A_526_617#_c_1235_n 9.07588e-19 $X=3.415 $Y=2.59 $X2=3.545
+ $Y2=3.455
cc_600 N_CI_c_747_n N_A_27_115#_c_1319_n 3.85943e-19 $X=1.325 $Y=2.22 $X2=1.035
+ $Y2=1.345
cc_601 N_CI_M1005_g N_A_27_115#_c_1321_n 2.68807e-19 $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_602 N_CI_M1014_g N_A_526_115#_c_1343_n 0.0151472f $X=3.415 $Y=1.075 $X2=3.545
+ $Y2=1.345
cc_603 N_CI_M1014_g N_A_526_115#_c_1346_n 2.68807e-19 $X=3.415 $Y=1.075 $X2=3.63
+ $Y2=0.825
cc_604 N_CON_c_925_n N_A_784_115#_M1015_d 0.0013709f $X=5.995 $Y=1.48 $X2=3.92
+ $Y2=0.575
cc_605 N_CON_c_928_n N_A_784_115#_M1015_d 0.00383935f $X=4.115 $Y=1.48 $X2=3.92
+ $Y2=0.575
cc_606 N_CON_c_929_n N_A_784_115#_M1015_d 0.00149447f $X=3.97 $Y=1.48 $X2=3.92
+ $Y2=0.575
cc_607 N_CON_c_914_n N_A_784_115#_M1018_g 0.00198469f $X=6.41 $Y=2.74 $X2=5.585
+ $Y2=0.945
cc_608 N_CON_c_925_n N_A_784_115#_M1018_g 0.0170447f $X=5.995 $Y=1.48 $X2=5.585
+ $Y2=0.945
cc_609 N_CON_M1013_g N_A_784_115#_c_1096_n 0.0136798f $X=3.845 $Y=4.585
+ $X2=3.845 $Y2=3.03
cc_610 N_CON_c_917_n N_A_784_115#_c_1097_n 0.00118003f $X=3.845 $Y=1.85
+ $X2=4.225 $Y2=2.22
cc_611 N_CON_c_918_n N_A_784_115#_c_1097_n 0.00732851f $X=3.97 $Y=1.85 $X2=4.225
+ $Y2=2.22
cc_612 N_CON_M1013_g N_A_784_115#_c_1098_n 0.00624765f $X=3.845 $Y=4.585
+ $X2=3.93 $Y2=2.22
cc_613 N_CON_c_917_n N_A_784_115#_c_1098_n 4.82273e-19 $X=3.845 $Y=1.85 $X2=3.93
+ $Y2=2.22
cc_614 N_CON_c_918_n N_A_784_115#_c_1098_n 0.00939629f $X=3.97 $Y=1.85 $X2=3.93
+ $Y2=2.22
cc_615 N_CON_c_906_n N_A_784_115#_c_1099_n 2.68807e-19 $X=3.845 $Y=1.685
+ $X2=4.06 $Y2=0.905
cc_616 N_CON_M1013_g N_A_784_115#_c_1113_n 0.0124031f $X=3.845 $Y=4.585 $X2=4.06
+ $Y2=3.42
cc_617 N_CON_c_906_n N_A_784_115#_c_1102_n 0.00148932f $X=3.845 $Y=1.685
+ $X2=4.31 $Y2=2.135
cc_618 N_CON_M1013_g N_A_784_115#_c_1102_n 7.13673e-19 $X=3.845 $Y=4.585
+ $X2=4.31 $Y2=2.135
cc_619 N_CON_c_917_n N_A_784_115#_c_1102_n 8.78503e-19 $X=3.845 $Y=1.85 $X2=4.31
+ $Y2=2.135
cc_620 N_CON_c_918_n N_A_784_115#_c_1102_n 0.0115992f $X=3.97 $Y=1.85 $X2=4.31
+ $Y2=2.135
cc_621 N_CON_c_925_n N_A_784_115#_c_1102_n 0.0156075f $X=5.995 $Y=1.48 $X2=4.31
+ $Y2=2.135
cc_622 N_CON_c_928_n N_A_784_115#_c_1102_n 0.00193898f $X=4.115 $Y=1.48 $X2=4.31
+ $Y2=2.135
cc_623 N_CON_c_929_n N_A_784_115#_c_1102_n 0.0253848f $X=3.97 $Y=1.48 $X2=4.31
+ $Y2=2.135
cc_624 N_CON_c_925_n N_A_784_115#_c_1103_n 0.00469291f $X=5.995 $Y=1.48 $X2=4.31
+ $Y2=0.99
cc_625 N_CON_c_928_n N_A_784_115#_c_1103_n 0.00462554f $X=4.115 $Y=1.48 $X2=4.31
+ $Y2=0.99
cc_626 N_CON_c_929_n N_A_784_115#_c_1103_n 0.00254859f $X=3.97 $Y=1.48 $X2=4.31
+ $Y2=0.99
cc_627 N_CON_c_915_n N_A_784_115#_c_1106_n 0.00451843f $X=6.41 $Y=2.74 $X2=5.585
+ $Y2=2.755
cc_628 N_CON_M1021_g N_S_c_1246_n 0.0112727f $X=6.535 $Y=0.945 $X2=5.8 $Y2=0.825
cc_629 N_CON_c_914_n N_S_c_1246_n 0.0216008f $X=6.41 $Y=2.74 $X2=5.8 $Y2=0.825
cc_630 N_CON_c_925_n N_S_c_1246_n 0.0230501f $X=5.995 $Y=1.48 $X2=5.8 $Y2=0.825
cc_631 CON N_S_c_1246_n 0.00260317f $X=6.14 $Y=1.48 $X2=5.8 $Y2=0.825
cc_632 N_CON_c_936_n N_S_c_1246_n 0.0121035f $X=6.41 $Y=1.48 $X2=5.8 $Y2=0.825
cc_633 N_CON_M1021_g N_S_c_1251_n 0.00130367f $X=6.535 $Y=0.945 $X2=5.925
+ $Y2=3.165
cc_634 N_CON_M1008_g N_S_c_1251_n 0.00437761f $X=6.535 $Y=5.085 $X2=5.925
+ $Y2=3.165
cc_635 N_CON_c_914_n N_S_c_1251_n 0.0278588f $X=6.41 $Y=2.74 $X2=5.925 $Y2=3.165
cc_636 N_CON_c_915_n N_S_c_1251_n 0.00305399f $X=6.41 $Y=2.74 $X2=5.925
+ $Y2=3.165
cc_637 N_CON_M1021_g N_S_c_1252_n 8.65886e-19 $X=6.535 $Y=0.945 $X2=5.925
+ $Y2=2.22
cc_638 N_CON_c_914_n N_S_c_1252_n 0.00863446f $X=6.41 $Y=2.74 $X2=5.925 $Y2=2.22
cc_639 N_CON_c_925_n N_S_c_1252_n 0.00384217f $X=5.995 $Y=1.48 $X2=5.925
+ $Y2=2.22
cc_640 CON N_S_c_1252_n 5.03075e-19 $X=6.14 $Y=1.48 $X2=5.925 $Y2=2.22
cc_641 N_CON_M1008_g N_S_c_1254_n 0.00293837f $X=6.535 $Y=5.085 $X2=5.925
+ $Y2=3.25
cc_642 N_CON_M1008_g S 0.0029718f $X=6.535 $Y=5.085 $X2=5.8 $Y2=3.365
cc_643 N_CON_M1008_g N_S_c_1256_n 0.022505f $X=6.535 $Y=5.085 $X2=5.8 $Y2=3.365
cc_644 N_CON_M1008_g CO 0.00944261f $X=6.535 $Y=5.085 $X2=6.75 $Y2=2.96
cc_645 N_CON_c_914_n CO 0.0017516f $X=6.41 $Y=2.74 $X2=6.75 $Y2=2.96
cc_646 N_CON_c_915_n CO 0.00612215f $X=6.41 $Y=2.74 $X2=6.75 $Y2=2.96
cc_647 N_CON_M1021_g N_CO_c_1300_n 0.0890511f $X=6.535 $Y=0.945 $X2=6.75
+ $Y2=0.825
cc_648 N_CON_c_914_n N_CO_c_1300_n 0.0950906f $X=6.41 $Y=2.74 $X2=6.75 $Y2=0.825
cc_649 CON N_CO_c_1300_n 0.00209642f $X=6.14 $Y=1.48 $X2=6.75 $Y2=0.825
cc_650 N_CON_c_936_n N_CO_c_1300_n 0.0122992f $X=6.41 $Y=1.48 $X2=6.75 $Y2=0.825
cc_651 N_CON_c_923_n N_A_27_115#_c_1319_n 0.00186751f $X=1.695 $Y=1.48 $X2=1.035
+ $Y2=1.345
cc_652 N_CON_c_932_n N_A_27_115#_c_1321_n 2.23682e-19 $X=1.55 $Y=0.825 $X2=1.12
+ $Y2=0.825
cc_653 N_CON_c_919_n A_368_115# 0.0100396f $X=3.825 $Y=1.48 $X2=1.84 $Y2=0.575
cc_654 N_CON_c_919_n N_A_526_115#_M1020_d 0.00434306f $X=3.825 $Y=1.48 $X2=2.63
+ $Y2=0.575
cc_655 N_CON_c_919_n N_A_526_115#_M1014_d 0.00424073f $X=3.825 $Y=1.48 $X2=3.49
+ $Y2=0.575
cc_656 N_CON_c_906_n N_A_526_115#_c_1343_n 3.23974e-19 $X=3.845 $Y=1.685
+ $X2=3.545 $Y2=1.345
cc_657 N_CON_c_918_n N_A_526_115#_c_1343_n 0.00122114f $X=3.97 $Y=1.85 $X2=3.545
+ $Y2=1.345
cc_658 N_CON_c_919_n N_A_526_115#_c_1343_n 0.0551297f $X=3.825 $Y=1.48 $X2=3.545
+ $Y2=1.345
cc_659 N_CON_c_928_n N_A_526_115#_c_1343_n 0.00103977f $X=4.115 $Y=1.48
+ $X2=3.545 $Y2=1.345
cc_660 N_CON_c_929_n N_A_526_115#_c_1343_n 0.00179176f $X=3.97 $Y=1.48 $X2=3.545
+ $Y2=1.345
cc_661 N_CON_c_919_n N_A_526_115#_c_1345_n 0.0147728f $X=3.825 $Y=1.48 $X2=2.855
+ $Y2=1.345
cc_662 N_CON_c_906_n N_A_526_115#_c_1346_n 2.68807e-19 $X=3.845 $Y=1.685
+ $X2=3.63 $Y2=0.825
cc_663 N_CON_c_925_n A_870_115# 0.0102308f $X=5.995 $Y=1.48 $X2=4.35 $Y2=0.575
cc_664 N_CON_c_925_n A_952_115# 0.0121403f $X=5.995 $Y=1.48 $X2=4.76 $Y2=0.575
cc_665 N_A_784_115#_c_1117_n A_870_617# 0.0106531f $X=5.33 $Y=3.335 $X2=4.35
+ $Y2=3.085
cc_666 N_A_784_115#_c_1117_n A_952_617# 0.00986639f $X=5.33 $Y=3.335 $X2=4.76
+ $Y2=3.085
cc_667 N_A_784_115#_M1018_g N_S_c_1246_n 0.0338104f $X=5.585 $Y=0.945 $X2=5.8
+ $Y2=0.825
cc_668 N_A_784_115#_M1018_g N_S_c_1251_n 0.00949101f $X=5.585 $Y=0.945 $X2=5.925
+ $Y2=3.165
cc_669 N_A_784_115#_M1001_g N_S_c_1251_n 0.00506137f $X=5.585 $Y=5.085 $X2=5.925
+ $Y2=3.165
cc_670 N_A_784_115#_c_1120_n N_S_c_1251_n 0.0113616f $X=5.415 $Y=3.25 $X2=5.925
+ $Y2=3.165
cc_671 N_A_784_115#_c_1105_n N_S_c_1251_n 0.0246408f $X=5.415 $Y=2.755 $X2=5.925
+ $Y2=3.165
cc_672 N_A_784_115#_c_1106_n N_S_c_1251_n 0.00346737f $X=5.585 $Y=2.755
+ $X2=5.925 $Y2=3.165
cc_673 N_A_784_115#_M1018_g N_S_c_1252_n 0.00698062f $X=5.585 $Y=0.945 $X2=5.925
+ $Y2=2.22
cc_674 N_A_784_115#_M1001_g N_S_c_1254_n 0.00358675f $X=5.585 $Y=5.085 $X2=5.925
+ $Y2=3.25
cc_675 N_A_784_115#_c_1117_n N_S_c_1254_n 0.00477774f $X=5.33 $Y=3.335 $X2=5.925
+ $Y2=3.25
cc_676 N_A_784_115#_c_1120_n N_S_c_1254_n 0.00558264f $X=5.415 $Y=3.25 $X2=5.925
+ $Y2=3.25
cc_677 N_A_784_115#_M1001_g S 0.0118598f $X=5.585 $Y=5.085 $X2=5.8 $Y2=3.365
cc_678 N_A_784_115#_c_1117_n S 0.00549343f $X=5.33 $Y=3.335 $X2=5.8 $Y2=3.365
cc_679 N_A_784_115#_c_1105_n S 0.00428732f $X=5.415 $Y=2.755 $X2=5.8 $Y2=3.365
cc_680 N_A_784_115#_c_1106_n S 0.00105962f $X=5.585 $Y=2.755 $X2=5.8 $Y2=3.365
cc_681 N_A_784_115#_M1001_g N_S_c_1256_n 0.0289488f $X=5.585 $Y=5.085 $X2=5.8
+ $Y2=3.365
cc_682 N_A_784_115#_c_1117_n N_S_c_1256_n 0.00473093f $X=5.33 $Y=3.335 $X2=5.8
+ $Y2=3.365
cc_683 N_A_784_115#_c_1099_n N_A_526_115#_c_1346_n 2.23682e-19 $X=4.06 $Y=0.905
+ $X2=3.63 $Y2=0.825
cc_684 N_S_c_1251_n CO 0.00370359f $X=5.925 $Y=3.165 $X2=6.75 $Y2=2.96
cc_685 N_S_c_1251_n N_CO_c_1300_n 0.0051304f $X=5.925 $Y=3.165 $X2=6.75
+ $Y2=0.825
cc_686 N_S_c_1254_n N_CO_c_1300_n 0.00509957f $X=5.925 $Y=3.25 $X2=6.75
+ $Y2=0.825
