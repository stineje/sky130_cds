* File: sky130_osu_sc_18T_hs__buf_1.pxi.spice
* Created: Fri Nov 12 13:47:48 2021
* 
x_PM_SKY130_OSU_SC_18T_HS__BUF_1%GND N_GND_M1003_d N_GND_M1003_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_HS__BUF_1%GND
x_PM_SKY130_OSU_SC_18T_HS__BUF_1%VDD N_VDD_M1002_d N_VDD_M1002_b N_VDD_c_29_p
+ N_VDD_c_30_p N_VDD_c_39_p VDD N_VDD_c_31_p PM_SKY130_OSU_SC_18T_HS__BUF_1%VDD
x_PM_SKY130_OSU_SC_18T_HS__BUF_1%A N_A_M1003_g N_A_M1002_g N_A_c_54_n N_A_c_55_n
+ A PM_SKY130_OSU_SC_18T_HS__BUF_1%A
x_PM_SKY130_OSU_SC_18T_HS__BUF_1%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1002_s N_A_27_115#_M1001_g N_A_27_115#_c_103_n
+ N_A_27_115#_M1000_g N_A_27_115#_c_92_n N_A_27_115#_c_93_n N_A_27_115#_c_94_n
+ N_A_27_115#_c_95_n N_A_27_115#_c_98_n N_A_27_115#_c_99_n N_A_27_115#_c_101_n
+ N_A_27_115#_c_102_n PM_SKY130_OSU_SC_18T_HS__BUF_1%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__BUF_1%Y N_Y_M1001_d N_Y_M1000_d N_Y_c_144_n
+ N_Y_c_150_n Y N_Y_c_147_n N_Y_c_149_n PM_SKY130_OSU_SC_18T_HS__BUF_1%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1003_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1003_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_A_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.075
cc_5 N_GND_M1003_b N_A_M1002_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_6 N_GND_M1003_b N_A_c_54_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_7 N_GND_M1003_b N_A_c_55_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_8 N_GND_M1003_b N_A_27_115#_M1001_g 0.0337861f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=1.075
cc_9 N_GND_c_3_p N_A_27_115#_M1001_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=1.075
cc_10 N_GND_c_4_p N_A_27_115#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=1.075
cc_11 N_GND_M1003_b N_A_27_115#_c_92_n 0.0597491f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.86
cc_12 N_GND_M1003_b N_A_27_115#_c_93_n 0.0562401f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=1.935
cc_13 N_GND_M1003_b N_A_27_115#_c_94_n 0.0168393f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.935
cc_14 N_GND_M1003_b N_A_27_115#_c_95_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_15 N_GND_c_2_p N_A_27_115#_c_95_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_16 N_GND_c_4_p N_A_27_115#_c_95_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_17 N_GND_M1003_b N_A_27_115#_c_98_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.455
cc_18 N_GND_M1003_b N_A_27_115#_c_99_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.935
cc_19 N_GND_c_3_p N_A_27_115#_c_99_n 0.00702738f $X=0.69 $Y=0.825 $X2=0.88
+ $Y2=1.935
cc_20 N_GND_M1003_b N_A_27_115#_c_101_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.935
cc_21 N_GND_M1003_b N_A_27_115#_c_102_n 0.00663593f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.935
cc_22 N_GND_M1003_b N_Y_c_144_n 0.00892292f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.825
cc_23 N_GND_c_4_p N_Y_c_144_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.12 $Y2=0.825
cc_24 N_GND_M1003_b Y 0.0164841f $X=-0.045 $Y=0 $X2=1.065 $Y2=2.275
cc_25 N_GND_M1003_b N_Y_c_147_n 0.0110015f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.48
cc_26 N_GND_c_3_p N_Y_c_147_n 0.00125659f $X=0.69 $Y=0.825 $X2=1.12 $Y2=1.48
cc_27 N_GND_M1003_b N_Y_c_149_n 0.00501078f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.96
cc_28 N_VDD_M1002_b N_A_M1002_g 0.0245629f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_29 N_VDD_c_29_p N_A_M1002_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475 $Y2=4.585
cc_30 N_VDD_c_30_p N_A_M1002_g 0.00354579f $X=0.69 $Y=4.135 $X2=0.475 $Y2=4.585
cc_31 N_VDD_c_31_p N_A_M1002_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=4.585
cc_32 N_VDD_M1002_d N_A_c_55_n 0.00628533f $X=0.55 $Y=3.085 $X2=0.635 $Y2=2.48
cc_33 N_VDD_M1002_b N_A_c_55_n 0.00328912f $X=-0.045 $Y=2.905 $X2=0.635 $Y2=2.48
cc_34 N_VDD_c_30_p N_A_c_55_n 0.00264661f $X=0.69 $Y=4.135 $X2=0.635 $Y2=2.48
cc_35 N_VDD_M1002_d A 0.00797576f $X=0.55 $Y=3.085 $X2=0.635 $Y2=3.33
cc_36 N_VDD_c_30_p A 0.00510982f $X=0.69 $Y=4.135 $X2=0.635 $Y2=3.33
cc_37 N_VDD_M1002_b N_A_27_115#_c_103_n 0.0194495f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=3.01
cc_38 N_VDD_c_30_p N_A_27_115#_c_103_n 0.00354579f $X=0.69 $Y=4.135 $X2=0.905
+ $Y2=3.01
cc_39 N_VDD_c_39_p N_A_27_115#_c_103_n 0.00606474f $X=1.02 $Y=6.44 $X2=0.905
+ $Y2=3.01
cc_40 N_VDD_c_31_p N_A_27_115#_c_103_n 0.00468827f $X=1.02 $Y=6.47 $X2=0.905
+ $Y2=3.01
cc_41 N_VDD_M1002_b N_A_27_115#_c_94_n 0.0187682f $X=-0.045 $Y=2.905 $X2=1.18
+ $Y2=2.935
cc_42 N_VDD_M1002_b N_A_27_115#_c_98_n 0.00996008f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.455
cc_43 N_VDD_c_29_p N_A_27_115#_c_98_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=3.455
cc_44 N_VDD_c_31_p N_A_27_115#_c_98_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26
+ $Y2=3.455
cc_45 N_VDD_M1002_b N_Y_c_150_n 0.00317324f $X=-0.045 $Y=2.905 $X2=1.12 $Y2=2.96
cc_46 N_VDD_c_39_p N_Y_c_150_n 0.00736239f $X=1.02 $Y=6.44 $X2=1.12 $Y2=2.96
cc_47 N_VDD_c_31_p N_Y_c_150_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.12 $Y2=2.96
cc_48 N_VDD_M1002_b N_Y_c_149_n 0.0107503f $X=-0.045 $Y=2.905 $X2=1.12 $Y2=2.96
cc_49 A N_A_27_115#_M1002_s 0.00414531f $X=0.635 $Y=3.33 $X2=0.135 $Y2=3.085
cc_50 N_A_M1003_g N_A_27_115#_M1001_g 0.0385412f $X=0.475 $Y=1.075 $X2=0.905
+ $Y2=1.075
cc_51 A N_A_27_115#_c_103_n 0.00419145f $X=0.635 $Y=3.33 $X2=0.905 $Y2=3.01
cc_52 N_A_M1003_g N_A_27_115#_c_92_n 0.00260138f $X=0.475 $Y=1.075 $X2=1.18
+ $Y2=2.86
cc_53 N_A_M1002_g N_A_27_115#_c_92_n 0.00209773f $X=0.475 $Y=4.585 $X2=1.18
+ $Y2=2.86
cc_54 N_A_c_54_n N_A_27_115#_c_92_n 0.0139096f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_55 N_A_c_55_n N_A_27_115#_c_92_n 0.00361737f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_56 N_A_M1002_g N_A_27_115#_c_94_n 0.0496795f $X=0.475 $Y=4.585 $X2=1.18
+ $Y2=2.935
cc_57 N_A_c_55_n N_A_27_115#_c_94_n 0.00468272f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.935
cc_58 N_A_M1003_g N_A_27_115#_c_95_n 0.0148408f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_59 N_A_M1003_g N_A_27_115#_c_98_n 0.0337582f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=3.455
cc_60 N_A_c_55_n N_A_27_115#_c_98_n 0.0548951f $X=0.635 $Y=2.48 $X2=0.26
+ $Y2=3.455
cc_61 A N_A_27_115#_c_98_n 0.0155137f $X=0.635 $Y=3.33 $X2=0.26 $Y2=3.455
cc_62 N_A_M1003_g N_A_27_115#_c_99_n 0.0207696f $X=0.475 $Y=1.075 $X2=0.88
+ $Y2=1.935
cc_63 N_A_c_54_n N_A_27_115#_c_99_n 0.00273049f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_64 N_A_c_55_n N_A_27_115#_c_99_n 0.00886797f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_65 N_A_M1003_g N_A_27_115#_c_102_n 6.59135e-19 $X=0.475 $Y=1.075 $X2=0.965
+ $Y2=1.935
cc_66 N_A_c_55_n N_Y_c_150_n 0.0135622f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_67 A N_Y_c_150_n 0.00731851f $X=0.635 $Y=3.33 $X2=1.12 $Y2=2.96
cc_68 N_A_M1003_g Y 0.00310306f $X=0.475 $Y=1.075 $X2=1.065 $Y2=2.275
cc_69 N_A_c_54_n Y 0.00441844f $X=0.635 $Y=2.48 $X2=1.065 $Y2=2.275
cc_70 N_A_c_55_n Y 0.0200396f $X=0.635 $Y=2.48 $X2=1.065 $Y2=2.275
cc_71 N_A_M1003_g N_Y_c_147_n 7.99941e-19 $X=0.475 $Y=1.075 $X2=1.12 $Y2=1.48
cc_72 N_A_c_55_n N_Y_c_149_n 0.00609526f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_73 N_A_27_115#_M1001_g N_Y_c_144_n 0.0057847f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_74 N_A_27_115#_c_93_n N_Y_c_144_n 0.00477112f $X=1.18 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_75 N_A_27_115#_c_102_n N_Y_c_144_n 7.32051e-19 $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_76 N_A_27_115#_c_103_n N_Y_c_150_n 0.00596111f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_77 N_A_27_115#_c_94_n N_Y_c_150_n 0.0134943f $X=1.18 $Y=2.935 $X2=1.12
+ $Y2=2.96
cc_78 N_A_27_115#_M1001_g Y 0.00406656f $X=0.905 $Y=1.075 $X2=1.065 $Y2=2.275
cc_79 N_A_27_115#_c_92_n Y 0.0310322f $X=1.18 $Y=2.86 $X2=1.065 $Y2=2.275
cc_80 N_A_27_115#_c_93_n Y 0.0161039f $X=1.18 $Y=1.935 $X2=1.065 $Y2=2.275
cc_81 N_A_27_115#_c_99_n Y 8.73078e-19 $X=0.88 $Y=1.935 $X2=1.065 $Y2=2.275
cc_82 N_A_27_115#_c_102_n Y 0.0121742f $X=0.965 $Y=1.935 $X2=1.065 $Y2=2.275
cc_83 N_A_27_115#_M1001_g N_Y_c_147_n 0.00668893f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=1.48
cc_84 N_A_27_115#_c_93_n N_Y_c_147_n 0.0014753f $X=1.18 $Y=1.935 $X2=1.12
+ $Y2=1.48
cc_85 N_A_27_115#_c_102_n N_Y_c_147_n 0.00278861f $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=1.48
cc_86 N_A_27_115#_c_103_n N_Y_c_149_n 0.0015856f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_87 N_A_27_115#_c_92_n N_Y_c_149_n 0.00226191f $X=1.18 $Y=2.86 $X2=1.12
+ $Y2=2.96
cc_88 N_A_27_115#_c_94_n N_Y_c_149_n 0.00513726f $X=1.18 $Y=2.935 $X2=1.12
+ $Y2=2.96
