* File: sky130_osu_sc_18T_ls__buf_6.pex.spice
* Created: Fri Nov 12 14:15:03 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_1 1 2 3 4 47 49 56 58 65 67 74 76
+ 83 85 86
r86 81 83 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.825
r87 76 81 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=3.185 $Y=0.152
+ $X2=3.27 $Y2=0.305
r88 72 74 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.825
r89 68 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0.152
+ $X2=1.55 $Y2=0.152
r90 63 86 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.152
r91 63 65 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.825
r92 59 85 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r93 58 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.152
r94 54 85 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r95 54 56 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r96 49 85 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r97 47 72 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.41 $Y2=0.305
r98 47 67 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.325 $Y2=0.152
r99 47 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.495 $Y2=0.152
r100 47 76 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.185 $Y2=0.152
r101 47 77 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.495 $Y2=0.152
r102 47 67 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r103 47 68 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r104 47 58 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r105 47 59 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r106 47 49 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r107 4 83 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.825
r108 3 74 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r109 2 65 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r110 1 56 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_2 1 2 3 4 37 39 45 49 55 59 65 69
+ 75 79 80 82
r60 75 78 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.27 $Y=3.455
+ $X2=3.27 $Y2=5.835
r61 73 78 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=6.355
+ $X2=3.27 $Y2=5.835
r62 70 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=2.41 $Y2=6.507
r63 70 72 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=3.06 $Y2=6.507
r64 69 73 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.27 $Y2=6.355
r65 69 72 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.06 $Y2=6.507
r66 65 68 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r67 63 82 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=6.507
r68 63 68 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=5.835
r69 60 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.55 $Y2=6.507
r70 60 62 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.7 $Y2=6.507
r71 59 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=2.41 $Y2=6.507
r72 59 62 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=1.7 $Y2=6.507
r73 55 58 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r74 53 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=6.507
r75 53 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=5.835
r76 50 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r77 50 52 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r78 49 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.55 $Y2=6.507
r79 49 52 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.02 $Y2=6.507
r80 45 48 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r81 43 79 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r82 43 48 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r83 39 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r84 39 41 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r85 37 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r86 37 82 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r87 37 62 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r88 37 52 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r89 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r90 4 78 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=5.835
r91 4 75 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=3.455
r92 3 68 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r93 3 65 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r94 2 58 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r95 2 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r96 1 48 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r97 1 45 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=3.33
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2.48
+ $X2=0.635 $Y2=3.33
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.48 $X2=0.635 $Y2=2.48
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.645
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.315
r45 7 12 994.766 $w=1.5e-07 $l=1.94e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.645
r46 3 11 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.315
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%A_27_115# 1 3 11 13 15 17 20 22 24 25 26
+ 27 28 31 33 35 36 38 42 44 46 47 49 53 56 57 59 60 62 66 68 70 80 81 82 83 84
+ 85 88 92 96 98 101
c177 57 0 1.33323e-19 $X=2.625 $Y=3.01
c178 53 0 1.33323e-19 $X=2.625 $Y=1.075
c179 44 0 1.33323e-19 $X=2.195 $Y=3.01
c180 42 0 1.33323e-19 $X=2.195 $Y=1.075
c181 33 0 1.33323e-19 $X=1.765 $Y=3.01
c182 31 0 1.33323e-19 $X=1.765 $Y=1.075
c183 22 0 1.33323e-19 $X=1.335 $Y=3.01
c184 20 0 1.33323e-19 $X=1.335 $Y=1.075
r185 97 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.935
+ $X2=0.26 $Y2=1.935
r186 96 101 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.965 $Y2=1.935
r187 96 97 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.345 $Y2=1.935
r188 92 94 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r189 90 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=1.935
r190 90 92 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=3.455
r191 86 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=1.935
r192 86 88 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r193 77 101 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.935 $X2=0.965 $Y2=1.935
r194 77 78 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=1.18 $Y2=1.935
r195 75 77 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.935
+ $X2=0.965 $Y2=1.935
r196 73 74 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.935
+ $X2=1.335 $Y2=2.935
r197 71 73 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.935
+ $X2=1.18 $Y2=2.935
r198 68 70 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.055 $Y=3.01
+ $X2=3.055 $Y2=4.585
r199 64 66 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.075
r200 63 85 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.935 $X2=2.625
+ $Y2=2.935
r201 62 68 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=3.055 $Y2=3.01
r202 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=2.7 $Y2=2.935
r203 61 84 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.845 $X2=2.625
+ $Y2=1.845
r204 60 64 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=3.055 $Y2=1.77
r205 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=2.7 $Y2=1.845
r206 57 85 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=2.935
r207 57 59 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=4.585
r208 56 85 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.86
+ $X2=2.625 $Y2=2.935
r209 55 84 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.92
+ $X2=2.625 $Y2=1.845
r210 55 56 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.625 $Y=1.92 $X2=2.625
+ $Y2=2.86
r211 51 84 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.845
r212 51 53 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.075
r213 50 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.935
+ $X2=2.195 $Y2=2.935
r214 49 85 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.625 $Y2=2.935
r215 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.27 $Y2=2.935
r216 48 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.195 $Y2=1.845
r217 47 84 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.625 $Y2=1.845
r218 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.27 $Y2=1.845
r219 44 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=2.935
r220 44 46 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=4.585
r221 40 82 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.845
r222 40 42 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r223 39 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.935
+ $X2=1.765 $Y2=2.935
r224 38 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=2.195 $Y2=2.935
r225 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=1.84 $Y2=2.935
r226 37 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.765 $Y2=1.845
r227 36 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.845
r228 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r229 33 81 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=2.935
r230 33 35 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=4.585
r231 29 80 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.845
r232 29 31 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r233 28 74 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.935
+ $X2=1.335 $Y2=2.935
r234 27 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.765 $Y2=2.935
r235 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.41 $Y2=2.935
r236 25 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.765 $Y2=1.845
r237 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.41 $Y2=1.845
r238 22 74 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=2.935
r239 22 24 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=4.585
r240 18 26 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.41 $Y2=1.845
r241 18 78 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.18 $Y2=1.935
r242 18 20 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r243 17 73 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.86
+ $X2=1.18 $Y2=2.935
r244 16 78 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=1.935
r245 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=2.86
r246 13 71 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=2.935
r247 13 15 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=4.585
r248 9 75 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.935
r249 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.075
r250 3 94 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r251 3 92 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r252 1 88 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%Y 1 2 3 7 8 9 26 32 40 46 54 60 67 68 70
+ 72 74 77 78 79 80 81 82 83
c124 83 0 1.33323e-19 $X=2.84 $Y=2.845
c125 82 0 1.33323e-19 $X=2.84 $Y=1.595
c126 81 0 2.66647e-19 $X=2.125 $Y=2.96
c127 79 0 2.66647e-19 $X=2.125 $Y=1.48
c128 68 0 1.33323e-19 $X=1.12 $Y=2.845
c129 67 0 1.33323e-19 $X=1.12 $Y=1.595
r130 83 95 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=2.845
+ $X2=2.84 $Y2=2.96
r131 82 93 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=1.48
r132 82 83 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=2.845
r133 81 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=2.96
+ $X2=1.98 $Y2=2.96
r134 80 95 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.84 $Y2=2.96
r135 80 81 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.125 $Y2=2.96
r136 79 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=1.48
+ $X2=1.98 $Y2=1.48
r137 78 93 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.84 $Y2=1.48
r138 78 79 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.125 $Y2=1.48
r139 77 91 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.845
+ $X2=1.98 $Y2=2.96
r140 76 89 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=1.48
r141 76 77 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=2.845
r142 75 87 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.96
+ $X2=1.12 $Y2=2.96
r143 74 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.98 $Y2=2.96
r144 74 75 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.265 $Y2=2.96
r145 73 85 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1.48
+ $X2=1.12 $Y2=1.48
r146 72 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.98 $Y2=1.48
r147 72 73 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.265 $Y2=1.48
r148 68 87 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.96
r149 68 70 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.27
r150 67 85 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=1.48
r151 67 70 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=2.27
r152 63 65 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r153 60 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=2.96
r154 60 63 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=3.455
r155 57 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=1.48
+ $X2=2.84 $Y2=1.48
r156 54 57 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.84 $Y=0.825
+ $X2=2.84 $Y2=1.48
r157 49 51 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r158 46 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=2.96
r159 46 49 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=3.455
r160 43 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=1.48
r161 40 43 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.98 $Y=0.825
+ $X2=1.98 $Y2=1.48
r162 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r163 32 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=2.96
r164 32 35 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=3.455
r165 29 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=1.48
r166 26 29 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.12 $Y=0.825
+ $X2=1.12 $Y2=1.48
r167 9 65 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r168 9 63 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r169 8 51 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r170 8 49 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r171 7 37 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r172 7 35 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r173 3 54 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r174 2 40 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r175 1 26 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
.ends

