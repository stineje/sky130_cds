* File: sky130_osu_sc_18T_ls__buf_4.spice
* Created: Fri Nov 12 14:14:55 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_ls__buf_4.pex.spice"
.subckt sky130_osu_sc_18T_ls__buf_4  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1004_d N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1000_d N_A_27_115#_M1001_g N_GND_M1001_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_A_27_115#_M1007_g N_GND_M1001_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1007_d N_A_27_115#_M1008_g N_GND_M1008_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g N_A_27_115#_M1003_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1002 N_Y_M1002_d N_A_27_115#_M1002_g N_VDD_M1003_d N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75001.5 A=0.45 P=6.3 MULT=1
MM1005 N_Y_M1002_d N_A_27_115#_M1005_g N_VDD_M1005_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1006 N_Y_M1006_d N_A_27_115#_M1006_g N_VDD_M1005_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.5
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1009 N_Y_M1006_d N_A_27_115#_M1009_g N_VDD_M1009_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75001.9
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX10_noxref N_GND_M1004_b N_VDD_M1003_b NWDIODE A=10.659 P=13.21
pX11_noxref noxref_6 A A PROBETYPE=1
pX12_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__buf_4.pxi.spice"
*
.ends
*
*
