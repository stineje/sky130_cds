* File: sky130_osu_sc_15T_ms__and2_2.spice
* Created: Fri Nov 12 14:40:11 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__and2_2.pex.spice"
.subckt sky130_osu_sc_15T_ms__and2_2  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1005 A_110_115# N_A_M1005_g N_A_27_115#_M1005_s N_GND_M1005_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1002 N_GND_M1002_d N_B_M1002_g A_110_115# N_GND_M1005_b NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.0777 PD=1.09 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1005_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1001_d N_A_27_115#_M1007_g N_GND_M1007_s N_GND_M1005_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_115#_M1006_d N_A_M1006_g N_VDD_M1006_s N_VDD_M1006_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001.5 A=0.3 P=4.3 MULT=1
MM1003 N_VDD_M1003_d N_B_M1003_g N_A_27_115#_M1006_d N_VDD_M1006_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1000 N_VDD_M1003_d N_A_27_115#_M1000_g N_Y_M1000_s N_VDD_M1006_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1004 N_VDD_M1004_d N_A_27_115#_M1004_g N_Y_M1000_s N_VDD_M1006_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001.5
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX8_noxref N_GND_M1005_b N_VDD_M1006_b NWDIODE A=6.94725 P=10.61
pX9_noxref noxref_8 A A PROBETYPE=1
pX10_noxref noxref_9 B B PROBETYPE=1
pX11_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__and2_2.pxi.spice"
*
.ends
*
*
