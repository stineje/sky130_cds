* File: sky130_osu_sc_12T_ms__aoi21_l.pex.spice
* Created: Fri Nov 12 15:21:12 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%GND 1 2 21 25 27 35 42 45
c45 21 0 6.36774e-20 $X=-0.05 $Y=0
r46 42 45 0.321969 $w=3e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.15 $X2=1.02
+ $Y2=0.15
r47 33 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.54 $Y=0.3
+ $X2=1.54 $Y2=0.735
r48 27 33 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.455 $Y=0.15
+ $X2=1.54 $Y2=0.3
r49 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.3
+ $X2=0.26 $Y2=0.735
r50 21 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.185
+ $X2=1.02 $Y2=0.185
r51 21 23 4.3533 $w=1.7e-07 $l=1.88944e-07 $layer=LI1_cond $X=0.172 $Y=0.15
+ $X2=0.26 $Y2=0.3
r52 21 28 3.16437 $w=3e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.15
+ $X2=0.345 $Y2=0.15
r53 21 27 16.7104 $w=2.98e-07 $l=4.35e-07 $layer=LI1_cond $X=1.02 $Y=0.15
+ $X2=1.455 $Y2=0.15
r54 21 28 25.93 $w=2.98e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.15
+ $X2=0.345 $Y2=0.15
r55 2 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.57 $X2=1.54 $Y2=0.735
r56 1 25 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.57 $X2=0.26 $Y2=0.735
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%VDD 1 13 15 21 25 29 32
r26 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r27 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r28 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r29 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287 $X2=1.02
+ $Y2=4.287
r30 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r31 19 21 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.63
r32 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r33 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r34 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r35 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r36 1 21 600 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.63
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%A0 2 3 5 8 12 18 21 27
c34 8 0 6.36774e-20 $X=0.475 $Y=3.235
r35 21 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=2.11
+ $X2=0.385 $Y2=2.11
r36 21 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.385 $Y=2.11
+ $X2=0.385 $Y2=2.285
r37 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.285 $X2=0.385 $Y2=2.285
r38 17 18 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.285
+ $X2=0.475 $Y2=2.285
r39 14 17 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.285
+ $X2=0.385 $Y2=2.285
r40 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.29
+ $X2=0.475 $Y2=1.29
r41 6 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.42
+ $X2=0.475 $Y2=2.285
r42 6 8 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=0.475 $Y=2.42
+ $X2=0.475 $Y2=3.235
r43 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.21 $X2=0.475
+ $Y2=1.29
r44 3 5 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=0.83
r45 2 14 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.15
+ $X2=0.295 $Y2=2.285
r46 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.37 $X2=0.295
+ $Y2=1.29
r47 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.37
+ $X2=0.295 $Y2=2.15
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%A1 3 7 10 15 20 23
c51 23 0 1.59493e-19 $X=0.725 $Y=2.48
r52 17 20 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.725 $Y=1.775
+ $X2=0.815 $Y2=1.775
r53 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.48
+ $X2=0.725 $Y2=2.48
r54 13 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.94
+ $X2=0.725 $Y2=1.775
r55 13 15 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.725 $Y=1.94
+ $X2=0.725 $Y2=2.48
r56 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=1.775 $X2=0.815 $Y2=1.775
r57 10 12 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.775
+ $X2=0.825 $Y2=1.94
r58 10 11 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.775
+ $X2=0.825 $Y2=1.61
r59 7 12 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=1.94
r60 3 11 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.835 $Y=0.83
+ $X2=0.835 $Y2=1.61
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%B0 3 5 7 9 12 15 20 22 24 27
c55 9 0 2.08793e-20 $X=1.47 $Y=2.37
c56 5 0 1.38614e-19 $X=1.335 $Y=2.52
r57 22 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.25 $Y=1.38
+ $X2=1.53 $Y2=1.38
r58 20 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.11
+ $X2=1.165 $Y2=2.11
r59 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.165 $Y=1.465
+ $X2=1.25 $Y2=1.38
r60 18 20 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.165 $Y=1.465
+ $X2=1.165 $Y2=2.11
r61 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.53
+ $Y=1.38 $X2=1.53 $Y2=1.38
r62 15 17 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.47 $Y=1.38 $X2=1.53
+ $Y2=1.38
r63 10 12 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.335 $Y=2.445
+ $X2=1.47 $Y2=2.445
r64 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=2.37 $X2=1.47
+ $Y2=2.445
r65 8 15 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=1.545
+ $X2=1.47 $Y2=1.38
r66 8 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=1.47 $Y=1.545
+ $X2=1.47 $Y2=2.37
r67 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.52
+ $X2=1.335 $Y2=2.445
r68 5 7 229.753 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.335 $Y=2.52
+ $X2=1.335 $Y2=3.235
r69 1 15 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.325 $Y=1.215
+ $X2=1.47 $Y2=1.38
r70 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.325 $Y=1.215
+ $X2=1.325 $Y2=0.75
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%A_27_521# 1 2 11 13 14 17
r15 15 17 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.12 $Y=3.23
+ $X2=1.12 $Y2=3.635
r16 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.145
+ $X2=1.12 $Y2=3.23
r17 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.145
+ $X2=0.345 $Y2=3.145
r18 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.23
+ $X2=0.345 $Y2=3.145
r19 9 11 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.26 $Y=3.23 $X2=0.26
+ $Y2=3.63
r20 2 17 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r21 1 11 600 $w=1.7e-07 $l=1.0857e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.63
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AOI21_L%Y 1 3 10 16 21 26 31 33
r50 29 31 0.0825816 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=1.05 $Y=1
+ $X2=1.165 $Y2=1
r51 24 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.625
+ $X2=1.55 $Y2=1.74
r52 24 26 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.55 $Y=1.625
+ $X2=1.55 $Y2=1.59
r53 23 26 0.481441 $w=1.7e-07 $l=5e-07 $layer=MET1_cond $X=1.55 $Y=1.09 $X2=1.55
+ $Y2=1.59
r54 21 23 0.0698602 $w=1.75e-07 $l=1.23386e-07 $layer=MET1_cond $X=1.465
+ $Y=1.002 $X2=1.55 $Y2=1.09
r55 21 31 0.271526 $w=1.75e-07 $l=3e-07 $layer=MET1_cond $X=1.465 $Y=1.002
+ $X2=1.165 $Y2=1.002
r56 16 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.74
+ $X2=1.55 $Y2=1.74
r57 16 19 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=1.55 $Y=1.74
+ $X2=1.55 $Y2=3.33
r58 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.05 $Y=1 $X2=1.05
+ $Y2=1
r59 10 13 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.05 $Y=0.735
+ $X2=1.05 $Y2=1
r60 3 19 300 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.33
r61 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.57 $X2=1.05 $Y2=0.735
.ends

