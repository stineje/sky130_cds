magic
tech sky130A
magscale 1 2
timestamp 1606864622
<< checkpaint >>
rect -1209 -1243 1753 2575
<< nwell >>
rect -9 581 638 1341
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 238 617 268 1217
rect 358 617 388 1217
rect 430 617 460 1217
rect 516 617 546 1217
<< nmoslvt >>
rect 80 115 110 315
rect 166 115 196 315
rect 238 115 268 315
rect 358 115 388 315
rect 430 115 460 315
rect 516 115 546 315
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 166 315
rect 110 131 121 267
rect 155 131 166 267
rect 110 115 166 131
rect 196 115 238 315
rect 268 267 358 315
rect 268 131 279 267
rect 347 131 358 267
rect 268 115 358 131
rect 388 115 430 315
rect 460 267 516 315
rect 460 131 471 267
rect 505 131 516 267
rect 460 115 516 131
rect 546 267 599 315
rect 546 131 557 267
rect 591 131 599 267
rect 546 115 599 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 657 35 1201
rect 69 657 80 1201
rect 27 617 80 657
rect 110 1201 166 1217
rect 110 793 121 1201
rect 155 793 166 1201
rect 110 617 166 793
rect 196 617 238 1217
rect 268 1201 358 1217
rect 268 657 279 1201
rect 347 657 358 1201
rect 268 617 358 657
rect 388 617 430 1217
rect 460 1201 516 1217
rect 460 793 471 1201
rect 505 793 516 1201
rect 460 617 516 793
rect 546 1201 599 1217
rect 546 658 557 1201
rect 591 658 599 1201
rect 546 617 599 658
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 279 131 347 267
rect 471 131 505 267
rect 557 131 591 267
<< pdiffc >>
rect 35 657 69 1201
rect 121 793 155 1201
rect 279 657 347 1201
rect 471 793 505 1201
rect 557 658 591 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 238 1217 268 1243
rect 358 1217 388 1243
rect 430 1217 460 1243
rect 516 1217 546 1243
rect 80 602 110 617
rect 166 602 196 617
rect 70 572 196 602
rect 70 355 100 572
rect 142 570 196 572
rect 142 536 152 570
rect 186 536 196 570
rect 142 520 196 536
rect 142 462 196 478
rect 142 428 152 462
rect 186 428 196 462
rect 142 412 196 428
rect 70 330 110 355
rect 80 315 110 330
rect 166 315 196 412
rect 238 403 268 617
rect 358 586 388 617
rect 334 570 388 586
rect 430 602 460 617
rect 516 602 546 617
rect 430 572 546 602
rect 334 536 344 570
rect 378 536 388 570
rect 334 520 388 536
rect 479 570 546 572
rect 479 536 489 570
rect 523 536 546 570
rect 479 520 546 536
rect 420 461 474 477
rect 420 432 430 461
rect 358 427 430 432
rect 464 427 474 461
rect 238 387 292 403
rect 238 353 248 387
rect 282 353 292 387
rect 238 337 292 353
rect 358 402 474 427
rect 238 315 268 337
rect 358 315 388 402
rect 516 360 546 520
rect 430 330 546 360
rect 430 315 460 330
rect 516 315 546 330
rect 80 89 110 115
rect 166 89 196 115
rect 238 89 268 115
rect 358 89 388 115
rect 430 89 460 115
rect 516 89 546 115
<< polycont >>
rect 152 536 186 570
rect 152 428 186 462
rect 344 536 378 570
rect 489 536 523 570
rect 430 427 464 461
rect 248 353 282 387
<< locali >>
rect 0 1311 638 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 638 1311
rect 35 1201 69 1217
rect 121 1201 155 1271
rect 121 777 155 793
rect 279 1201 347 1217
rect 35 462 69 657
rect 152 649 200 683
rect 268 657 279 675
rect 471 1201 505 1271
rect 471 777 505 793
rect 557 1201 591 1217
rect 152 570 186 649
rect 268 641 347 657
rect 136 536 152 570
rect 186 536 202 570
rect 268 535 302 641
rect 344 570 378 586
rect 344 462 378 536
rect 35 428 152 462
rect 186 428 378 462
rect 412 461 446 649
rect 489 570 523 575
rect 489 520 523 536
rect 35 267 69 428
rect 412 427 430 461
rect 464 427 480 461
rect 557 387 591 658
rect 232 353 248 387
rect 282 353 591 387
rect 35 115 69 131
rect 121 267 155 283
rect 121 61 155 131
rect 279 279 296 283
rect 330 279 347 283
rect 279 267 347 279
rect 279 115 347 131
rect 471 267 505 283
rect 471 61 505 131
rect 557 267 591 353
rect 557 115 591 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 638 61
rect 0 0 638 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 200 649 234 683
rect 412 649 446 683
rect 268 501 302 535
rect 489 575 523 609
rect 296 279 330 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1311 638 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 638 1311
rect 0 1271 638 1277
rect 188 683 246 689
rect 400 683 458 689
rect 188 649 200 683
rect 234 649 412 683
rect 446 649 458 683
rect 188 643 246 649
rect 400 643 458 649
rect 477 609 535 615
rect 455 575 489 609
rect 523 575 535 609
rect 477 569 535 575
rect 256 535 314 541
rect 256 501 268 535
rect 302 501 314 535
rect 256 495 314 501
rect 268 319 302 495
rect 268 313 342 319
rect 268 279 296 313
rect 330 279 342 313
rect 284 273 342 279
rect 0 55 638 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 638 55
rect 0 0 638 21
<< labels >>
rlabel metal1 218 666 218 666 1 A
port 1 n
rlabel metal1 285 486 285 486 1 Y
port 2 n
rlabel metal1 506 592 506 592 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
