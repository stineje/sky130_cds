* File: sky130_osu_sc_15T_hs__or2_8.pxi.spice
* Created: Fri Nov 12 14:32:56 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__OR2_8%GND N_GND_M1007_s N_GND_M1002_d N_GND_M1008_s
+ N_GND_M1013_s N_GND_M1015_s N_GND_M1017_s N_GND_M1007_b N_GND_c_2_p
+ N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p N_GND_c_24_p N_GND_c_32_p N_GND_c_38_p
+ N_GND_c_45_p N_GND_c_52_p N_GND_c_59_p N_GND_c_65_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_15T_HS__OR2_8%GND
x_PM_SKY130_OSU_SC_15T_HS__OR2_8%VDD N_VDD_M1005_d N_VDD_M1001_d N_VDD_M1006_d
+ N_VDD_M1012_d N_VDD_M1019_d N_VDD_M1010_b N_VDD_c_140_p N_VDD_c_146_p
+ N_VDD_c_153_p N_VDD_c_159_p N_VDD_c_165_p N_VDD_c_170_p N_VDD_c_176_p
+ N_VDD_c_181_p N_VDD_c_187_p N_VDD_c_192_p VDD N_VDD_c_141_p
+ PM_SKY130_OSU_SC_15T_HS__OR2_8%VDD
x_PM_SKY130_OSU_SC_15T_HS__OR2_8%B N_B_M1007_g N_B_M1010_g N_B_c_225_n
+ N_B_c_226_n B PM_SKY130_OSU_SC_15T_HS__OR2_8%B
x_PM_SKY130_OSU_SC_15T_HS__OR2_8%A N_A_M1002_g N_A_M1005_g N_A_c_253_n
+ N_A_c_254_n A PM_SKY130_OSU_SC_15T_HS__OR2_8%A
x_PM_SKY130_OSU_SC_15T_HS__OR2_8%A_27_565# N_A_27_565#_M1007_d
+ N_A_27_565#_M1010_s N_A_27_565#_M1004_g N_A_27_565#_c_362_n
+ N_A_27_565#_M1000_g N_A_27_565#_c_296_n N_A_27_565#_c_297_n
+ N_A_27_565#_M1008_g N_A_27_565#_c_367_n N_A_27_565#_M1001_g
+ N_A_27_565#_c_302_n N_A_27_565#_c_304_n N_A_27_565#_c_305_n
+ N_A_27_565#_M1009_g N_A_27_565#_c_374_n N_A_27_565#_M1003_g
+ N_A_27_565#_c_310_n N_A_27_565#_c_311_n N_A_27_565#_M1013_g
+ N_A_27_565#_c_379_n N_A_27_565#_M1006_g N_A_27_565#_c_316_n
+ N_A_27_565#_c_318_n N_A_27_565#_M1014_g N_A_27_565#_c_323_n
+ N_A_27_565#_c_385_n N_A_27_565#_M1011_g N_A_27_565#_c_324_n
+ N_A_27_565#_c_325_n N_A_27_565#_M1015_g N_A_27_565#_c_390_n
+ N_A_27_565#_M1012_g N_A_27_565#_c_330_n N_A_27_565#_c_332_n
+ N_A_27_565#_M1016_g N_A_27_565#_c_396_n N_A_27_565#_M1018_g
+ N_A_27_565#_c_337_n N_A_27_565#_c_338_n N_A_27_565#_M1017_g
+ N_A_27_565#_c_401_n N_A_27_565#_M1019_g N_A_27_565#_c_343_n
+ N_A_27_565#_c_344_n N_A_27_565#_c_345_n N_A_27_565#_c_346_n
+ N_A_27_565#_c_347_n N_A_27_565#_c_348_n N_A_27_565#_c_349_n
+ N_A_27_565#_c_350_n N_A_27_565#_c_351_n N_A_27_565#_c_352_n
+ N_A_27_565#_c_353_n N_A_27_565#_c_354_n N_A_27_565#_c_412_n
+ N_A_27_565#_c_416_n N_A_27_565#_c_418_n N_A_27_565#_c_355_n
+ N_A_27_565#_c_356_n N_A_27_565#_c_359_n N_A_27_565#_c_361_n
+ PM_SKY130_OSU_SC_15T_HS__OR2_8%A_27_565#
x_PM_SKY130_OSU_SC_15T_HS__OR2_8%Y N_Y_M1004_d N_Y_M1009_d N_Y_M1014_d
+ N_Y_M1016_d N_Y_M1000_s N_Y_M1003_s N_Y_M1011_s N_Y_M1018_s N_Y_c_538_n
+ N_Y_c_542_n N_Y_c_543_n N_Y_c_548_n N_Y_c_549_n N_Y_c_554_n N_Y_c_555_n
+ N_Y_c_559_n N_Y_c_560_n N_Y_c_563_n Y N_Y_c_565_n N_Y_c_568_n N_Y_c_569_n
+ N_Y_c_570_n N_Y_c_573_n N_Y_c_576_n N_Y_c_577_n N_Y_c_578_n N_Y_c_581_n
+ N_Y_c_582_n N_Y_c_583_n N_Y_c_584_n N_Y_c_587_n N_Y_c_588_n
+ PM_SKY130_OSU_SC_15T_HS__OR2_8%Y
cc_1 N_GND_M1007_b N_B_M1007_g 0.0919998f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_B_M1007_g 0.00866533f $X=0.26 $Y=0.865 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_B_M1007_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.895
cc_4 N_GND_c_4_p N_B_M1007_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.475 $Y2=0.895
cc_5 N_GND_M1007_b N_B_M1010_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_6 N_GND_M1007_b N_B_c_225_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.415
cc_7 N_GND_M1007_b N_B_c_226_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.415
cc_8 N_GND_M1007_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.7
cc_9 N_GND_M1007_b N_A_M1002_g 0.0494465f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.895
cc_10 N_GND_c_3_p N_A_M1002_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.895
cc_11 N_GND_c_11_p N_A_M1002_g 0.00388248f $X=1.12 $Y=0.865 $X2=0.905 $Y2=0.895
cc_12 N_GND_c_4_p N_A_M1002_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.905 $Y2=0.895
cc_13 N_GND_M1007_b N_A_M1005_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_14 N_GND_M1007_b N_A_c_253_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.125
cc_15 N_GND_M1007_b N_A_c_254_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.125
cc_16 N_GND_M1007_b N_A_27_565#_M1004_g 0.0255964f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.895
cc_17 N_GND_c_11_p N_A_27_565#_M1004_g 0.00388248f $X=1.12 $Y=0.865 $X2=1.335
+ $Y2=0.895
cc_18 N_GND_c_18_p N_A_27_565#_M1004_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.895
cc_19 N_GND_c_4_p N_A_27_565#_M1004_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.335
+ $Y2=0.895
cc_20 N_GND_M1007_b N_A_27_565#_c_296_n 0.0466273f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.55
cc_21 N_GND_M1007_b N_A_27_565#_c_297_n 0.00727817f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.625
cc_22 N_GND_M1007_b N_A_27_565#_M1008_g 0.0245289f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.895
cc_23 N_GND_c_18_p N_A_27_565#_M1008_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.895
cc_24 N_GND_c_24_p N_A_27_565#_M1008_g 0.00390533f $X=1.98 $Y=0.865 $X2=1.765
+ $Y2=0.895
cc_25 N_GND_c_4_p N_A_27_565#_M1008_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.765
+ $Y2=0.895
cc_26 N_GND_M1007_b N_A_27_565#_c_302_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_27 N_GND_c_24_p N_A_27_565#_c_302_n 0.00256938f $X=1.98 $Y=0.865 $X2=2.12
+ $Y2=1.585
cc_28 N_GND_M1007_b N_A_27_565#_c_304_n 0.0447518f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.585
cc_29 N_GND_M1007_b N_A_27_565#_c_305_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.625
cc_30 N_GND_M1007_b N_A_27_565#_M1009_g 0.0245289f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.895
cc_31 N_GND_c_24_p N_A_27_565#_M1009_g 0.00390533f $X=1.98 $Y=0.865 $X2=2.195
+ $Y2=0.895
cc_32 N_GND_c_32_p N_A_27_565#_M1009_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.895
cc_33 N_GND_c_4_p N_A_27_565#_M1009_g 0.00468827f $X=4.42 $Y=0.19 $X2=2.195
+ $Y2=0.895
cc_34 N_GND_M1007_b N_A_27_565#_c_310_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.585
cc_35 N_GND_M1007_b N_A_27_565#_c_311_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.625
cc_36 N_GND_M1007_b N_A_27_565#_M1013_g 0.0245289f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.895
cc_37 N_GND_c_32_p N_A_27_565#_M1013_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.895
cc_38 N_GND_c_38_p N_A_27_565#_M1013_g 0.00390533f $X=2.84 $Y=0.865 $X2=2.625
+ $Y2=0.895
cc_39 N_GND_c_4_p N_A_27_565#_M1013_g 0.00468827f $X=4.42 $Y=0.19 $X2=2.625
+ $Y2=0.895
cc_40 N_GND_M1007_b N_A_27_565#_c_316_n 0.0181078f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.585
cc_41 N_GND_c_38_p N_A_27_565#_c_316_n 0.00256938f $X=2.84 $Y=0.865 $X2=2.98
+ $Y2=1.585
cc_42 N_GND_M1007_b N_A_27_565#_c_318_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.625
cc_43 N_GND_M1007_b N_A_27_565#_M1014_g 0.0245289f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.895
cc_44 N_GND_c_38_p N_A_27_565#_M1014_g 0.00390533f $X=2.84 $Y=0.865 $X2=3.055
+ $Y2=0.895
cc_45 N_GND_c_45_p N_A_27_565#_M1014_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.055
+ $Y2=0.895
cc_46 N_GND_c_4_p N_A_27_565#_M1014_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.055
+ $Y2=0.895
cc_47 N_GND_M1007_b N_A_27_565#_c_323_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.55
cc_48 N_GND_M1007_b N_A_27_565#_c_324_n 0.0180386f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.585
cc_49 N_GND_M1007_b N_A_27_565#_c_325_n 0.0118833f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.625
cc_50 N_GND_M1007_b N_A_27_565#_M1015_g 0.0245289f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=0.895
cc_51 N_GND_c_45_p N_A_27_565#_M1015_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.485
+ $Y2=0.895
cc_52 N_GND_c_52_p N_A_27_565#_M1015_g 0.00390533f $X=3.7 $Y=0.865 $X2=3.485
+ $Y2=0.895
cc_53 N_GND_c_4_p N_A_27_565#_M1015_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.485
+ $Y2=0.895
cc_54 N_GND_M1007_b N_A_27_565#_c_330_n 0.0181078f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.585
cc_55 N_GND_c_52_p N_A_27_565#_c_330_n 0.00256938f $X=3.7 $Y=0.865 $X2=3.84
+ $Y2=1.585
cc_56 N_GND_M1007_b N_A_27_565#_c_332_n 0.013058f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.625
cc_57 N_GND_M1007_b N_A_27_565#_M1016_g 0.0245289f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=0.895
cc_58 N_GND_c_52_p N_A_27_565#_M1016_g 0.00390533f $X=3.7 $Y=0.865 $X2=3.915
+ $Y2=0.895
cc_59 N_GND_c_59_p N_A_27_565#_M1016_g 0.00606474f $X=4.475 $Y=0.152 $X2=3.915
+ $Y2=0.895
cc_60 N_GND_c_4_p N_A_27_565#_M1016_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.915
+ $Y2=0.895
cc_61 N_GND_M1007_b N_A_27_565#_c_337_n 0.0369419f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=1.585
cc_62 N_GND_M1007_b N_A_27_565#_c_338_n 0.0268552f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=2.625
cc_63 N_GND_M1007_b N_A_27_565#_M1017_g 0.0341369f $X=-0.045 $Y=0 $X2=4.345
+ $Y2=0.895
cc_64 N_GND_c_59_p N_A_27_565#_M1017_g 0.00606474f $X=4.475 $Y=0.152 $X2=4.345
+ $Y2=0.895
cc_65 N_GND_c_65_p N_A_27_565#_M1017_g 0.00866533f $X=4.56 $Y=0.865 $X2=4.345
+ $Y2=0.895
cc_66 N_GND_c_4_p N_A_27_565#_M1017_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.345
+ $Y2=0.895
cc_67 N_GND_M1007_b N_A_27_565#_c_343_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.625
cc_68 N_GND_M1007_b N_A_27_565#_c_344_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.625
cc_69 N_GND_M1007_b N_A_27_565#_c_345_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.585
cc_70 N_GND_M1007_b N_A_27_565#_c_346_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.625
cc_71 N_GND_M1007_b N_A_27_565#_c_347_n 0.00873941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.585
cc_72 N_GND_M1007_b N_A_27_565#_c_348_n 0.00735657f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.625
cc_73 N_GND_M1007_b N_A_27_565#_c_349_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.585
cc_74 N_GND_M1007_b N_A_27_565#_c_350_n 0.00151234f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.625
cc_75 N_GND_M1007_b N_A_27_565#_c_351_n 0.00873941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.585
cc_76 N_GND_M1007_b N_A_27_565#_c_352_n 0.00735657f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.625
cc_77 N_GND_M1007_b N_A_27_565#_c_353_n 0.00873941f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=1.585
cc_78 N_GND_M1007_b N_A_27_565#_c_354_n 0.00735657f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=2.625
cc_79 N_GND_M1007_b N_A_27_565#_c_355_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.285
cc_80 N_GND_M1007_b N_A_27_565#_c_356_n 0.00953944f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.865
cc_81 N_GND_c_3_p N_A_27_565#_c_356_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.865
cc_82 N_GND_c_4_p N_A_27_565#_c_356_n 0.00475776f $X=4.42 $Y=0.19 $X2=0.69
+ $Y2=0.865
cc_83 N_GND_M1007_b N_A_27_565#_c_359_n 0.0190355f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_84 N_GND_c_11_p N_A_27_565#_c_359_n 0.00702738f $X=1.12 $Y=0.865 $X2=1.43
+ $Y2=1.675
cc_85 N_GND_M1007_b N_A_27_565#_c_361_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.675
cc_86 N_GND_M1007_b N_Y_c_538_n 0.00558158f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.865
cc_87 N_GND_c_18_p N_Y_c_538_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.865
cc_88 N_GND_c_24_p N_Y_c_538_n 8.14297e-19 $X=1.98 $Y=0.865 $X2=1.55 $Y2=0.865
cc_89 N_GND_c_4_p N_Y_c_538_n 0.00475776f $X=4.42 $Y=0.19 $X2=1.55 $Y2=0.865
cc_90 N_GND_M1007_b N_Y_c_542_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_91 N_GND_M1007_b N_Y_c_543_n 0.00656459f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.865
cc_92 N_GND_c_24_p N_Y_c_543_n 8.14297e-19 $X=1.98 $Y=0.865 $X2=2.41 $Y2=0.865
cc_93 N_GND_c_32_p N_Y_c_543_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.865
cc_94 N_GND_c_38_p N_Y_c_543_n 8.14297e-19 $X=2.84 $Y=0.865 $X2=2.41 $Y2=0.865
cc_95 N_GND_c_4_p N_Y_c_543_n 0.00475776f $X=4.42 $Y=0.19 $X2=2.41 $Y2=0.865
cc_96 N_GND_M1007_b N_Y_c_548_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.33
cc_97 N_GND_M1007_b N_Y_c_549_n 0.00656459f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.865
cc_98 N_GND_c_38_p N_Y_c_549_n 8.14297e-19 $X=2.84 $Y=0.865 $X2=3.27 $Y2=0.865
cc_99 N_GND_c_45_p N_Y_c_549_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.865
cc_100 N_GND_c_52_p N_Y_c_549_n 8.14297e-19 $X=3.7 $Y=0.865 $X2=3.27 $Y2=0.865
cc_101 N_GND_c_4_p N_Y_c_549_n 0.00475776f $X=4.42 $Y=0.19 $X2=3.27 $Y2=0.865
cc_102 N_GND_M1007_b N_Y_c_554_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.33
cc_103 N_GND_M1007_b N_Y_c_555_n 0.00656459f $X=-0.045 $Y=0 $X2=4.13 $Y2=0.865
cc_104 N_GND_c_52_p N_Y_c_555_n 8.14297e-19 $X=3.7 $Y=0.865 $X2=4.13 $Y2=0.865
cc_105 N_GND_c_59_p N_Y_c_555_n 0.0075556f $X=4.475 $Y=0.152 $X2=4.13 $Y2=0.865
cc_106 N_GND_c_4_p N_Y_c_555_n 0.00475776f $X=4.42 $Y=0.19 $X2=4.13 $Y2=0.865
cc_107 N_GND_M1007_b N_Y_c_559_n 0.0152877f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.33
cc_108 N_GND_M1007_b N_Y_c_560_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.335
cc_109 N_GND_c_11_p N_Y_c_560_n 0.00134236f $X=1.12 $Y=0.865 $X2=1.55 $Y2=1.335
cc_110 N_GND_c_24_p N_Y_c_560_n 7.53951e-19 $X=1.98 $Y=0.865 $X2=1.55 $Y2=1.335
cc_111 N_GND_M1007_b N_Y_c_563_n 0.00509006f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.215
cc_112 N_GND_M1007_b Y 0.0305055f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.96
cc_113 N_GND_M1008_s N_Y_c_565_n 0.00418405f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.22
cc_114 N_GND_M1007_b N_Y_c_565_n 0.00793787f $X=-0.045 $Y=0 $X2=2.265 $Y2=1.22
cc_115 N_GND_c_24_p N_Y_c_565_n 0.0142303f $X=1.98 $Y=0.865 $X2=2.265 $Y2=1.22
cc_116 N_GND_M1007_b N_Y_c_568_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.33
cc_117 N_GND_M1007_b N_Y_c_569_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.215
cc_118 N_GND_M1013_s N_Y_c_570_n 0.00418405f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.22
cc_119 N_GND_M1007_b N_Y_c_570_n 0.00793787f $X=-0.045 $Y=0 $X2=3.125 $Y2=1.22
cc_120 N_GND_c_38_p N_Y_c_570_n 0.0142303f $X=2.84 $Y=0.865 $X2=3.125 $Y2=1.22
cc_121 N_GND_M1007_b N_Y_c_573_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.22
cc_122 N_GND_c_24_p N_Y_c_573_n 7.53951e-19 $X=1.98 $Y=0.865 $X2=2.555 $Y2=1.22
cc_123 N_GND_c_38_p N_Y_c_573_n 7.53951e-19 $X=2.84 $Y=0.865 $X2=2.555 $Y2=1.22
cc_124 N_GND_M1007_b N_Y_c_576_n 0.0144211f $X=-0.045 $Y=0 $X2=3.125 $Y2=2.33
cc_125 N_GND_M1007_b N_Y_c_577_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.33
cc_126 N_GND_M1007_b N_Y_c_578_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.335
cc_127 N_GND_c_38_p N_Y_c_578_n 7.53951e-19 $X=2.84 $Y=0.865 $X2=3.27 $Y2=1.335
cc_128 N_GND_c_52_p N_Y_c_578_n 8.22956e-19 $X=3.7 $Y=0.865 $X2=3.27 $Y2=1.335
cc_129 N_GND_M1007_b N_Y_c_581_n 0.0358528f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.215
cc_130 N_GND_M1007_b N_Y_c_582_n 0.018807f $X=-0.045 $Y=0 $X2=3.985 $Y2=2.33
cc_131 N_GND_M1007_b N_Y_c_583_n 0.00584404f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.33
cc_132 N_GND_M1007_b N_Y_c_584_n 0.00409378f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.335
cc_133 N_GND_c_52_p N_Y_c_584_n 7.53951e-19 $X=3.7 $Y=0.865 $X2=4.13 $Y2=1.335
cc_134 N_GND_c_65_p N_Y_c_584_n 0.00134792f $X=4.56 $Y=0.865 $X2=4.13 $Y2=1.335
cc_135 N_GND_M1007_b N_Y_c_587_n 0.06145f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.215
cc_136 N_GND_M1015_s N_Y_c_588_n 0.00418405f $X=3.56 $Y=0.575 $X2=4.13 $Y2=1.22
cc_137 N_GND_M1007_b N_Y_c_588_n 0.00806676f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.22
cc_138 N_GND_c_52_p N_Y_c_588_n 0.0140638f $X=3.7 $Y=0.865 $X2=4.13 $Y2=1.22
cc_139 N_VDD_M1010_b N_B_M1010_g 0.0264002f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_140 N_VDD_c_140_p N_B_M1010_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_141 N_VDD_c_141_p N_B_M1010_g 0.00429146f $X=4.42 $Y=5.36 $X2=0.475 $Y2=3.825
cc_142 N_VDD_M1010_b N_B_c_226_n 0.00375034f $X=-0.045 $Y=2.645 $X2=0.27
+ $Y2=2.415
cc_143 N_VDD_M1010_b B 0.0108395f $X=-0.045 $Y=2.645 $X2=0.27 $Y2=2.7
cc_144 N_VDD_M1010_b N_A_M1005_g 0.0199048f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_145 N_VDD_c_140_p N_A_M1005_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905
+ $Y2=3.825
cc_146 N_VDD_c_146_p N_A_M1005_g 0.00362996f $X=1.12 $Y=3.885 $X2=0.905
+ $Y2=3.825
cc_147 N_VDD_c_141_p N_A_M1005_g 0.00429146f $X=4.42 $Y=5.36 $X2=0.905 $Y2=3.825
cc_148 N_VDD_M1010_b N_A_c_254_n 0.00153494f $X=-0.045 $Y=2.645 $X2=0.95
+ $Y2=2.125
cc_149 N_VDD_M1005_d A 0.0077995f $X=0.98 $Y=2.825 $X2=0.95 $Y2=3.07
cc_150 N_VDD_c_146_p A 0.00247404f $X=1.12 $Y=3.885 $X2=0.95 $Y2=3.07
cc_151 N_VDD_M1010_b N_A_27_565#_c_362_n 0.0174876f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.7
cc_152 N_VDD_c_146_p N_A_27_565#_c_362_n 0.00362996f $X=1.12 $Y=3.885 $X2=1.335
+ $Y2=2.7
cc_153 N_VDD_c_153_p N_A_27_565#_c_362_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335
+ $Y2=2.7
cc_154 N_VDD_c_141_p N_A_27_565#_c_362_n 0.00429146f $X=4.42 $Y=5.36 $X2=1.335
+ $Y2=2.7
cc_155 N_VDD_M1010_b N_A_27_565#_c_297_n 0.00427883f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_156 N_VDD_M1010_b N_A_27_565#_c_367_n 0.0173909f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.7
cc_157 N_VDD_c_146_p N_A_27_565#_c_367_n 3.67508e-19 $X=1.12 $Y=3.885 $X2=1.765
+ $Y2=2.7
cc_158 N_VDD_c_153_p N_A_27_565#_c_367_n 0.00500229f $X=1.895 $Y=5.397 $X2=1.765
+ $Y2=2.7
cc_159 N_VDD_c_159_p N_A_27_565#_c_367_n 0.00382402f $X=1.98 $Y=3.205 $X2=1.765
+ $Y2=2.7
cc_160 N_VDD_c_141_p N_A_27_565#_c_367_n 0.00430409f $X=4.42 $Y=5.36 $X2=1.765
+ $Y2=2.7
cc_161 N_VDD_M1010_b N_A_27_565#_c_305_n 0.00396043f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.625
cc_162 N_VDD_c_159_p N_A_27_565#_c_305_n 0.00379272f $X=1.98 $Y=3.205 $X2=2.12
+ $Y2=2.625
cc_163 N_VDD_M1010_b N_A_27_565#_c_374_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.7
cc_164 N_VDD_c_159_p N_A_27_565#_c_374_n 0.00362996f $X=1.98 $Y=3.205 $X2=2.195
+ $Y2=2.7
cc_165 N_VDD_c_165_p N_A_27_565#_c_374_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.195
+ $Y2=2.7
cc_166 N_VDD_c_141_p N_A_27_565#_c_374_n 0.00429146f $X=4.42 $Y=5.36 $X2=2.195
+ $Y2=2.7
cc_167 N_VDD_M1010_b N_A_27_565#_c_311_n 0.00448664f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.625
cc_168 N_VDD_M1010_b N_A_27_565#_c_379_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.7
cc_169 N_VDD_c_165_p N_A_27_565#_c_379_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.625
+ $Y2=2.7
cc_170 N_VDD_c_170_p N_A_27_565#_c_379_n 0.00362996f $X=2.84 $Y=3.205 $X2=2.625
+ $Y2=2.7
cc_171 N_VDD_c_141_p N_A_27_565#_c_379_n 0.00429146f $X=4.42 $Y=5.36 $X2=2.625
+ $Y2=2.7
cc_172 N_VDD_M1010_b N_A_27_565#_c_318_n 0.00396043f $X=-0.045 $Y=2.645 $X2=2.98
+ $Y2=2.625
cc_173 N_VDD_c_170_p N_A_27_565#_c_318_n 0.00379272f $X=2.84 $Y=3.205 $X2=2.98
+ $Y2=2.625
cc_174 N_VDD_M1010_b N_A_27_565#_c_385_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.055
+ $Y2=2.7
cc_175 N_VDD_c_170_p N_A_27_565#_c_385_n 0.00362996f $X=2.84 $Y=3.205 $X2=3.055
+ $Y2=2.7
cc_176 N_VDD_c_176_p N_A_27_565#_c_385_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.055
+ $Y2=2.7
cc_177 N_VDD_c_141_p N_A_27_565#_c_385_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.055
+ $Y2=2.7
cc_178 N_VDD_M1010_b N_A_27_565#_c_325_n 0.00448664f $X=-0.045 $Y=2.645 $X2=3.41
+ $Y2=2.625
cc_179 N_VDD_M1010_b N_A_27_565#_c_390_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.485
+ $Y2=2.7
cc_180 N_VDD_c_176_p N_A_27_565#_c_390_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.485
+ $Y2=2.7
cc_181 N_VDD_c_181_p N_A_27_565#_c_390_n 0.00362996f $X=3.7 $Y=3.205 $X2=3.485
+ $Y2=2.7
cc_182 N_VDD_c_141_p N_A_27_565#_c_390_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.485
+ $Y2=2.7
cc_183 N_VDD_M1010_b N_A_27_565#_c_332_n 0.00396043f $X=-0.045 $Y=2.645 $X2=3.84
+ $Y2=2.625
cc_184 N_VDD_c_181_p N_A_27_565#_c_332_n 0.00379272f $X=3.7 $Y=3.205 $X2=3.84
+ $Y2=2.625
cc_185 N_VDD_M1010_b N_A_27_565#_c_396_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.915
+ $Y2=2.7
cc_186 N_VDD_c_181_p N_A_27_565#_c_396_n 0.00362996f $X=3.7 $Y=3.205 $X2=3.915
+ $Y2=2.7
cc_187 N_VDD_c_187_p N_A_27_565#_c_396_n 0.00496961f $X=4.475 $Y=5.397 $X2=3.915
+ $Y2=2.7
cc_188 N_VDD_c_141_p N_A_27_565#_c_396_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.915
+ $Y2=2.7
cc_189 N_VDD_M1010_b N_A_27_565#_c_338_n 0.00840215f $X=-0.045 $Y=2.645 $X2=4.27
+ $Y2=2.625
cc_190 N_VDD_M1010_b N_A_27_565#_c_401_n 0.0212947f $X=-0.045 $Y=2.645 $X2=4.345
+ $Y2=2.7
cc_191 N_VDD_c_187_p N_A_27_565#_c_401_n 0.00496961f $X=4.475 $Y=5.397 $X2=4.345
+ $Y2=2.7
cc_192 N_VDD_c_192_p N_A_27_565#_c_401_n 0.00751602f $X=4.56 $Y=3.205 $X2=4.345
+ $Y2=2.7
cc_193 N_VDD_c_141_p N_A_27_565#_c_401_n 0.00429146f $X=4.42 $Y=5.36 $X2=4.345
+ $Y2=2.7
cc_194 N_VDD_M1010_b N_A_27_565#_c_343_n 0.0021704f $X=-0.045 $Y=2.645 $X2=1.352
+ $Y2=2.625
cc_195 N_VDD_M1010_b N_A_27_565#_c_344_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=1.765 $Y2=2.625
cc_196 N_VDD_M1010_b N_A_27_565#_c_346_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.195 $Y2=2.625
cc_197 N_VDD_M1010_b N_A_27_565#_c_348_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.625 $Y2=2.625
cc_198 N_VDD_M1010_b N_A_27_565#_c_350_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.055 $Y2=2.625
cc_199 N_VDD_M1010_b N_A_27_565#_c_352_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.485 $Y2=2.625
cc_200 N_VDD_M1010_b N_A_27_565#_c_354_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.915 $Y2=2.625
cc_201 N_VDD_M1010_b N_A_27_565#_c_412_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.545
cc_202 N_VDD_c_140_p N_A_27_565#_c_412_n 0.00452684f $X=1.035 $Y=5.397 $X2=0.26
+ $Y2=3.545
cc_203 N_VDD_c_141_p N_A_27_565#_c_412_n 0.00435496f $X=4.42 $Y=5.36 $X2=0.26
+ $Y2=3.545
cc_204 N_VDD_M1010_b N_A_27_565#_c_355_n 0.00106577f $X=-0.045 $Y=2.645 $X2=0.61
+ $Y2=3.285
cc_205 N_VDD_M1010_b N_Y_c_542_n 0.00410619f $X=-0.045 $Y=2.645 $X2=1.55
+ $Y2=2.33
cc_206 N_VDD_c_153_p N_Y_c_542_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.33
cc_207 N_VDD_c_141_p N_Y_c_542_n 0.00434939f $X=4.42 $Y=5.36 $X2=1.55 $Y2=2.33
cc_208 N_VDD_M1010_b N_Y_c_548_n 0.0042387f $X=-0.045 $Y=2.645 $X2=2.41 $Y2=2.33
cc_209 N_VDD_c_165_p N_Y_c_548_n 0.0045126f $X=2.755 $Y=5.397 $X2=2.41 $Y2=2.33
cc_210 N_VDD_c_141_p N_Y_c_548_n 0.00434939f $X=4.42 $Y=5.36 $X2=2.41 $Y2=2.33
cc_211 N_VDD_M1010_b N_Y_c_554_n 0.0042387f $X=-0.045 $Y=2.645 $X2=3.27 $Y2=2.33
cc_212 N_VDD_c_176_p N_Y_c_554_n 0.00464147f $X=3.615 $Y=5.397 $X2=3.27 $Y2=2.33
cc_213 N_VDD_c_141_p N_Y_c_554_n 0.00434939f $X=4.42 $Y=5.36 $X2=3.27 $Y2=2.33
cc_214 N_VDD_M1010_b N_Y_c_559_n 0.0042387f $X=-0.045 $Y=2.645 $X2=4.13 $Y2=2.33
cc_215 N_VDD_c_187_p N_Y_c_559_n 0.00475585f $X=4.475 $Y=5.397 $X2=4.13 $Y2=2.33
cc_216 N_VDD_c_141_p N_Y_c_559_n 0.00434939f $X=4.42 $Y=5.36 $X2=4.13 $Y2=2.33
cc_217 N_VDD_c_159_p N_Y_c_568_n 0.00634153f $X=1.98 $Y=3.205 $X2=2.265 $Y2=2.33
cc_218 N_VDD_c_170_p N_Y_c_576_n 0.00634153f $X=2.84 $Y=3.205 $X2=3.125 $Y2=2.33
cc_219 N_VDD_c_181_p N_Y_c_582_n 0.00634153f $X=3.7 $Y=3.205 $X2=3.985 $Y2=2.33
cc_220 N_B_M1007_g N_A_M1002_g 0.0430073f $X=0.475 $Y=0.895 $X2=0.905 $Y2=0.895
cc_221 N_B_c_225_n N_A_M1005_g 0.112923f $X=0.475 $Y=2.415 $X2=0.905 $Y2=3.825
cc_222 N_B_M1007_g N_A_c_253_n 0.0148656f $X=0.475 $Y=0.895 $X2=0.95 $Y2=2.125
cc_223 N_B_M1007_g N_A_c_254_n 0.00121111f $X=0.475 $Y=0.895 $X2=0.95 $Y2=2.125
cc_224 N_B_M1010_g N_A_27_565#_c_416_n 0.0142177f $X=0.475 $Y=3.825 $X2=0.525
+ $Y2=3.37
cc_225 B N_A_27_565#_c_416_n 0.00520961f $X=0.27 $Y=2.7 $X2=0.525 $Y2=3.37
cc_226 N_B_c_226_n N_A_27_565#_c_418_n 0.00369517f $X=0.27 $Y=2.415 $X2=0.345
+ $Y2=3.37
cc_227 B N_A_27_565#_c_418_n 0.00431991f $X=0.27 $Y=2.7 $X2=0.345 $Y2=3.37
cc_228 N_B_M1007_g N_A_27_565#_c_355_n 0.0231435f $X=0.475 $Y=0.895 $X2=0.61
+ $Y2=3.285
cc_229 N_B_M1010_g N_A_27_565#_c_355_n 0.026563f $X=0.475 $Y=3.825 $X2=0.61
+ $Y2=3.285
cc_230 N_B_c_225_n N_A_27_565#_c_355_n 0.00764878f $X=0.475 $Y=2.415 $X2=0.61
+ $Y2=3.285
cc_231 N_B_c_226_n N_A_27_565#_c_355_n 0.0350086f $X=0.27 $Y=2.415 $X2=0.61
+ $Y2=3.285
cc_232 B N_A_27_565#_c_355_n 0.00758489f $X=0.27 $Y=2.7 $X2=0.61 $Y2=3.285
cc_233 N_B_M1007_g N_A_27_565#_c_356_n 0.00996235f $X=0.475 $Y=0.895 $X2=0.69
+ $Y2=0.865
cc_234 N_B_M1007_g N_A_27_565#_c_361_n 0.0113001f $X=0.475 $Y=0.895 $X2=0.65
+ $Y2=1.675
cc_235 N_A_M1002_g N_A_27_565#_M1004_g 0.0337969f $X=0.905 $Y=0.895 $X2=1.335
+ $Y2=0.895
cc_236 A N_A_27_565#_c_362_n 0.00374181f $X=0.95 $Y=3.07 $X2=1.335 $Y2=2.7
cc_237 N_A_M1005_g N_A_27_565#_c_296_n 0.00914307f $X=0.905 $Y=3.825 $X2=1.37
+ $Y2=2.55
cc_238 N_A_c_253_n N_A_27_565#_c_296_n 0.0204279f $X=0.95 $Y=2.125 $X2=1.37
+ $Y2=2.55
cc_239 N_A_c_254_n N_A_27_565#_c_296_n 0.00375034f $X=0.95 $Y=2.125 $X2=1.37
+ $Y2=2.55
cc_240 N_A_M1002_g N_A_27_565#_c_304_n 0.0119161f $X=0.905 $Y=0.895 $X2=1.84
+ $Y2=1.585
cc_241 N_A_M1005_g N_A_27_565#_c_343_n 0.0554147f $X=0.905 $Y=3.825 $X2=1.352
+ $Y2=2.625
cc_242 N_A_c_254_n N_A_27_565#_c_343_n 0.00358357f $X=0.95 $Y=2.125 $X2=1.352
+ $Y2=2.625
cc_243 N_A_M1005_g N_A_27_565#_c_416_n 0.00457566f $X=0.905 $Y=3.825 $X2=0.525
+ $Y2=3.37
cc_244 N_A_M1002_g N_A_27_565#_c_355_n 0.00429604f $X=0.905 $Y=0.895 $X2=0.61
+ $Y2=3.285
cc_245 N_A_M1005_g N_A_27_565#_c_355_n 0.00776428f $X=0.905 $Y=3.825 $X2=0.61
+ $Y2=3.285
cc_246 N_A_c_253_n N_A_27_565#_c_355_n 0.0021255f $X=0.95 $Y=2.125 $X2=0.61
+ $Y2=3.285
cc_247 N_A_c_254_n N_A_27_565#_c_355_n 0.0822139f $X=0.95 $Y=2.125 $X2=0.61
+ $Y2=3.285
cc_248 A N_A_27_565#_c_355_n 0.00866797f $X=0.95 $Y=3.07 $X2=0.61 $Y2=3.285
cc_249 N_A_M1002_g N_A_27_565#_c_356_n 0.00996235f $X=0.905 $Y=0.895 $X2=0.69
+ $Y2=0.865
cc_250 N_A_M1002_g N_A_27_565#_c_359_n 0.0163305f $X=0.905 $Y=0.895 $X2=1.43
+ $Y2=1.675
cc_251 N_A_c_253_n N_A_27_565#_c_359_n 0.00276813f $X=0.95 $Y=2.125 $X2=1.43
+ $Y2=1.675
cc_252 N_A_c_254_n N_A_27_565#_c_359_n 0.0114342f $X=0.95 $Y=2.125 $X2=1.43
+ $Y2=1.675
cc_253 A A_110_565# 0.0123256f $X=0.95 $Y=3.07 $X2=0.55 $Y2=2.825
cc_254 N_A_c_254_n N_Y_c_542_n 0.0206732f $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.33
cc_255 A N_Y_c_542_n 0.00659455f $X=0.95 $Y=3.07 $X2=1.55 $Y2=2.33
cc_256 N_A_M1002_g N_Y_c_560_n 8.23842e-19 $X=0.905 $Y=0.895 $X2=1.55 $Y2=1.335
cc_257 N_A_c_253_n N_Y_c_563_n 3.73261e-19 $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.215
cc_258 N_A_c_254_n N_Y_c_563_n 0.0059581f $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.215
cc_259 N_A_M1002_g Y 6.73508e-19 $X=0.905 $Y=0.895 $X2=1.555 $Y2=1.96
cc_260 N_A_c_254_n Y 0.00825539f $X=0.95 $Y=2.125 $X2=1.555 $Y2=1.96
cc_261 N_A_27_565#_c_416_n A_110_565# 0.00613297f $X=0.525 $Y=3.37 $X2=0.55
+ $Y2=2.825
cc_262 N_A_27_565#_c_355_n A_110_565# 0.00377193f $X=0.61 $Y=3.285 $X2=0.55
+ $Y2=2.825
cc_263 N_A_27_565#_M1004_g N_Y_c_538_n 0.00339663f $X=1.335 $Y=0.895 $X2=1.55
+ $Y2=0.865
cc_264 N_A_27_565#_M1008_g N_Y_c_538_n 0.00339663f $X=1.765 $Y=0.895 $X2=1.55
+ $Y2=0.865
cc_265 N_A_27_565#_c_304_n N_Y_c_538_n 0.00171364f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=0.865
cc_266 N_A_27_565#_c_359_n N_Y_c_538_n 0.00520269f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.865
cc_267 N_A_27_565#_c_362_n N_Y_c_542_n 0.00234922f $X=1.335 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_268 N_A_27_565#_c_296_n N_Y_c_542_n 0.00744772f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_269 N_A_27_565#_c_297_n N_Y_c_542_n 0.0156814f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_270 N_A_27_565#_c_367_n N_Y_c_542_n 0.00401146f $X=1.765 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_271 N_A_27_565#_c_304_n N_Y_c_542_n 0.00182797f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.33
cc_272 N_A_27_565#_c_359_n N_Y_c_542_n 0.00273485f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_273 N_A_27_565#_M1009_g N_Y_c_543_n 0.00339663f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=0.865
cc_274 N_A_27_565#_c_310_n N_Y_c_543_n 0.00280419f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=0.865
cc_275 N_A_27_565#_M1013_g N_Y_c_543_n 0.00339663f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=0.865
cc_276 N_A_27_565#_c_374_n N_Y_c_548_n 0.00401146f $X=2.195 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_277 N_A_27_565#_c_310_n N_Y_c_548_n 0.00250559f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.33
cc_278 N_A_27_565#_c_311_n N_Y_c_548_n 0.021445f $X=2.55 $Y=2.625 $X2=2.41
+ $Y2=2.33
cc_279 N_A_27_565#_c_379_n N_Y_c_548_n 0.00401146f $X=2.625 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_280 N_A_27_565#_c_323_n N_Y_c_548_n 0.00361281f $X=3.055 $Y=2.55 $X2=2.41
+ $Y2=2.33
cc_281 N_A_27_565#_M1014_g N_Y_c_549_n 0.00339663f $X=3.055 $Y=0.895 $X2=3.27
+ $Y2=0.865
cc_282 N_A_27_565#_c_324_n N_Y_c_549_n 0.00280419f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=0.865
cc_283 N_A_27_565#_M1015_g N_Y_c_549_n 0.00339663f $X=3.485 $Y=0.895 $X2=3.27
+ $Y2=0.865
cc_284 N_A_27_565#_c_323_n N_Y_c_554_n 0.00721971f $X=3.055 $Y=2.55 $X2=3.27
+ $Y2=2.33
cc_285 N_A_27_565#_c_385_n N_Y_c_554_n 0.00401146f $X=3.055 $Y=2.7 $X2=3.27
+ $Y2=2.33
cc_286 N_A_27_565#_c_324_n N_Y_c_554_n 0.00250559f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=2.33
cc_287 N_A_27_565#_c_325_n N_Y_c_554_n 0.021445f $X=3.41 $Y=2.625 $X2=3.27
+ $Y2=2.33
cc_288 N_A_27_565#_c_390_n N_Y_c_554_n 0.00401146f $X=3.485 $Y=2.7 $X2=3.27
+ $Y2=2.33
cc_289 N_A_27_565#_M1016_g N_Y_c_555_n 0.00339663f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=0.865
cc_290 N_A_27_565#_c_337_n N_Y_c_555_n 0.00280419f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=0.865
cc_291 N_A_27_565#_M1017_g N_Y_c_555_n 0.00339663f $X=4.345 $Y=0.895 $X2=4.13
+ $Y2=0.865
cc_292 N_A_27_565#_c_396_n N_Y_c_559_n 0.00401146f $X=3.915 $Y=2.7 $X2=4.13
+ $Y2=2.33
cc_293 N_A_27_565#_c_337_n N_Y_c_559_n 0.00250559f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=2.33
cc_294 N_A_27_565#_c_338_n N_Y_c_559_n 0.0206674f $X=4.27 $Y=2.625 $X2=4.13
+ $Y2=2.33
cc_295 N_A_27_565#_c_401_n N_Y_c_559_n 0.00401146f $X=4.345 $Y=2.7 $X2=4.13
+ $Y2=2.33
cc_296 N_A_27_565#_M1004_g N_Y_c_560_n 0.00542903f $X=1.335 $Y=0.895 $X2=1.55
+ $Y2=1.335
cc_297 N_A_27_565#_M1008_g N_Y_c_560_n 0.00259902f $X=1.765 $Y=0.895 $X2=1.55
+ $Y2=1.335
cc_298 N_A_27_565#_c_359_n N_Y_c_560_n 0.00238892f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=1.335
cc_299 N_A_27_565#_c_296_n N_Y_c_563_n 0.00821104f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.215
cc_300 N_A_27_565#_c_297_n N_Y_c_563_n 0.00186325f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.215
cc_301 N_A_27_565#_c_304_n N_Y_c_563_n 0.00194187f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.215
cc_302 N_A_27_565#_c_359_n N_Y_c_563_n 0.00181779f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.215
cc_303 N_A_27_565#_M1004_g Y 0.00251111f $X=1.335 $Y=0.895 $X2=1.555 $Y2=1.96
cc_304 N_A_27_565#_c_296_n Y 0.00892438f $X=1.37 $Y=2.55 $X2=1.555 $Y2=1.96
cc_305 N_A_27_565#_M1008_g Y 0.00251111f $X=1.765 $Y=0.895 $X2=1.555 $Y2=1.96
cc_306 N_A_27_565#_c_304_n Y 0.0131034f $X=1.84 $Y=1.585 $X2=1.555 $Y2=1.96
cc_307 N_A_27_565#_c_359_n Y 0.0147088f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_308 N_A_27_565#_M1008_g N_Y_c_565_n 0.0130095f $X=1.765 $Y=0.895 $X2=2.265
+ $Y2=1.22
cc_309 N_A_27_565#_c_302_n N_Y_c_565_n 0.00213861f $X=2.12 $Y=1.585 $X2=2.265
+ $Y2=1.22
cc_310 N_A_27_565#_M1009_g N_Y_c_565_n 0.0130095f $X=2.195 $Y=0.895 $X2=2.265
+ $Y2=1.22
cc_311 N_A_27_565#_c_304_n N_Y_c_568_n 0.0121767f $X=1.84 $Y=1.585 $X2=2.265
+ $Y2=2.33
cc_312 N_A_27_565#_c_344_n N_Y_c_568_n 0.0158479f $X=1.765 $Y=2.625 $X2=2.265
+ $Y2=2.33
cc_313 N_A_27_565#_M1009_g N_Y_c_569_n 0.00251111f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=2.215
cc_314 N_A_27_565#_c_310_n N_Y_c_569_n 0.0177725f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_315 N_A_27_565#_M1013_g N_Y_c_569_n 0.00251111f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=2.215
cc_316 N_A_27_565#_c_323_n N_Y_c_569_n 0.00843025f $X=3.055 $Y=2.55 $X2=2.41
+ $Y2=2.215
cc_317 N_A_27_565#_M1013_g N_Y_c_570_n 0.0130095f $X=2.625 $Y=0.895 $X2=3.125
+ $Y2=1.22
cc_318 N_A_27_565#_c_316_n N_Y_c_570_n 0.00213861f $X=2.98 $Y=1.585 $X2=3.125
+ $Y2=1.22
cc_319 N_A_27_565#_M1014_g N_Y_c_570_n 0.0136594f $X=3.055 $Y=0.895 $X2=3.125
+ $Y2=1.22
cc_320 N_A_27_565#_M1009_g N_Y_c_573_n 0.00259902f $X=2.195 $Y=0.895 $X2=2.555
+ $Y2=1.22
cc_321 N_A_27_565#_M1013_g N_Y_c_573_n 0.00259902f $X=2.625 $Y=0.895 $X2=2.555
+ $Y2=1.22
cc_322 N_A_27_565#_c_323_n N_Y_c_576_n 0.0155956f $X=3.055 $Y=2.55 $X2=3.125
+ $Y2=2.33
cc_323 N_A_27_565#_c_347_n N_Y_c_576_n 0.00894336f $X=2.625 $Y=1.585 $X2=3.125
+ $Y2=2.33
cc_324 N_A_27_565#_c_348_n N_Y_c_576_n 0.00903839f $X=2.625 $Y=2.625 $X2=3.125
+ $Y2=2.33
cc_325 N_A_27_565#_c_310_n N_Y_c_577_n 0.00140336f $X=2.55 $Y=1.585 $X2=2.555
+ $Y2=2.33
cc_326 N_A_27_565#_c_323_n N_Y_c_577_n 0.0012308f $X=3.055 $Y=2.55 $X2=2.555
+ $Y2=2.33
cc_327 N_A_27_565#_c_345_n N_Y_c_577_n 0.00140336f $X=2.195 $Y=1.585 $X2=2.555
+ $Y2=2.33
cc_328 N_A_27_565#_c_346_n N_Y_c_577_n 0.00372651f $X=2.195 $Y=2.625 $X2=2.555
+ $Y2=2.33
cc_329 N_A_27_565#_M1014_g N_Y_c_578_n 0.00262362f $X=3.055 $Y=0.895 $X2=3.27
+ $Y2=1.335
cc_330 N_A_27_565#_M1015_g N_Y_c_578_n 0.00394441f $X=3.485 $Y=0.895 $X2=3.27
+ $Y2=1.335
cc_331 N_A_27_565#_M1016_g N_Y_c_578_n 2.43068e-19 $X=3.915 $Y=0.895 $X2=3.27
+ $Y2=1.335
cc_332 N_A_27_565#_M1014_g N_Y_c_581_n 0.00251111f $X=3.055 $Y=0.895 $X2=3.27
+ $Y2=2.215
cc_333 N_A_27_565#_c_323_n N_Y_c_581_n 0.0108556f $X=3.055 $Y=2.55 $X2=3.27
+ $Y2=2.215
cc_334 N_A_27_565#_c_324_n N_Y_c_581_n 0.0177725f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=2.215
cc_335 N_A_27_565#_M1015_g N_Y_c_581_n 0.00251111f $X=3.485 $Y=0.895 $X2=3.27
+ $Y2=2.215
cc_336 N_A_27_565#_c_351_n N_Y_c_582_n 0.0121767f $X=3.485 $Y=1.585 $X2=3.985
+ $Y2=2.33
cc_337 N_A_27_565#_c_352_n N_Y_c_582_n 0.0158479f $X=3.485 $Y=2.625 $X2=3.985
+ $Y2=2.33
cc_338 N_A_27_565#_c_323_n N_Y_c_583_n 0.00618817f $X=3.055 $Y=2.55 $X2=3.415
+ $Y2=2.33
cc_339 N_A_27_565#_c_324_n N_Y_c_583_n 0.00268861f $X=3.41 $Y=1.585 $X2=3.415
+ $Y2=2.33
cc_340 N_A_27_565#_c_325_n N_Y_c_583_n 0.00357274f $X=3.41 $Y=2.625 $X2=3.415
+ $Y2=2.33
cc_341 N_A_27_565#_M1016_g N_Y_c_584_n 0.00259902f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=1.335
cc_342 N_A_27_565#_M1017_g N_Y_c_584_n 0.00954936f $X=4.345 $Y=0.895 $X2=4.13
+ $Y2=1.335
cc_343 N_A_27_565#_M1016_g N_Y_c_587_n 0.00251111f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=2.215
cc_344 N_A_27_565#_c_337_n N_Y_c_587_n 0.0184054f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=2.215
cc_345 N_A_27_565#_M1017_g N_Y_c_587_n 0.00251111f $X=4.345 $Y=0.895 $X2=4.13
+ $Y2=2.215
cc_346 N_A_27_565#_c_353_n N_Y_c_587_n 0.00140336f $X=3.915 $Y=1.585 $X2=4.13
+ $Y2=2.215
cc_347 N_A_27_565#_c_354_n N_Y_c_587_n 0.00372651f $X=3.915 $Y=2.625 $X2=4.13
+ $Y2=2.215
cc_348 N_A_27_565#_M1015_g N_Y_c_588_n 8.84842e-19 $X=3.485 $Y=0.895 $X2=4.13
+ $Y2=1.22
cc_349 N_A_27_565#_c_330_n N_Y_c_588_n 0.00213861f $X=3.84 $Y=1.585 $X2=4.13
+ $Y2=1.22
cc_350 N_A_27_565#_M1016_g N_Y_c_588_n 0.0130426f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=1.22
