* File: sky130_osu_sc_12T_ms__dff_1.spice
* Created: Fri Nov 12 15:22:21 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ms__dff_1.pex.spice"
.subckt sky130_osu_sc_12T_ms__dff_1  GND VDD D CK ON Q
* 
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A_75_248#_M1004_g N_A_32_115#_M1004_s N_GND_M1004_b
+ NSHORT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75004.1 A=0.078 P=1.34 MULT=1
MM1003 A_201_115# N_D_M1003_g N_GND_M1004_d N_GND_M1004_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75003.7 A=0.078 P=1.34 MULT=1
MM1021 N_A_75_248#_M1021_d N_A_243_89#_M1021_g A_201_115# N_GND_M1004_b NSHORT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75001 SB=75003.3 A=0.078 P=1.34 MULT=1
MM1016 A_393_115# N_CK_M1016_g N_A_75_248#_M1021_d N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.6 SB=75002.7 A=0.078 P=1.34 MULT=1
MM1010 N_GND_M1010_d N_A_32_115#_M1010_g A_393_115# N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1011 A_551_115# N_A_32_115#_M1011_g N_GND_M1010_d N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1009 N_A_623_115#_M1009_d N_CK_M1009_g A_551_115# N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75002.7 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1001 A_743_115# N_A_243_89#_M1001_g N_A_623_115#_M1009_d N_GND_M1004_b NSHORT
+ L=0.15 W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1
+ R=3.46667 SA=75003.3 SB=75001 A=0.078 P=1.34 MULT=1
MM1023 N_GND_M1023_d N_A_785_89#_M1023_g A_743_115# N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75003.7 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1024 N_A_243_89#_M1024_d N_CK_M1024_g N_GND_M1023_d N_GND_M1004_b NSHORT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75004.1 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1006 N_A_785_89#_M1006_d N_A_623_115#_M1006_g N_GND_M1006_s N_GND_M1004_b
+ NSHORT L=0.15 W=0.52 AD=0.1378 AS=0.1378 PD=1.57 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_A_785_89#_M1007_g N_ON_M1007_s N_GND_M1004_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1025 N_Q_M1025_d N_ON_M1025_g N_GND_M1007_d N_GND_M1004_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1019 N_VDD_M1019_d N_A_75_248#_M1019_g N_A_32_115#_M1019_s N_VDD_M1019_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1018 A_201_521# N_D_M1018_g N_VDD_M1019_d N_VDD_M1019_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1012 N_A_75_248#_M1012_d N_CK_M1012_g A_201_521# N_VDD_M1019_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1008 A_393_521# N_A_243_89#_M1008_g N_A_75_248#_M1012_d N_VDD_M1019_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.6 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1002 N_VDD_M1002_d N_A_32_115#_M1002_g A_393_521# N_VDD_M1019_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1005 A_551_521# N_A_32_115#_M1005_g N_VDD_M1002_d N_VDD_M1019_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1000 N_A_623_115#_M1000_d N_A_243_89#_M1000_g A_551_521# N_VDD_M1019_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.7 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1017 A_743_521# N_CK_M1017_g N_A_623_115#_M1000_d N_VDD_M1019_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75003.3 SB=75001 A=0.189 P=2.82 MULT=1
MM1013 N_VDD_M1013_d N_A_785_89#_M1013_g A_743_521# N_VDD_M1019_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_243_89#_M1014_d N_CK_M1014_g N_VDD_M1013_d N_VDD_M1019_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1020 N_A_785_89#_M1020_d N_A_623_115#_M1020_g N_VDD_M1020_s N_VDD_M1019_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1022 N_VDD_M1022_d N_A_785_89#_M1022_g N_ON_M1022_s N_VDD_M1019_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_Q_M1015_d N_ON_M1015_g N_VDD_M1022_d N_VDD_M1019_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref N_GND_M1004_b N_VDD_M1019_b NWDIODE A=15.0895 P=18.77
pX27_noxref noxref_20 D D PROBETYPE=1
pX28_noxref noxref_21 CK CK PROBETYPE=1
pX29_noxref noxref_22 ON ON PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
c_1311 A_551_521# 0 1.57671e-19 $X=2.755 $Y=2.605
*
.include "sky130_osu_sc_12T_ms__dff_1.pxi.spice"
*
.ends
*
*
