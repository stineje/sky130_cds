* File: sky130_osu_sc_12T_ls__tbufi_l.spice
* Created: Fri Nov 12 15:40:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__tbufi_l.pex.spice"
.subckt sky130_osu_sc_12T_ls__tbufi_l  GND VDD OE A Y
* 
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_OE_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NSHORT
+ L=0.15 W=0.36 AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75001 A=0.054 P=1.02 MULT=1
MM1000 A_196_115# N_OE_M1000_g N_GND_M1002_d N_GND_M1002_b NSHORT L=0.15 W=0.36
+ AD=0.0378 AS=0.0504 PD=0.57 PS=0.64 NRD=16.656 NRS=0 M=1 R=2.4 SA=75000.6
+ SB=75000.6 A=0.054 P=1.02 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_196_115# N_GND_M1002_b NSHORT L=0.15 W=0.36
+ AD=0.0954 AS=0.0378 PD=1.25 PS=0.57 NRD=0 NRS=16.656 M=1 R=2.4 SA=75001
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1001 N_VDD_M1001_d N_OE_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1003 A_196_605# N_A_27_115#_M1003_g N_VDD_M1001_d N_VDD_M1001_b PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g A_196_605# N_VDD_M1001_b PHIGHVT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=3.2448 P=7.22
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__tbufi_l.pxi.spice"
*
.ends
*
*
