* File: sky130_osu_sc_12T_ms__dlat_l.pex.spice
* Created: Fri Nov 12 15:23:38 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%GND 1 2 3 4 59 63 65 75 77 84 86 93 112
+ 114
c121 75 0 1.5259e-19 $X=2.035 $Y=0.74
r122 112 114 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r123 91 93 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.365 $Y=0.305
+ $X2=4.365 $Y2=0.74
r124 82 84 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.985 $Y=0.305
+ $X2=2.985 $Y2=0.74
r125 78 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.152
+ $X2=2.035 $Y2=0.152
r126 73 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.035 $Y=0.305
+ $X2=2.035 $Y2=0.152
r127 73 75 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.035 $Y=0.305
+ $X2=2.035 $Y2=0.74
r128 65 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.152
+ $X2=2.035 $Y2=0.152
r129 61 63 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.285 $Y=0.305
+ $X2=0.285 $Y2=0.74
r130 59 114 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r131 59 112 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r132 59 91 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.365 $Y2=0.305
r133 59 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.28 $Y2=0.152
r134 59 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.985 $Y=0.152
+ $X2=2.985 $Y2=0.305
r135 59 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.152
+ $X2=2.9 $Y2=0.152
r136 59 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.152
+ $X2=3.07 $Y2=0.152
r137 59 61 4.36583 $w=1.7e-07 $l=1.96746e-07 $layer=LI1_cond $X=0.185 $Y=0.152
+ $X2=0.285 $Y2=0.305
r138 59 66 3.19241 $w=3.05e-07 $l=1.85e-07 $layer=LI1_cond $X=0.185 $Y=0.152
+ $X2=0.37 $Y2=0.152
r139 59 86 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.28 $Y2=0.152
r140 59 87 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.07 $Y2=0.152
r141 59 77 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.9 $Y2=0.152
r142 59 78 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.12 $Y2=0.152
r143 59 65 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.95 $Y2=0.152
r144 59 66 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.37 $Y2=0.152
r145 4 93 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.575 $X2=4.365 $Y2=0.74
r146 3 84 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.575 $X2=2.985 $Y2=0.74
r147 2 75 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.575 $X2=2.035 $Y2=0.74
r148 1 63 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%VDD 1 2 3 4 45 49 51 59 61 67 69 75 86
+ 89 93
r63 89 93 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=4.42 $Y2=4.287
r64 86 93 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=4.25
+ $X2=4.42 $Y2=4.25
r65 80 89 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r66 73 86 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.365 $Y=4.135
+ $X2=4.365 $Y2=4.287
r67 73 75 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.365 $Y=4.135
+ $X2=4.365 $Y2=3.615
r68 70 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=4.287
+ $X2=2.985 $Y2=4.287
r69 70 72 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=3.07 $Y=4.287
+ $X2=3.74 $Y2=4.287
r70 69 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=4.287
+ $X2=4.365 $Y2=4.287
r71 69 72 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=4.28 $Y=4.287
+ $X2=3.74 $Y2=4.287
r72 65 84 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.985 $Y=4.135
+ $X2=2.985 $Y2=4.287
r73 65 67 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.985 $Y=4.135
+ $X2=2.985 $Y2=3.275
r74 62 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=4.287
+ $X2=2.035 $Y2=4.287
r75 62 64 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=2.12 $Y=4.287
+ $X2=2.38 $Y2=4.287
r76 61 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=4.287
+ $X2=2.985 $Y2=4.287
r77 61 64 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=2.9 $Y=4.287
+ $X2=2.38 $Y2=4.287
r78 57 82 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.035 $Y=4.135
+ $X2=2.035 $Y2=4.287
r79 57 59 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.035 $Y=4.135
+ $X2=2.035 $Y2=3.275
r80 54 56 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r81 52 80 3.19971 $w=3.05e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=4.287
+ $X2=0.185 $Y2=4.287
r82 52 54 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=0.37 $Y=4.287
+ $X2=1.02 $Y2=4.287
r83 51 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=4.287
+ $X2=2.035 $Y2=4.287
r84 51 56 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.95 $Y=4.287
+ $X2=1.7 $Y2=4.287
r85 47 80 4.35853 $w=1.7e-07 $l=1.95714e-07 $layer=LI1_cond $X=0.285 $Y=4.135
+ $X2=0.185 $Y2=4.287
r86 47 49 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.285 $Y=4.135
+ $X2=0.285 $Y2=3.275
r87 45 86 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=4.135 $X2=4.42 $Y2=4.22
r88 45 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r89 45 84 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r90 45 64 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r91 45 56 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r92 45 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r93 45 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r94 4 75 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=4.225
+ $Y=3.025 $X2=4.365 $Y2=3.615
r95 3 67 300 $w=1.7e-07 $l=7.29829e-07 $layer=licon1_PDIFF $count=2 $X=2.86
+ $Y=2.605 $X2=2.985 $Y2=3.275
r96 2 59 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=1.895
+ $Y=2.605 $X2=2.035 $Y2=3.275
r97 1 49 300 $w=1.7e-07 $l=7.29829e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.605 $X2=0.285 $Y2=3.275
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%D 1 3 11 15 17 19 22 25 31 35 38 39 40
+ 43 47 50 55 62 65 66 72 77 78 80
c127 62 0 1.24842e-20 $X=1.26 $Y=0.74
c128 38 0 1.57671e-19 $X=0.58 $Y=2.62
c129 22 0 3.47982e-21 $X=3.2 $Y=3.235
c130 15 0 1.65121e-19 $X=0.5 $Y=3.235
r131 76 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.26 $Y=1.34
+ $X2=1.405 $Y2=1.34
r132 76 77 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.26 $Y=1.34
+ $X2=1.115 $Y2=1.34
r133 66 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.85 $Y=1.37
+ $X2=2.995 $Y2=1.37
r134 66 78 1.39137 $w=1.7e-07 $l=1.445e-06 $layer=MET1_cond $X=2.85 $Y=1.37
+ $X2=1.405 $Y2=1.37
r135 65 69 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.725 $Y=1.37
+ $X2=0.58 $Y2=1.37
r136 65 77 0.375524 $w=1.7e-07 $l=3.9e-07 $layer=MET1_cond $X=0.725 $Y=1.37
+ $X2=1.115 $Y2=1.37
r137 60 62 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.16 $Y=0.74 $X2=1.26
+ $Y2=0.74
r138 55 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.44 $Y=1.74
+ $X2=0.44 $Y2=1.74
r139 55 58 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.51 $Y=1.74
+ $X2=0.51 $Y2=1.905
r140 55 56 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.51 $Y=1.74
+ $X2=0.51 $Y2=1.575
r141 50 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.995 $Y=1.37
+ $X2=2.995 $Y2=1.37
r142 47 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.26 $Y=1.34
+ $X2=1.26 $Y2=1.34
r143 45 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=0.905
+ $X2=1.26 $Y2=0.74
r144 45 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.26 $Y=0.905
+ $X2=1.26 $Y2=1.34
r145 41 43 16.4393 $w=3.38e-07 $l=4.85e-07 $layer=LI1_cond $X=1.16 $Y=2.79
+ $X2=1.16 $Y2=3.275
r146 39 41 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.99 $Y=2.705
+ $X2=1.16 $Y2=2.79
r147 39 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.99 $Y=2.705
+ $X2=0.665 $Y2=2.705
r148 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.58 $Y=2.62
+ $X2=0.665 $Y2=2.705
r149 38 58 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.58 $Y=2.62
+ $X2=0.58 $Y2=1.905
r150 35 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.58 $Y=1.37
+ $X2=0.58 $Y2=1.37
r151 35 56 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.58 $Y=1.37
+ $X2=0.58 $Y2=1.575
r152 29 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=1.37 $X2=2.995 $Y2=1.37
r153 29 31 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.995 $Y=1.37
+ $X2=3.2 $Y2=1.37
r154 25 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.44
+ $Y=1.74 $X2=0.44 $Y2=1.74
r155 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.44 $Y=1.74
+ $X2=0.44 $Y2=1.905
r156 25 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.44 $Y=1.74
+ $X2=0.44 $Y2=1.575
r157 20 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.535
+ $X2=3.2 $Y2=1.37
r158 20 22 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=3.2 $Y=1.535
+ $X2=3.2 $Y2=3.235
r159 17 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.205
+ $X2=3.2 $Y2=1.37
r160 17 19 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.2 $Y=1.205
+ $X2=3.2 $Y2=0.835
r161 15 27 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.5 $Y=3.235
+ $X2=0.5 $Y2=1.905
r162 11 26 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.5 $Y=0.835
+ $X2=0.5 $Y2=1.575
r163 3 43 300 $w=1.7e-07 $l=7.74371e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.605 $X2=1.16 $Y2=3.275
r164 1 60 182 $w=1.7e-07 $l=2.96226e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.575 $X2=1.16 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%CK 3 6 10 11 13 16 18 19 22 25 26 31 33
+ 34 36 43 47 48 53
c146 36 0 1.35605e-19 $X=2.395 $Y=2.11
c147 34 0 1.65121e-19 $X=1.005 $Y=2.11
c148 22 0 4.60524e-20 $X=1.4 $Y=2.285
r149 48 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.545 $Y=2.11
+ $X2=1.4 $Y2=2.11
r150 47 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.25 $Y=2.11
+ $X2=2.395 $Y2=2.11
r151 47 48 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=2.25 $Y=2.11
+ $X2=1.545 $Y2=2.11
r152 43 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.4 $Y=2.11 $X2=1.4
+ $Y2=2.11
r153 43 45 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.4 $Y=2.11
+ $X2=1.4 $Y2=2.285
r154 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.395 $Y=2.11
+ $X2=2.395 $Y2=2.11
r155 36 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.395 $Y=2.11
+ $X2=2.395 $Y2=2.285
r156 33 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.11
+ $X2=1.4 $Y2=2.11
r157 33 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.315 $Y=2.11
+ $X2=1.005 $Y2=2.11
r158 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.92 $Y=2.025
+ $X2=1.005 $Y2=2.11
r159 29 31 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.92 $Y=2.025
+ $X2=0.92 $Y2=1.37
r160 28 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=2.285 $X2=2.395 $Y2=2.285
r161 25 26 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.277 $Y=1.205
+ $X2=2.277 $Y2=1.355
r162 22 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=2.285 $X2=1.4 $Y2=2.285
r163 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=2.285
+ $X2=1.4 $Y2=2.45
r164 18 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.92
+ $Y=1.37 $X2=0.92 $Y2=1.37
r165 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.37
+ $X2=0.92 $Y2=1.205
r166 16 28 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=2.305 $Y=2.12
+ $X2=2.352 $Y2=2.285
r167 16 26 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.305 $Y=2.12
+ $X2=2.305 $Y2=1.355
r168 11 28 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=2.25 $Y=2.45
+ $X2=2.352 $Y2=2.285
r169 11 13 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.25 $Y=2.45
+ $X2=2.25 $Y2=3.235
r170 10 25 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.25 $Y=0.835
+ $X2=2.25 $Y2=1.205
r171 6 24 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.46 $Y=3.235
+ $X2=1.46 $Y2=2.45
r172 3 19 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.86 $Y=0.835
+ $X2=0.86 $Y2=1.205
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%A_157_349# 1 3 11 13 14 17 20 25 31 35
+ 40 44 48 51 55 56
c136 56 0 1.35605e-19 $X=2.32 $Y=1.74
c137 55 0 3.47982e-21 $X=2.465 $Y=1.74
c138 51 0 4.60524e-20 $X=1.545 $Y=1.725
c139 20 0 1.24842e-20 $X=1.4 $Y=1.74
r140 55 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.465 $Y=1.74
+ $X2=2.32 $Y2=1.74
r141 51 53 0.0981889 $w=2.26e-07 $l=1.52315e-07 $layer=MET1_cond $X=1.545
+ $Y=1.725 $X2=1.4 $Y2=1.74
r142 51 56 0.959157 $w=1.4e-07 $l=7.75e-07 $layer=MET1_cond $X=1.545 $Y=1.725
+ $X2=2.32 $Y2=1.725
r143 46 48 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.465 $Y=2.705
+ $X2=2.735 $Y2=2.705
r144 43 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.465 $Y=1.74
+ $X2=2.465 $Y2=1.74
r145 43 44 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=2.465 $Y=1.725
+ $X2=2.735 $Y2=1.725
r146 40 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.62
+ $X2=2.735 $Y2=2.705
r147 39 44 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.735 $Y=1.825
+ $X2=2.735 $Y2=1.725
r148 39 40 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.735 $Y=1.825
+ $X2=2.735 $Y2=2.62
r149 35 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.465 $Y=2.935
+ $X2=2.465 $Y2=3.615
r150 33 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=2.79
+ $X2=2.465 $Y2=2.705
r151 33 35 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.465 $Y=2.79
+ $X2=2.465 $Y2=2.935
r152 29 43 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.465 $Y=1.625
+ $X2=2.465 $Y2=1.725
r153 29 31 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.465 $Y=1.625
+ $X2=2.465 $Y2=0.74
r154 25 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.4 $Y=1.74 $X2=1.4
+ $Y2=1.74
r155 20 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=1.74 $X2=1.4 $Y2=1.74
r156 20 22 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=1.4 $Y=1.74 $X2=1.4
+ $Y2=1.825
r157 20 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.74
+ $X2=1.4 $Y2=1.575
r158 17 21 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.46 $Y=0.835
+ $X2=1.46 $Y2=1.575
r159 13 22 15.0071 $w=1.6e-07 $l=1.35e-07 $layer=POLY_cond $X=1.265 $Y=1.825
+ $X2=1.4 $Y2=1.825
r160 13 14 152.942 $w=1.6e-07 $l=3.3e-07 $layer=POLY_cond $X=1.265 $Y=1.825
+ $X2=0.935 $Y2=1.825
r161 9 14 26.9672 $w=1.6e-07 $l=1.11355e-07 $layer=POLY_cond $X=0.86 $Y=1.905
+ $X2=0.935 $Y2=1.825
r162 9 11 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.86 $Y=1.905
+ $X2=0.86 $Y2=3.235
r163 3 37 400 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=2.605 $X2=2.465 $Y2=3.615
r164 3 35 400 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=2.605 $X2=2.465 $Y2=2.935
r165 1 31 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%A_349_89# 1 3 11 15 17 21 25 28 31 32 35
+ 37 41 45 51 56 57 58 60 61 62 67
c167 67 0 7.28655e-20 $X=4.035 $Y=1.74
c168 61 0 1.62658e-19 $X=3.9 $Y=1.74
c169 35 0 1.5259e-19 $X=1.882 $Y=1.812
c170 25 0 1.33411e-19 $X=4.15 $Y=3.445
r171 61 67 0.0969593 $w=2.3e-07 $l=1.35e-07 $layer=MET1_cond $X=3.9 $Y=1.74
+ $X2=4.035 $Y2=1.74
r172 61 62 0.962882 $w=1.7e-07 $l=1e-06 $layer=MET1_cond $X=3.9 $Y=1.74 $X2=2.9
+ $Y2=1.74
r173 59 62 0.0704148 $w=1.7e-07 $l=1.15888e-07 $layer=MET1_cond $X=2.827
+ $Y=1.825 $X2=2.9 $Y2=1.74
r174 59 60 0.664026 $w=1.45e-07 $l=5.7e-07 $layer=MET1_cond $X=2.827 $Y=1.825
+ $X2=2.827 $Y2=2.395
r175 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.025 $Y=2.48
+ $X2=1.88 $Y2=2.48
r176 57 60 0.0704148 $w=1.7e-07 $l=1.15521e-07 $layer=MET1_cond $X=2.755 $Y=2.48
+ $X2=2.827 $Y2=2.395
r177 57 58 0.702904 $w=1.7e-07 $l=7.3e-07 $layer=MET1_cond $X=2.755 $Y=2.48
+ $X2=2.025 $Y2=2.48
r178 51 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.035 $Y=1.74
+ $X2=4.035 $Y2=1.74
r179 49 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=1.74
+ $X2=3.415 $Y2=1.74
r180 49 51 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.5 $Y=1.74
+ $X2=4.035 $Y2=1.74
r181 45 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.415 $Y=2.935
+ $X2=3.415 $Y2=3.615
r182 43 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.825
+ $X2=3.415 $Y2=1.74
r183 43 45 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.415 $Y=1.825
+ $X2=3.415 $Y2=2.935
r184 39 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.655
+ $X2=3.415 $Y2=1.74
r185 39 41 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.415 $Y=1.655
+ $X2=3.415 $Y2=0.74
r186 37 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.88 $Y=2.48
+ $X2=1.88 $Y2=2.48
r187 35 55 5.01943 $w=1.75e-07 $l=7.2e-08 $layer=LI1_cond $X=1.882 $Y=1.812
+ $X2=1.882 $Y2=1.74
r188 35 37 42.3356 $w=1.73e-07 $l=6.68e-07 $layer=LI1_cond $X=1.882 $Y=1.812
+ $X2=1.882 $Y2=2.48
r189 34 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=1.74 $X2=4.035 $Y2=1.74
r190 31 32 43.105 $w=2e-07 $l=1.3e-07 $layer=POLY_cond $X=4.125 $Y=2.36
+ $X2=4.125 $Y2=2.49
r191 28 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.74 $X2=1.88 $Y2=1.74
r192 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.74
+ $X2=1.88 $Y2=1.905
r193 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.74
+ $X2=1.88 $Y2=1.575
r194 25 32 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=4.15 $Y=3.445
+ $X2=4.15 $Y2=2.49
r195 19 34 105.348 $w=2.27e-07 $l=5.12113e-07 $layer=POLY_cond $X=4.15 $Y=1.27
+ $X2=4.062 $Y2=1.74
r196 19 21 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.15 $Y=1.27
+ $X2=4.15 $Y2=0.755
r197 17 34 40.5863 $w=2.27e-07 $l=1.83016e-07 $layer=POLY_cond $X=4.1 $Y=1.905
+ $X2=4.062 $Y2=1.74
r198 17 31 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.1 $Y=1.905
+ $X2=4.1 $Y2=2.36
r199 15 30 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.82 $Y=3.235
+ $X2=1.82 $Y2=1.905
r200 11 29 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.82 $Y=0.835
+ $X2=1.82 $Y2=1.575
r201 3 47 400 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=2.605 $X2=3.415 $Y2=3.615
r202 3 45 400 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=2.605 $X2=3.415 $Y2=2.935
r203 1 41 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.575 $X2=3.415 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%ON 1 3 11 15 18 23 25 27 29 30 31 34 38
+ 41 43
c75 25 0 1.62658e-19 $X=3.935 $Y=2.195
c76 18 0 7.28655e-20 $X=4.52 $Y=2.015
r77 40 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=2.11
+ $X2=3.935 $Y2=2.11
r78 38 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.52 $Y=2.015
+ $X2=4.52 $Y2=1.745
r79 36 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=4.52 $Y=2.025
+ $X2=4.52 $Y2=2.015
r80 34 41 5.51377 $w=1.73e-07 $l=8.7e-08 $layer=LI1_cond $X=4.517 $Y=1.658
+ $X2=4.517 $Y2=1.745
r81 33 34 10.9642 $w=1.73e-07 $l=1.73e-07 $layer=LI1_cond $X=4.517 $Y=1.485
+ $X2=4.517 $Y2=1.658
r82 32 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.11
+ $X2=3.935 $Y2=2.11
r83 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=2.11
+ $X2=4.52 $Y2=2.025
r84 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=2.11
+ $X2=4.02 $Y2=2.11
r85 29 33 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.43 $Y=1.4
+ $X2=4.517 $Y2=1.485
r86 29 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.43 $Y=1.4 $X2=4.02
+ $Y2=1.4
r87 25 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=2.195
+ $X2=3.935 $Y2=2.11
r88 25 27 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=3.935 $Y=2.195
+ $X2=3.935 $Y2=3.615
r89 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=1.315
+ $X2=4.02 $Y2=1.4
r90 21 23 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.935 $Y=1.315
+ $X2=3.935 $Y2=0.74
r91 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=2.015 $X2=4.52 $Y2=2.015
r92 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.015
+ $X2=4.52 $Y2=2.18
r93 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.015
+ $X2=4.52 $Y2=1.85
r94 15 20 648.649 $w=1.5e-07 $l=1.265e-06 $layer=POLY_cond $X=4.58 $Y=3.445
+ $X2=4.58 $Y2=2.18
r95 11 19 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=4.58 $Y=0.755
+ $X2=4.58 $Y2=1.85
r96 3 27 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=3.025 $X2=3.935 $Y2=3.615
r97 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.81
+ $Y=0.575 $X2=3.935 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DLAT_L%Q 1 3 11 15 20 22 23 26
c21 26 0 1.33411e-19 $X=4.795 $Y=2.48
r22 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.795 $Y=2.48
+ $X2=4.795 $Y2=2.48
r23 22 24 5.06963 $w=2.33e-07 $l=8.5e-08 $layer=LI1_cond $X=4.827 $Y=2.48
+ $X2=4.827 $Y2=2.565
r24 22 23 5.06963 $w=2.33e-07 $l=8.5e-08 $layer=LI1_cond $X=4.827 $Y=2.48
+ $X2=4.827 $Y2=2.395
r25 20 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.86 $Y=1.145
+ $X2=4.86 $Y2=2.395
r26 19 20 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.827 $Y=0.975
+ $X2=4.827 $Y2=1.145
r27 15 24 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=4.795 $Y=3.615
+ $X2=4.795 $Y2=2.565
r28 11 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.795 $Y=0.74
+ $X2=4.795 $Y2=0.975
r29 3 15 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=4.655
+ $Y=3.025 $X2=4.795 $Y2=3.615
r30 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.575 $X2=4.795 $Y2=0.74
.ends

