* File: sky130_osu_sc_18T_ls__aoi22_l.pex.spice
* Created: Fri Nov 12 14:14:30 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%GND 1 2 27 31 33 44 56 58
c44 27 0 6.36774e-20 $X=-0.045 $Y=0
r45 56 58 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r46 42 52 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.152
r47 42 44 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.825
r48 33 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=0.152
+ $X2=1.91 $Y2=0.152
r49 29 31 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r50 27 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r51 27 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r52 27 29 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r53 27 34 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r54 27 33 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.825 $Y2=0.152
r55 27 34 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r56 2 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.77
+ $Y=0.575 $X2=1.91 $Y2=0.825
r57 1 31 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%VDD 1 17 19 26 34 39 43
r30 39 43 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r31 34 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.47 $X2=1.7
+ $Y2=6.47
r32 32 34 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r33 30 37 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r34 30 32 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r35 26 29 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=4.475
+ $X2=0.69 $Y2=5.835
r36 24 37 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r37 24 29 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r38 21 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r39 19 37 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r40 19 21 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r41 17 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r42 17 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r43 17 21 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r44 1 29 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r45 1 26 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%A0 2 3 5 8 12 18 21 27
c35 8 0 6.36774e-20 $X=0.475 $Y=4.585
r36 24 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=3.33
+ $X2=0.385 $Y2=3.33
r37 21 24 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.385 $Y=2.765
+ $X2=0.385 $Y2=3.33
r38 17 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.765 $X2=0.385 $Y2=2.765
r39 17 18 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.765
+ $X2=0.475 $Y2=2.765
r40 14 17 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.765
+ $X2=0.385 $Y2=2.765
r41 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.77
+ $X2=0.475 $Y2=1.77
r42 6 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=2.765
r43 6 8 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=4.585
r44 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.69 $X2=0.475
+ $Y2=1.77
r45 3 5 197.62 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.475 $Y=1.69
+ $X2=0.475 $Y2=1.075
r46 2 14 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.63
+ $X2=0.295 $Y2=2.765
r47 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.85 $X2=0.295
+ $Y2=1.77
r48 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.85
+ $X2=0.295 $Y2=2.63
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%A1 3 5 7 12 18
r43 15 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.96
+ $X2=0.725 $Y2=2.96
r44 12 15 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.725 $Y=2.255
+ $X2=0.725 $Y2=2.96
r45 10 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=2.255 $X2=0.725 $Y2=2.255
r46 5 10 63.0864 $w=2.95e-07 $l=3.7229e-07 $layer=POLY_cond $X=0.905 $Y=2.57
+ $X2=0.78 $Y2=2.255
r47 5 7 1033.22 $w=1.5e-07 $l=2.015e-06 $layer=POLY_cond $X=0.905 $Y=2.57
+ $X2=0.905 $Y2=4.585
r48 1 10 38.578 $w=2.95e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.835 $Y=2.09
+ $X2=0.78 $Y2=2.255
r49 1 3 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=0.835 $Y=2.09
+ $X2=0.835 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%B0 3 7 10 15 17 21
r44 17 19 3.63576 $w=3.02e-07 $l=9e-08 $layer=LI1_cond $X=1.165 $Y=1.9 $X2=1.255
+ $Y2=1.9
r45 15 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.59
+ $X2=1.165 $Y2=2.59
r46 13 17 4.10007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=2.065
+ $X2=1.165 $Y2=1.9
r47 13 15 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.165 $Y=2.065
+ $X2=1.165 $Y2=2.59
r48 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.9 $X2=1.255 $Y2=1.9
r49 10 12 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.9
+ $X2=1.265 $Y2=2.065
r50 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.9
+ $X2=1.265 $Y2=1.735
r51 7 12 1292.17 $w=1.5e-07 $l=2.52e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.065
r52 3 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=1.735
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%B1 3 7 10 14 19
r26 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.935 $Y=2.225
+ $X2=1.935 $Y2=2.225
r27 12 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=2.225 $X2=1.935 $Y2=2.225
r28 10 12 26.0127 $w=3.15e-07 $l=1.7e-07 $layer=POLY_cond $X=1.765 $Y=2.205
+ $X2=1.935 $Y2=2.205
r29 9 10 10.7111 $w=3.15e-07 $l=7e-08 $layer=POLY_cond $X=1.695 $Y=2.205
+ $X2=1.765 $Y2=2.205
r30 5 10 20.1192 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.765 $Y=2.39
+ $X2=1.765 $Y2=2.205
r31 5 7 1125.52 $w=1.5e-07 $l=2.195e-06 $layer=POLY_cond $X=1.765 $Y=2.39
+ $X2=1.765 $Y2=4.585
r32 1 9 20.1192 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.695 $Y=2.02
+ $X2=1.695 $Y2=2.205
r33 1 3 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.695 $Y=2.02
+ $X2=1.695 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%A_27_617# 1 2 3 15 19 20 27 28
r23 31 34 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=5.835
r24 29 34 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.98 $Y=5.915 $X2=1.98
+ $Y2=5.835
r25 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.895 $Y=6
+ $X2=1.98 $Y2=5.915
r26 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=6 $X2=1.205
+ $Y2=6
r27 24 26 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=5.835
r28 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=5.915
+ $X2=1.205 $Y2=6
r29 22 26 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=5.915 $X2=1.12
+ $Y2=5.835
r30 21 24 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=4.055 $X2=1.12
+ $Y2=4.135
r31 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.97
+ $X2=1.12 $Y2=4.055
r32 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.97
+ $X2=0.345 $Y2=3.97
r33 15 17 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r34 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=4.055
+ $X2=0.345 $Y2=3.97
r35 13 15 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=4.055 $X2=0.26
+ $Y2=4.135
r36 3 34 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r37 3 31 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=4.135
r38 2 26 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r39 2 24 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=4.135
r40 1 17 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r41 1 15 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%Y 1 3 10 17 23 27 28 32 38
c40 32 0 5.84789e-20 $X=1.605 $Y=1.7
r41 38 39 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.595 $Y=1.85
+ $X2=1.595 $Y2=1.735
r42 32 39 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.605 $Y=1.7
+ $X2=1.605 $Y2=1.735
r43 29 32 0.129989 $w=1.7e-07 $l=1.35e-07 $layer=MET1_cond $X=1.605 $Y=1.565
+ $X2=1.605 $Y2=1.7
r44 28 35 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.23 $Y=1.48
+ $X2=1.085 $Y2=1.48
r45 27 29 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.52 $Y=1.48
+ $X2=1.605 $Y2=1.565
r46 27 28 0.279236 $w=1.7e-07 $l=2.9e-07 $layer=MET1_cond $X=1.52 $Y=1.48
+ $X2=1.23 $Y2=1.48
r47 25 26 9.11234 $w=2.13e-07 $l=1.7e-07 $layer=LI1_cond $X=1.572 $Y=3.16
+ $X2=1.572 $Y2=3.33
r48 23 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.595 $Y=1.85
+ $X2=1.595 $Y2=1.85
r49 23 25 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.595 $Y=1.85
+ $X2=1.595 $Y2=3.16
r50 17 19 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=5.495
r51 17 26 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=3.33
r52 13 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=1.48
+ $X2=1.085 $Y2=1.48
r53 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.085 $Y=0.825
+ $X2=1.085 $Y2=1.48
r54 3 19 240 $w=1.7e-07 $l=2.47901e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.495
r55 3 17 240 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=4.135
r56 1 10 91 $w=1.7e-07 $l=3.2596e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.085 $Y2=0.825
.ends

