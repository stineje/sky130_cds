magic
tech sky130A
magscale 1 2
timestamp 1646761201
<< checkpaint >>
rect -1529 2461 2577 2597
rect -1760 -1129 6260 2461
rect -1529 -1260 2577 -1129
<< nwell >>
rect 0 1084 255 1085
rect -269 711 1317 1084
rect -269 524 1310 711
<< nmoslvt >>
rect -180 110 -150 258
rect -94 110 -64 258
rect 96 110 126 258
rect 182 110 212 258
rect 254 110 284 258
rect 374 110 404 258
rect 446 110 476 258
rect 532 110 562 258
rect 740 110 770 258
rect 826 110 856 258
rect 1016 110 1046 258
rect 1102 110 1132 258
rect 1188 110 1218 258
<< pmos >>
rect -180 560 -150 960
rect -108 560 -78 960
rect 96 560 126 960
rect 182 560 212 960
rect 254 560 284 960
rect 374 560 404 960
rect 446 560 476 960
rect 532 560 562 960
rect 740 560 770 960
rect 826 560 856 960
rect 1016 560 1046 960
rect 1102 560 1132 960
rect 1188 560 1218 960
<< ndiff >>
rect -233 210 -180 258
rect -233 126 -225 210
rect -191 126 -180 210
rect -233 110 -180 126
rect -150 210 -94 258
rect -150 126 -139 210
rect -105 126 -94 210
rect -150 110 -94 126
rect -64 210 -11 258
rect -64 126 -53 210
rect -19 126 -11 210
rect -64 110 -11 126
rect 43 210 96 258
rect 43 126 51 210
rect 85 126 96 210
rect 43 110 96 126
rect 126 210 182 258
rect 126 126 137 210
rect 171 126 182 210
rect 126 110 182 126
rect 212 110 254 258
rect 284 210 374 258
rect 284 126 295 210
rect 363 126 374 210
rect 284 110 374 126
rect 404 110 446 258
rect 476 210 532 258
rect 476 126 487 210
rect 521 126 532 210
rect 476 110 532 126
rect 562 210 615 258
rect 562 126 573 210
rect 607 126 615 210
rect 562 110 615 126
rect 687 210 740 258
rect 687 126 695 210
rect 729 126 740 210
rect 687 110 740 126
rect 770 210 826 258
rect 770 126 781 210
rect 815 126 826 210
rect 770 110 826 126
rect 856 210 909 258
rect 856 126 867 210
rect 901 126 909 210
rect 856 110 909 126
rect 963 210 1016 258
rect 963 126 971 210
rect 1005 126 1016 210
rect 963 110 1016 126
rect 1046 210 1102 258
rect 1046 126 1057 210
rect 1091 126 1102 210
rect 1046 110 1102 126
rect 1132 210 1188 258
rect 1132 126 1143 210
rect 1177 126 1188 210
rect 1132 110 1188 126
rect 1218 210 1271 258
rect 1218 126 1229 210
rect 1263 126 1271 210
rect 1218 110 1271 126
<< pdiff >>
rect -233 949 -180 960
rect -233 600 -225 949
rect -191 600 -180 949
rect -233 560 -180 600
rect -150 560 -108 960
rect -78 949 -25 960
rect -78 736 -67 949
rect -33 736 -25 949
rect -78 560 -25 736
rect 43 949 96 960
rect 43 668 51 949
rect 85 668 96 949
rect 43 560 96 668
rect 126 949 182 960
rect 126 668 137 949
rect 171 668 182 949
rect 126 560 182 668
rect 212 560 254 960
rect 284 949 374 960
rect 284 600 295 949
rect 363 600 374 949
rect 284 560 374 600
rect 404 560 446 960
rect 476 949 532 960
rect 476 600 487 949
rect 521 600 532 949
rect 476 560 532 600
rect 562 949 615 960
rect 562 600 573 949
rect 607 600 615 949
rect 562 560 615 600
rect 687 949 740 960
rect 687 600 695 949
rect 729 600 740 949
rect 687 560 740 600
rect 770 949 826 960
rect 770 600 781 949
rect 815 600 826 949
rect 770 560 826 600
rect 856 949 909 960
rect 856 600 867 949
rect 901 600 909 949
rect 856 560 909 600
rect 963 949 1016 960
rect 963 668 971 949
rect 1005 668 1016 949
rect 963 560 1016 668
rect 1046 560 1102 960
rect 1132 949 1188 960
rect 1132 736 1143 949
rect 1177 736 1188 949
rect 1132 560 1188 736
rect 1218 949 1271 960
rect 1218 600 1229 949
rect 1263 600 1271 949
rect 1218 560 1271 600
<< ndiffc >>
rect -225 126 -191 210
rect -139 126 -105 210
rect -53 126 -19 210
rect 51 126 85 210
rect 137 126 171 210
rect 295 126 363 210
rect 487 126 521 210
rect 573 126 607 210
rect 695 126 729 210
rect 781 126 815 210
rect 867 126 901 210
rect 971 126 1005 210
rect 1057 126 1091 210
rect 1143 126 1177 210
rect 1229 126 1263 210
<< pdiffc >>
rect -225 600 -191 949
rect -67 736 -33 949
rect 51 668 85 949
rect 137 668 171 949
rect 295 600 363 949
rect 487 600 521 949
rect 573 600 607 949
rect 695 600 729 949
rect 781 600 815 949
rect 867 600 901 949
rect 971 668 1005 949
rect 1143 736 1177 949
rect 1229 600 1263 949
<< psubdiff >>
rect -233 22 -209 56
rect -175 22 -151 56
rect -97 22 -73 56
rect -39 22 -15 56
rect 88 22 112 56
rect 146 22 170 56
rect 224 22 248 56
rect 282 22 306 56
rect 360 22 384 56
rect 418 22 442 56
rect 496 22 520 56
rect 554 22 578 56
rect 632 22 656 56
rect 690 22 714 56
rect 768 22 792 56
rect 826 22 850 56
rect 963 22 987 56
rect 1021 22 1045 56
rect 1099 22 1123 56
rect 1157 22 1181 56
<< nsubdiff >>
rect -233 1014 -209 1048
rect -175 1014 -151 1048
rect -97 1014 -73 1048
rect -39 1014 -15 1048
rect 88 1014 112 1048
rect 146 1014 170 1048
rect 224 1014 248 1048
rect 282 1014 306 1048
rect 360 1014 384 1048
rect 418 1014 442 1048
rect 496 1014 520 1048
rect 554 1014 578 1048
rect 632 1014 656 1048
rect 690 1014 714 1048
rect 768 1014 792 1048
rect 826 1014 850 1048
rect 963 1014 987 1048
rect 1021 1014 1045 1048
rect 1099 1014 1123 1048
rect 1157 1014 1181 1048
<< psubdiffcont >>
rect -209 22 -175 56
rect -73 22 -39 56
rect 112 22 146 56
rect 248 22 282 56
rect 384 22 418 56
rect 520 22 554 56
rect 656 22 690 56
rect 792 22 826 56
rect 987 22 1021 56
rect 1123 22 1157 56
<< nsubdiffcont >>
rect -209 1014 -175 1048
rect -73 1014 -39 1048
rect 112 1014 146 1048
rect 248 1014 282 1048
rect 384 1014 418 1048
rect 520 1014 554 1048
rect 656 1014 690 1048
rect 792 1014 826 1048
rect 987 1014 1021 1048
rect 1123 1014 1157 1048
<< poly >>
rect -180 960 -150 986
rect -108 960 -78 986
rect 96 960 126 986
rect 182 960 212 986
rect 254 960 284 986
rect 374 960 404 986
rect 446 960 476 986
rect 532 960 562 986
rect 740 960 770 986
rect 826 960 856 986
rect 1016 960 1046 986
rect 1102 960 1132 986
rect 1188 960 1218 986
rect -180 394 -150 560
rect -108 527 -78 560
rect 96 538 126 560
rect -108 511 -35 527
rect -108 477 -79 511
rect -45 477 -35 511
rect -108 461 -35 477
rect 86 504 126 538
rect -204 378 -150 394
rect -204 344 -194 378
rect -160 344 -150 378
rect -204 328 -150 344
rect -180 258 -150 328
rect -94 258 -64 461
rect 86 346 116 504
rect 182 461 212 560
rect 254 529 284 560
rect 374 529 404 560
rect 254 513 308 529
rect 254 479 264 513
rect 298 479 308 513
rect 254 463 308 479
rect 350 513 404 529
rect 350 479 360 513
rect 394 479 404 513
rect 350 463 404 479
rect 158 445 212 461
rect 158 411 168 445
rect 202 411 212 445
rect 350 418 380 463
rect 158 395 212 411
rect 86 330 140 346
rect 86 296 96 330
rect 130 296 140 330
rect 86 280 140 296
rect 96 258 126 280
rect 182 258 212 395
rect 254 388 380 418
rect 446 420 476 560
rect 532 529 562 560
rect 740 544 770 560
rect 532 513 603 529
rect 532 499 559 513
rect 543 479 559 499
rect 593 479 603 513
rect 543 463 603 479
rect 730 514 770 544
rect 446 404 500 420
rect 254 258 284 388
rect 446 370 456 404
rect 490 370 500 404
rect 446 354 500 370
rect 350 330 404 346
rect 350 296 360 330
rect 394 296 404 330
rect 350 280 404 296
rect 374 258 404 280
rect 446 258 476 354
rect 543 306 573 463
rect 730 420 760 514
rect 826 420 856 560
rect 1016 511 1046 560
rect 963 495 1046 511
rect 963 461 973 495
rect 1007 461 1046 495
rect 963 445 1046 461
rect 1102 453 1132 560
rect 1188 535 1218 560
rect 1188 505 1225 535
rect 705 404 760 420
rect 705 370 715 404
rect 749 370 760 404
rect 705 354 760 370
rect 802 404 856 420
rect 802 370 812 404
rect 846 370 856 404
rect 802 354 856 370
rect 532 276 573 306
rect 730 303 760 354
rect 532 258 562 276
rect 730 273 770 303
rect 740 258 770 273
rect 826 258 856 354
rect 1016 258 1046 445
rect 1099 437 1153 453
rect 1099 403 1109 437
rect 1143 403 1153 437
rect 1099 387 1153 403
rect 1102 258 1132 387
rect 1195 363 1225 505
rect 1195 347 1249 363
rect 1195 327 1205 347
rect 1188 313 1205 327
rect 1239 313 1249 347
rect 1188 297 1249 313
rect 1188 258 1218 297
rect -180 84 -150 110
rect -94 84 -64 110
rect 96 84 126 110
rect 182 84 212 110
rect 254 84 284 110
rect 374 84 404 110
rect 446 84 476 110
rect 532 84 562 110
rect 740 84 770 110
rect 826 84 856 110
rect 1016 84 1046 110
rect 1102 84 1132 110
rect 1188 84 1218 110
<< polycont >>
rect -79 477 -45 511
rect -194 344 -160 378
rect 264 479 298 513
rect 360 479 394 513
rect 168 411 202 445
rect 96 296 130 330
rect 559 479 593 513
rect 456 370 490 404
rect 360 296 394 330
rect 973 461 1007 495
rect 715 370 749 404
rect 812 370 846 404
rect 1109 403 1143 437
rect 1205 313 1239 347
<< locali >>
rect -267 1054 1317 1075
rect -267 1014 -209 1054
rect -175 1014 -73 1054
rect -39 1014 112 1054
rect 146 1014 248 1054
rect 282 1014 384 1054
rect 418 1014 520 1054
rect 554 1014 656 1054
rect 690 1014 792 1054
rect 826 1014 987 1054
rect 1021 1014 1123 1054
rect 1157 1014 1317 1054
rect -225 949 -191 960
rect -67 949 -33 1014
rect -67 720 -33 736
rect 51 949 85 960
rect 28 668 51 734
rect 28 651 85 668
rect 137 949 171 1014
rect 137 652 171 668
rect 295 949 363 960
rect -225 478 -191 600
rect -147 378 -113 518
rect -79 511 -45 592
rect -79 461 -45 477
rect -210 344 -194 378
rect -160 344 -113 378
rect 28 404 62 651
rect 295 597 363 600
rect -225 210 -191 226
rect -225 56 -191 126
rect 28 239 62 370
rect 96 563 363 597
rect 487 949 521 1014
rect 487 584 521 600
rect 573 949 607 960
rect 573 597 607 600
rect 695 949 729 960
rect 573 563 661 597
rect 96 330 130 563
rect 360 513 394 529
rect 248 479 264 513
rect 298 479 314 513
rect 168 395 202 411
rect 280 330 314 479
rect 360 478 394 479
rect 559 513 593 529
rect 559 478 593 479
rect 627 404 661 563
rect 695 552 729 600
rect 781 949 815 1014
rect 781 584 815 600
rect 867 949 901 960
rect 971 949 1005 960
rect 1143 949 1177 1014
rect 1143 720 1177 736
rect 1229 949 1263 960
rect 1005 668 1075 686
rect 971 652 1075 668
rect 901 592 914 609
rect 867 575 914 592
rect 695 513 729 518
rect 695 479 846 513
rect 812 404 846 479
rect 440 370 456 404
rect 490 370 506 404
rect 573 370 661 404
rect 699 370 715 404
rect 749 370 765 404
rect 573 330 607 370
rect 812 330 846 370
rect 130 296 239 330
rect 280 296 360 330
rect 394 296 607 330
rect 96 280 130 296
rect 205 246 239 296
rect -139 210 -105 222
rect -139 110 -105 126
rect -53 210 -19 226
rect 28 210 85 239
rect 28 205 51 210
rect -53 56 -19 126
rect 51 110 85 126
rect 137 210 171 226
rect 205 212 363 246
rect 137 56 171 126
rect 295 210 363 212
rect 295 110 363 126
rect 487 210 521 226
rect 487 56 521 126
rect 573 210 607 296
rect 573 110 607 126
rect 695 296 846 330
rect 695 210 729 296
rect 880 262 914 575
rect 973 495 1007 518
rect 973 445 1007 461
rect 1041 347 1075 652
rect 1109 478 1143 592
rect 1229 478 1263 600
rect 1109 437 1143 444
rect 1109 387 1143 403
rect 1041 313 1205 347
rect 1239 313 1255 347
rect 867 228 914 262
rect 695 110 729 126
rect 781 210 815 226
rect 781 56 815 126
rect 867 210 901 228
rect 867 110 901 126
rect 971 210 1005 226
rect 971 56 1005 126
rect 1057 210 1091 313
rect 1057 110 1091 126
rect 1143 210 1177 226
rect 1143 56 1177 126
rect 1229 210 1263 222
rect 1229 110 1263 126
rect -267 16 -209 56
rect -175 16 -73 56
rect -39 16 112 56
rect 146 16 248 56
rect 282 16 384 56
rect 418 16 520 56
rect 554 16 656 56
rect 690 16 792 56
rect 826 16 987 56
rect 1021 16 1123 56
rect 1157 16 1317 56
rect -267 -5 1317 16
<< viali >>
rect -209 1048 -175 1054
rect -209 1020 -175 1048
rect -73 1048 -39 1054
rect -73 1020 -39 1048
rect 112 1048 146 1054
rect 112 1020 146 1048
rect 248 1048 282 1054
rect 248 1020 282 1048
rect 384 1048 418 1054
rect 384 1020 418 1048
rect 520 1048 554 1054
rect 520 1020 554 1048
rect 656 1048 690 1054
rect 656 1020 690 1048
rect 792 1048 826 1054
rect 792 1020 826 1048
rect 987 1048 1021 1054
rect 987 1020 1021 1048
rect 1123 1048 1157 1054
rect 1123 1020 1157 1048
rect -79 592 -45 626
rect -225 444 -191 478
rect -147 518 -113 552
rect 28 370 62 404
rect -139 222 -105 256
rect 168 445 202 479
rect 360 444 394 478
rect 559 444 593 478
rect 867 600 901 626
rect 867 592 901 600
rect 695 518 729 552
rect 456 370 490 404
rect 715 370 749 404
rect 973 518 1007 552
rect 1109 592 1143 626
rect 1109 444 1143 478
rect 1229 444 1263 478
rect 1229 222 1263 256
rect -209 22 -175 50
rect -209 16 -175 22
rect -73 22 -39 50
rect -73 16 -39 22
rect 112 22 146 50
rect 112 16 146 22
rect 248 22 282 50
rect 248 16 282 22
rect 384 22 418 50
rect 384 16 418 22
rect 520 22 554 50
rect 520 16 554 22
rect 656 22 690 50
rect 656 16 690 22
rect 792 22 826 50
rect 792 16 826 22
rect 987 22 1021 50
rect 987 16 1021 22
rect 1123 22 1157 50
rect 1123 16 1157 22
<< metal1 >>
rect -267 1054 1317 1075
rect -267 1020 -209 1054
rect -175 1020 -73 1054
rect -39 1020 112 1054
rect 146 1020 248 1054
rect 282 1020 384 1054
rect 418 1020 520 1054
rect 554 1020 656 1054
rect 690 1020 792 1054
rect 826 1020 987 1054
rect 1021 1020 1123 1054
rect 1157 1020 1317 1054
rect -267 1014 1317 1020
rect -91 626 -33 632
rect 855 626 913 632
rect 1097 629 1155 632
rect -112 592 -79 626
rect -45 592 -33 626
rect 832 592 867 626
rect 901 592 913 626
rect -91 586 -33 592
rect 855 586 913 592
rect 1078 626 1155 629
rect 1078 592 1109 626
rect 1143 592 1155 626
rect 1078 591 1155 592
rect 1097 586 1155 591
rect -159 552 -101 558
rect 683 552 741 558
rect -181 518 -147 552
rect -113 518 -101 552
rect 676 551 695 552
rect 661 519 695 551
rect 676 518 695 519
rect 729 518 741 552
rect 867 552 901 586
rect 961 552 1019 558
rect 867 518 973 552
rect 1007 518 1041 552
rect -159 512 -101 518
rect 683 512 741 518
rect 961 512 1019 518
rect -237 478 -179 484
rect 156 479 215 485
rect 156 478 168 479
rect -237 444 -225 478
rect -191 445 168 478
rect 202 445 235 479
rect 348 478 406 484
rect 547 478 605 484
rect 1097 478 1155 484
rect -191 444 215 445
rect -237 438 -179 444
rect -139 262 -105 444
rect 156 439 215 444
rect 348 444 360 478
rect 394 444 559 478
rect 593 444 609 478
rect 1076 444 1109 478
rect 1143 444 1155 478
rect 348 438 406 444
rect 547 438 605 444
rect 1097 438 1155 444
rect 1217 478 1275 484
rect 1217 444 1229 478
rect 1263 444 1275 478
rect 1217 438 1275 444
rect 15 404 74 410
rect 15 370 28 404
rect 62 397 74 404
rect 444 404 503 410
rect 444 397 456 404
rect 62 370 456 397
rect 490 401 503 404
rect 703 404 761 410
rect 703 401 715 404
rect 490 373 715 401
rect 490 370 503 373
rect 15 369 503 370
rect 15 364 74 369
rect 444 364 503 369
rect 703 370 715 373
rect 749 370 761 404
rect 703 364 761 370
rect 1229 262 1263 438
rect -151 256 -93 262
rect -151 222 -139 256
rect -105 222 -93 256
rect -151 216 -93 222
rect 1217 256 1275 262
rect 1217 222 1229 256
rect 1263 222 1275 256
rect 1217 216 1275 222
rect -267 50 1317 56
rect -267 16 -209 50
rect -175 16 -73 50
rect -39 16 112 50
rect 146 16 248 50
rect 282 16 384 50
rect 418 16 520 50
rect 554 16 656 50
rect 690 16 792 50
rect 826 16 987 50
rect 1021 16 1123 50
rect 1157 16 1317 50
rect -267 -5 1317 16
<< labels >>
rlabel viali -130 535 -130 535 1 SE
rlabel viali -61 608 -61 608 1 E
rlabel viali 576 461 576 461 1 CK
rlabel viali 1246 461 1246 461 1 ECK
rlabel viali 712 535 712 535 1 Q
rlabel viali 1125 462 1125 462 1 CKa
rlabel nwell -191 1035 -190 1035 1 vdd
rlabel nwell -56 1036 -55 1036 1 vdd
rlabel nwell 129 1036 130 1036 1 vdd
rlabel viali 264 1035 264 1035 1 vdd
rlabel viali 401 1037 401 1037 1 vdd
rlabel viali 538 1037 538 1037 1 vdd
rlabel nwell 674 1037 674 1038 1 vdd
rlabel nwell 809 1038 809 1039 1 vdd
rlabel nwell 1004 1037 1004 1038 1 vdd
rlabel nwell 1141 1037 1141 1038 1 vdd
rlabel viali -192 36 -192 36 1 gnd
rlabel viali -56 34 -56 34 1 gnd
rlabel viali 129 34 129 34 1 gnd
rlabel viali 265 34 265 34 1 gnd
rlabel viali 400 35 400 35 1 gnd
rlabel viali 536 33 536 33 1 gnd
rlabel viali 673 33 673 33 1 gnd
rlabel viali 810 34 810 34 1 gnd
rlabel viali 1005 34 1005 34 1 gnd
rlabel viali 1139 35 1139 35 1 gnd
<< end >>
