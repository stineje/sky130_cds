* File: sky130_osu_sc_15T_hs__buf_4.pxi.spice
* Created: Fri Nov 12 14:28:17 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__BUF_4%GND N_GND_M1006_d N_GND_M1003_s N_GND_M1009_s
+ N_GND_M1006_b N_GND_c_2_p N_GND_c_12_p N_GND_c_21_p N_GND_c_3_p N_GND_c_27_p
+ GND N_GND_c_22_p PM_SKY130_OSU_SC_15T_HS__BUF_4%GND
x_PM_SKY130_OSU_SC_15T_HS__BUF_4%VDD N_VDD_M1007_d N_VDD_M1001_s N_VDD_M1005_s
+ N_VDD_M1007_b N_VDD_c_60_p N_VDD_c_61_p N_VDD_c_70_p N_VDD_c_75_p N_VDD_c_82_p
+ N_VDD_c_87_p VDD N_VDD_c_62_p PM_SKY130_OSU_SC_15T_HS__BUF_4%VDD
x_PM_SKY130_OSU_SC_15T_HS__BUF_4%A N_A_M1006_g N_A_M1007_g N_A_c_107_n
+ N_A_c_108_n A PM_SKY130_OSU_SC_15T_HS__BUF_4%A
x_PM_SKY130_OSU_SC_15T_HS__BUF_4%A_27_115# N_A_27_115#_M1006_s
+ N_A_27_115#_M1007_s N_A_27_115#_M1002_g N_A_27_115#_c_174_n
+ N_A_27_115#_M1000_g N_A_27_115#_c_145_n N_A_27_115#_M1003_g
+ N_A_27_115#_c_178_n N_A_27_115#_M1001_g N_A_27_115#_c_149_n
+ N_A_27_115#_c_151_n N_A_27_115#_c_152_n N_A_27_115#_c_153_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_186_n N_A_27_115#_M1004_g
+ N_A_27_115#_c_158_n N_A_27_115#_c_159_n N_A_27_115#_M1009_g
+ N_A_27_115#_c_191_n N_A_27_115#_M1005_g N_A_27_115#_c_164_n
+ N_A_27_115#_c_165_n N_A_27_115#_c_166_n N_A_27_115#_c_169_n
+ N_A_27_115#_c_170_n N_A_27_115#_c_172_n N_A_27_115#_c_173_n
+ PM_SKY130_OSU_SC_15T_HS__BUF_4%A_27_115#
x_PM_SKY130_OSU_SC_15T_HS__BUF_4%Y N_Y_M1002_d N_Y_M1008_d N_Y_M1000_d
+ N_Y_M1004_d N_Y_c_260_n N_Y_c_280_n N_Y_c_264_n N_Y_c_283_n N_Y_c_268_n
+ N_Y_c_271_n Y N_Y_c_273_n N_Y_c_287_n N_Y_c_276_n N_Y_c_279_n
+ PM_SKY130_OSU_SC_15T_HS__BUF_4%Y
cc_1 N_GND_M1006_b N_A_M1006_g 0.0645215f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_A_M1006_g 0.00388248f $X=0.69 $Y=0.865 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_A_M1006_g 0.00607478f $X=1.635 $Y=0.152 $X2=0.475 $Y2=0.895
cc_4 N_GND_M1006_b N_A_M1007_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_5 N_GND_M1006_b N_A_c_107_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.22
cc_6 N_GND_M1006_b N_A_c_108_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.22
cc_7 N_GND_M1006_b N_A_27_115#_M1002_g 0.0255945f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.895
cc_8 N_GND_c_2_p N_A_27_115#_M1002_g 0.00388248f $X=0.69 $Y=0.865 $X2=0.905
+ $Y2=0.895
cc_9 N_GND_c_3_p N_A_27_115#_M1002_g 0.00607478f $X=1.635 $Y=0.152 $X2=0.905
+ $Y2=0.895
cc_10 N_GND_M1006_b N_A_27_115#_c_145_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.6
cc_11 N_GND_M1006_b N_A_27_115#_M1003_g 0.024527f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.895
cc_12 N_GND_c_12_p N_A_27_115#_M1003_g 0.00390533f $X=1.55 $Y=0.865 $X2=1.335
+ $Y2=0.895
cc_13 N_GND_c_3_p N_A_27_115#_M1003_g 0.00607478f $X=1.635 $Y=0.152 $X2=1.335
+ $Y2=0.895
cc_14 N_GND_M1006_b N_A_27_115#_c_149_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.585
cc_15 N_GND_c_12_p N_A_27_115#_c_149_n 0.00256938f $X=1.55 $Y=0.865 $X2=1.69
+ $Y2=1.585
cc_16 N_GND_M1006_b N_A_27_115#_c_151_n 0.0479019f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.585
cc_17 N_GND_M1006_b N_A_27_115#_c_152_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.675
cc_18 N_GND_M1006_b N_A_27_115#_c_153_n 0.0244408f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.675
cc_19 N_GND_M1006_b N_A_27_115#_M1008_g 0.0245289f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.895
cc_20 N_GND_c_12_p N_A_27_115#_M1008_g 0.00390533f $X=1.55 $Y=0.865 $X2=1.765
+ $Y2=0.895
cc_21 N_GND_c_21_p N_A_27_115#_M1008_g 0.00606474f $X=2.325 $Y=0.152 $X2=1.765
+ $Y2=0.895
cc_22 N_GND_c_22_p N_A_27_115#_M1008_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765
+ $Y2=0.895
cc_23 N_GND_M1006_b N_A_27_115#_c_158_n 0.0385034f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_24 N_GND_M1006_b N_A_27_115#_c_159_n 0.0221499f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.675
cc_25 N_GND_M1006_b N_A_27_115#_M1009_g 0.0341369f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.895
cc_26 N_GND_c_21_p N_A_27_115#_M1009_g 0.00606474f $X=2.325 $Y=0.152 $X2=2.195
+ $Y2=0.895
cc_27 N_GND_c_27_p N_A_27_115#_M1009_g 0.00866533f $X=2.41 $Y=0.865 $X2=2.195
+ $Y2=0.895
cc_28 N_GND_c_22_p N_A_27_115#_M1009_g 0.00468827f $X=1.7 $Y=0.19 $X2=2.195
+ $Y2=0.895
cc_29 N_GND_M1006_b N_A_27_115#_c_164_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.585
cc_30 N_GND_M1006_b N_A_27_115#_c_165_n 0.00890086f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.675
cc_31 N_GND_M1006_b N_A_27_115#_c_166_n 0.0191786f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_32 N_GND_c_3_p N_A_27_115#_c_166_n 0.00895373f $X=1.635 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_33 N_GND_c_22_p N_A_27_115#_c_166_n 0.00136847f $X=1.7 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_34 N_GND_M1006_b N_A_27_115#_c_169_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.205
cc_35 N_GND_M1006_b N_A_27_115#_c_170_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.675
cc_36 N_GND_c_2_p N_A_27_115#_c_170_n 0.00702738f $X=0.69 $Y=0.865 $X2=0.88
+ $Y2=1.675
cc_37 N_GND_M1006_b N_A_27_115#_c_172_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.675
cc_38 N_GND_M1006_b N_A_27_115#_c_173_n 0.00592383f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.675
cc_39 N_GND_M1006_b N_Y_c_260_n 0.00643585f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.865
cc_40 N_GND_c_12_p N_Y_c_260_n 8.14297e-19 $X=1.55 $Y=0.865 $X2=1.12 $Y2=0.865
cc_41 N_GND_c_3_p N_Y_c_260_n 0.00893077f $X=1.635 $Y=0.152 $X2=1.12 $Y2=0.865
cc_42 N_GND_c_22_p N_Y_c_260_n 0.00136371f $X=1.7 $Y=0.19 $X2=1.12 $Y2=0.865
cc_43 N_GND_M1006_b N_Y_c_264_n 0.00656459f $X=-0.045 $Y=0 $X2=1.98 $Y2=0.865
cc_44 N_GND_c_12_p N_Y_c_264_n 8.14297e-19 $X=1.55 $Y=0.865 $X2=1.98 $Y2=0.865
cc_45 N_GND_c_21_p N_Y_c_264_n 0.00754406f $X=2.325 $Y=0.152 $X2=1.98 $Y2=0.865
cc_46 N_GND_c_22_p N_Y_c_264_n 0.00475776f $X=1.7 $Y=0.19 $X2=1.98 $Y2=0.865
cc_47 N_GND_M1006_b N_Y_c_268_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.335
cc_48 N_GND_c_2_p N_Y_c_268_n 0.00134236f $X=0.69 $Y=0.865 $X2=1.12 $Y2=1.335
cc_49 N_GND_c_12_p N_Y_c_268_n 7.53951e-19 $X=1.55 $Y=0.865 $X2=1.12 $Y2=1.335
cc_50 N_GND_M1006_b N_Y_c_271_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.585
cc_51 N_GND_M1006_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=2.01
cc_52 N_GND_M1003_s N_Y_c_273_n 0.00418405f $X=1.41 $Y=0.575 $X2=1.835 $Y2=1.22
cc_53 N_GND_M1006_b N_Y_c_273_n 0.00793787f $X=-0.045 $Y=0 $X2=1.835 $Y2=1.22
cc_54 N_GND_c_12_p N_Y_c_273_n 0.0142303f $X=1.55 $Y=0.865 $X2=1.835 $Y2=1.22
cc_55 N_GND_M1006_b N_Y_c_276_n 0.00409378f $X=-0.045 $Y=0 $X2=1.98 $Y2=1.335
cc_56 N_GND_c_12_p N_Y_c_276_n 7.53951e-19 $X=1.55 $Y=0.865 $X2=1.98 $Y2=1.335
cc_57 N_GND_c_27_p N_Y_c_276_n 0.00134236f $X=2.41 $Y=0.865 $X2=1.98 $Y2=1.335
cc_58 N_GND_M1006_b N_Y_c_279_n 0.0651512f $X=-0.045 $Y=0 $X2=1.98 $Y2=2.585
cc_59 N_VDD_M1007_b N_A_M1007_g 0.024954f $X=-0.045 $Y=2.645 $X2=0.475 $Y2=3.825
cc_60 N_VDD_c_60_p N_A_M1007_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475 $Y2=3.825
cc_61 N_VDD_c_61_p N_A_M1007_g 0.00362996f $X=0.69 $Y=3.885 $X2=0.475 $Y2=3.825
cc_62 N_VDD_c_62_p N_A_M1007_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.475 $Y2=3.825
cc_63 N_VDD_M1007_d N_A_c_108_n 0.00628533f $X=0.55 $Y=2.825 $X2=0.635 $Y2=2.22
cc_64 N_VDD_M1007_b N_A_c_108_n 0.00328912f $X=-0.045 $Y=2.645 $X2=0.635
+ $Y2=2.22
cc_65 N_VDD_c_61_p N_A_c_108_n 0.00264661f $X=0.69 $Y=3.885 $X2=0.635 $Y2=2.22
cc_66 N_VDD_M1007_d A 0.00797576f $X=0.55 $Y=2.825 $X2=0.635 $Y2=3.07
cc_67 N_VDD_c_61_p A 0.00510982f $X=0.69 $Y=3.885 $X2=0.635 $Y2=3.07
cc_68 N_VDD_M1007_b N_A_27_115#_c_174_n 0.01464f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=2.75
cc_69 N_VDD_c_61_p N_A_27_115#_c_174_n 0.00362996f $X=0.69 $Y=3.885 $X2=0.905
+ $Y2=2.75
cc_70 N_VDD_c_70_p N_A_27_115#_c_174_n 0.00496961f $X=1.465 $Y=5.397 $X2=0.905
+ $Y2=2.75
cc_71 N_VDD_c_62_p N_A_27_115#_c_174_n 0.00429146f $X=1.7 $Y=5.36 $X2=0.905
+ $Y2=2.75
cc_72 N_VDD_M1007_b N_A_27_115#_c_178_n 0.0144912f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.75
cc_73 N_VDD_c_61_p N_A_27_115#_c_178_n 3.67508e-19 $X=0.69 $Y=3.885 $X2=1.335
+ $Y2=2.75
cc_74 N_VDD_c_70_p N_A_27_115#_c_178_n 0.00500229f $X=1.465 $Y=5.397 $X2=1.335
+ $Y2=2.75
cc_75 N_VDD_c_75_p N_A_27_115#_c_178_n 0.00382402f $X=1.55 $Y=3.205 $X2=1.335
+ $Y2=2.75
cc_76 N_VDD_c_62_p N_A_27_115#_c_178_n 0.00430409f $X=1.7 $Y=5.36 $X2=1.335
+ $Y2=2.75
cc_77 N_VDD_M1007_b N_A_27_115#_c_152_n 0.00647677f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.675
cc_78 N_VDD_c_75_p N_A_27_115#_c_152_n 0.00364479f $X=1.55 $Y=3.205 $X2=1.69
+ $Y2=2.675
cc_79 N_VDD_M1007_b N_A_27_115#_c_153_n 0.0113915f $X=-0.045 $Y=2.645 $X2=1.41
+ $Y2=2.675
cc_80 N_VDD_M1007_b N_A_27_115#_c_186_n 0.0141812f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.75
cc_81 N_VDD_c_75_p N_A_27_115#_c_186_n 0.00362996f $X=1.55 $Y=3.205 $X2=1.765
+ $Y2=2.75
cc_82 N_VDD_c_82_p N_A_27_115#_c_186_n 0.00496961f $X=2.325 $Y=5.397 $X2=1.765
+ $Y2=2.75
cc_83 N_VDD_c_62_p N_A_27_115#_c_186_n 0.00429146f $X=1.7 $Y=5.36 $X2=1.765
+ $Y2=2.75
cc_84 N_VDD_M1007_b N_A_27_115#_c_159_n 0.0134369f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.675
cc_85 N_VDD_M1007_b N_A_27_115#_c_191_n 0.017048f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.75
cc_86 N_VDD_c_82_p N_A_27_115#_c_191_n 0.00496961f $X=2.325 $Y=5.397 $X2=2.195
+ $Y2=2.75
cc_87 N_VDD_c_87_p N_A_27_115#_c_191_n 0.00751602f $X=2.41 $Y=3.205 $X2=2.195
+ $Y2=2.75
cc_88 N_VDD_c_62_p N_A_27_115#_c_191_n 0.00429146f $X=1.7 $Y=5.36 $X2=2.195
+ $Y2=2.75
cc_89 N_VDD_M1007_b N_A_27_115#_c_165_n 0.00167153f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.675
cc_90 N_VDD_M1007_b N_A_27_115#_c_169_n 0.0103979f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.205
cc_91 N_VDD_c_60_p N_A_27_115#_c_169_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.205
cc_92 N_VDD_c_62_p N_A_27_115#_c_169_n 0.00435496f $X=1.7 $Y=5.36 $X2=0.26
+ $Y2=3.205
cc_93 N_VDD_M1007_b N_Y_c_280_n 0.00333732f $X=-0.045 $Y=2.645 $X2=1.12 $Y2=2.7
cc_94 N_VDD_c_70_p N_Y_c_280_n 0.0045126f $X=1.465 $Y=5.397 $X2=1.12 $Y2=2.7
cc_95 N_VDD_c_62_p N_Y_c_280_n 0.00434939f $X=1.7 $Y=5.36 $X2=1.12 $Y2=2.7
cc_96 N_VDD_M1007_b N_Y_c_283_n 0.00381442f $X=-0.045 $Y=2.645 $X2=1.98 $Y2=2.7
cc_97 N_VDD_c_82_p N_Y_c_283_n 0.00474282f $X=2.325 $Y=5.397 $X2=1.98 $Y2=2.7
cc_98 N_VDD_c_62_p N_Y_c_283_n 0.00434939f $X=1.7 $Y=5.36 $X2=1.98 $Y2=2.7
cc_99 N_VDD_M1007_b N_Y_c_271_n 0.00409378f $X=-0.045 $Y=2.645 $X2=1.12
+ $Y2=2.585
cc_100 N_VDD_M1007_b N_Y_c_287_n 0.00520877f $X=-0.045 $Y=2.645 $X2=1.835
+ $Y2=2.7
cc_101 N_VDD_c_75_p N_Y_c_287_n 0.0090257f $X=1.55 $Y=3.205 $X2=1.835 $Y2=2.7
cc_102 N_VDD_M1007_b N_Y_c_279_n 0.00409378f $X=-0.045 $Y=2.645 $X2=1.98
+ $Y2=2.585
cc_103 A N_A_27_115#_M1007_s 0.00414531f $X=0.635 $Y=3.07 $X2=0.135 $Y2=2.825
cc_104 N_A_M1006_g N_A_27_115#_M1002_g 0.0415224f $X=0.475 $Y=0.895 $X2=0.905
+ $Y2=0.895
cc_105 A N_A_27_115#_c_174_n 0.00419145f $X=0.635 $Y=3.07 $X2=0.905 $Y2=2.75
cc_106 N_A_M1006_g N_A_27_115#_c_145_n 0.00260138f $X=0.475 $Y=0.895 $X2=1.18
+ $Y2=2.6
cc_107 N_A_M1007_g N_A_27_115#_c_145_n 0.00209773f $X=0.475 $Y=3.825 $X2=1.18
+ $Y2=2.6
cc_108 N_A_c_107_n N_A_27_115#_c_145_n 0.0139096f $X=0.635 $Y=2.22 $X2=1.18
+ $Y2=2.6
cc_109 N_A_c_108_n N_A_27_115#_c_145_n 0.00361737f $X=0.635 $Y=2.22 $X2=1.18
+ $Y2=2.6
cc_110 N_A_M1007_g N_A_27_115#_c_153_n 0.0506363f $X=0.475 $Y=3.825 $X2=1.41
+ $Y2=2.675
cc_111 N_A_c_108_n N_A_27_115#_c_153_n 0.00477416f $X=0.635 $Y=2.22 $X2=1.41
+ $Y2=2.675
cc_112 N_A_M1006_g N_A_27_115#_c_166_n 0.0183389f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=0.865
cc_113 N_A_M1006_g N_A_27_115#_c_169_n 0.0341146f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=3.205
cc_114 N_A_c_108_n N_A_27_115#_c_169_n 0.0548951f $X=0.635 $Y=2.22 $X2=0.26
+ $Y2=3.205
cc_115 A N_A_27_115#_c_169_n 0.0155137f $X=0.635 $Y=3.07 $X2=0.26 $Y2=3.205
cc_116 N_A_M1006_g N_A_27_115#_c_170_n 0.0207696f $X=0.475 $Y=0.895 $X2=0.88
+ $Y2=1.675
cc_117 N_A_c_107_n N_A_27_115#_c_170_n 0.00273049f $X=0.635 $Y=2.22 $X2=0.88
+ $Y2=1.675
cc_118 N_A_c_108_n N_A_27_115#_c_170_n 0.00886797f $X=0.635 $Y=2.22 $X2=0.88
+ $Y2=1.675
cc_119 N_A_M1006_g N_A_27_115#_c_173_n 6.59135e-19 $X=0.475 $Y=0.895 $X2=0.965
+ $Y2=1.675
cc_120 N_A_c_108_n N_Y_c_280_n 0.0135622f $X=0.635 $Y=2.22 $X2=1.12 $Y2=2.7
cc_121 A N_Y_c_280_n 0.00731851f $X=0.635 $Y=3.07 $X2=1.12 $Y2=2.7
cc_122 N_A_M1006_g N_Y_c_268_n 8.23842e-19 $X=0.475 $Y=0.895 $X2=1.12 $Y2=1.335
cc_123 N_A_c_108_n N_Y_c_271_n 0.00677552f $X=0.635 $Y=2.22 $X2=1.12 $Y2=2.585
cc_124 N_A_M1006_g Y 0.00310306f $X=0.475 $Y=0.895 $X2=1.055 $Y2=2.01
cc_125 N_A_c_107_n Y 0.00441844f $X=0.635 $Y=2.22 $X2=1.055 $Y2=2.01
cc_126 N_A_c_108_n Y 0.0200396f $X=0.635 $Y=2.22 $X2=1.055 $Y2=2.01
cc_127 N_A_27_115#_M1002_g N_Y_c_260_n 0.00339663f $X=0.905 $Y=0.895 $X2=1.12
+ $Y2=0.865
cc_128 N_A_27_115#_M1003_g N_Y_c_260_n 0.00339663f $X=1.335 $Y=0.895 $X2=1.12
+ $Y2=0.865
cc_129 N_A_27_115#_c_151_n N_Y_c_260_n 0.0030245f $X=1.41 $Y=1.585 $X2=1.12
+ $Y2=0.865
cc_130 N_A_27_115#_c_173_n N_Y_c_260_n 7.50437e-19 $X=0.965 $Y=1.675 $X2=1.12
+ $Y2=0.865
cc_131 N_A_27_115#_c_174_n N_Y_c_280_n 0.00163525f $X=0.905 $Y=2.75 $X2=1.12
+ $Y2=2.7
cc_132 N_A_27_115#_c_178_n N_Y_c_280_n 0.00258898f $X=1.335 $Y=2.75 $X2=1.12
+ $Y2=2.7
cc_133 N_A_27_115#_c_153_n N_Y_c_280_n 0.0126676f $X=1.41 $Y=2.675 $X2=1.12
+ $Y2=2.7
cc_134 N_A_27_115#_M1008_g N_Y_c_264_n 0.00339663f $X=1.765 $Y=0.895 $X2=1.98
+ $Y2=0.865
cc_135 N_A_27_115#_c_158_n N_Y_c_264_n 0.00280419f $X=2.12 $Y=1.585 $X2=1.98
+ $Y2=0.865
cc_136 N_A_27_115#_M1009_g N_Y_c_264_n 0.00339663f $X=2.195 $Y=0.895 $X2=1.98
+ $Y2=0.865
cc_137 N_A_27_115#_c_186_n N_Y_c_283_n 0.00258898f $X=1.765 $Y=2.75 $X2=1.98
+ $Y2=2.7
cc_138 N_A_27_115#_c_159_n N_Y_c_283_n 0.013404f $X=2.12 $Y=2.675 $X2=1.98
+ $Y2=2.7
cc_139 N_A_27_115#_c_191_n N_Y_c_283_n 0.00258898f $X=2.195 $Y=2.75 $X2=1.98
+ $Y2=2.7
cc_140 N_A_27_115#_M1002_g N_Y_c_268_n 0.00541983f $X=0.905 $Y=0.895 $X2=1.12
+ $Y2=1.335
cc_141 N_A_27_115#_M1003_g N_Y_c_268_n 0.00259902f $X=1.335 $Y=0.895 $X2=1.12
+ $Y2=1.335
cc_142 N_A_27_115#_c_173_n N_Y_c_268_n 0.00278861f $X=0.965 $Y=1.675 $X2=1.12
+ $Y2=1.335
cc_143 N_A_27_115#_c_174_n N_Y_c_271_n 0.00120715f $X=0.905 $Y=2.75 $X2=1.12
+ $Y2=2.585
cc_144 N_A_27_115#_c_145_n N_Y_c_271_n 0.00215118f $X=1.18 $Y=2.6 $X2=1.12
+ $Y2=2.585
cc_145 N_A_27_115#_c_178_n N_Y_c_271_n 0.00113627f $X=1.335 $Y=2.75 $X2=1.12
+ $Y2=2.585
cc_146 N_A_27_115#_c_153_n N_Y_c_271_n 0.0038035f $X=1.41 $Y=2.675 $X2=1.12
+ $Y2=2.585
cc_147 N_A_27_115#_M1002_g Y 0.00251111f $X=0.905 $Y=0.895 $X2=1.055 $Y2=2.01
cc_148 N_A_27_115#_c_145_n Y 0.0314621f $X=1.18 $Y=2.6 $X2=1.055 $Y2=2.01
cc_149 N_A_27_115#_M1003_g Y 0.00251111f $X=1.335 $Y=0.895 $X2=1.055 $Y2=2.01
cc_150 N_A_27_115#_c_151_n Y 0.0166018f $X=1.41 $Y=1.585 $X2=1.055 $Y2=2.01
cc_151 N_A_27_115#_c_170_n Y 8.73078e-19 $X=0.88 $Y=1.675 $X2=1.055 $Y2=2.01
cc_152 N_A_27_115#_c_173_n Y 0.0121742f $X=0.965 $Y=1.675 $X2=1.055 $Y2=2.01
cc_153 N_A_27_115#_M1003_g N_Y_c_273_n 0.0130095f $X=1.335 $Y=0.895 $X2=1.835
+ $Y2=1.22
cc_154 N_A_27_115#_c_149_n N_Y_c_273_n 0.00213861f $X=1.69 $Y=1.585 $X2=1.835
+ $Y2=1.22
cc_155 N_A_27_115#_M1008_g N_Y_c_273_n 0.0130095f $X=1.765 $Y=0.895 $X2=1.835
+ $Y2=1.22
cc_156 N_A_27_115#_c_178_n N_Y_c_287_n 0.00639369f $X=1.335 $Y=2.75 $X2=1.835
+ $Y2=2.7
cc_157 N_A_27_115#_c_152_n N_Y_c_287_n 0.0125005f $X=1.69 $Y=2.675 $X2=1.835
+ $Y2=2.7
cc_158 N_A_27_115#_c_153_n N_Y_c_287_n 0.00580646f $X=1.41 $Y=2.675 $X2=1.835
+ $Y2=2.7
cc_159 N_A_27_115#_c_186_n N_Y_c_287_n 0.00639369f $X=1.765 $Y=2.75 $X2=1.835
+ $Y2=2.7
cc_160 N_A_27_115#_c_165_n N_Y_c_287_n 0.00580646f $X=1.765 $Y=2.675 $X2=1.835
+ $Y2=2.7
cc_161 N_A_27_115#_M1008_g N_Y_c_276_n 0.00259902f $X=1.765 $Y=0.895 $X2=1.98
+ $Y2=1.335
cc_162 N_A_27_115#_M1009_g N_Y_c_276_n 0.00939545f $X=2.195 $Y=0.895 $X2=1.98
+ $Y2=1.335
cc_163 N_A_27_115#_c_151_n N_Y_c_279_n 0.013329f $X=1.41 $Y=1.585 $X2=1.98
+ $Y2=2.585
cc_164 N_A_27_115#_M1008_g N_Y_c_279_n 0.00251111f $X=1.765 $Y=0.895 $X2=1.98
+ $Y2=2.585
cc_165 N_A_27_115#_c_186_n N_Y_c_279_n 0.00113627f $X=1.765 $Y=2.75 $X2=1.98
+ $Y2=2.585
cc_166 N_A_27_115#_c_158_n N_Y_c_279_n 0.0170354f $X=2.12 $Y=1.585 $X2=1.98
+ $Y2=2.585
cc_167 N_A_27_115#_c_159_n N_Y_c_279_n 0.00966211f $X=2.12 $Y=2.675 $X2=1.98
+ $Y2=2.585
cc_168 N_A_27_115#_M1009_g N_Y_c_279_n 0.00251111f $X=2.195 $Y=0.895 $X2=1.98
+ $Y2=2.585
cc_169 N_A_27_115#_c_191_n N_Y_c_279_n 0.0031083f $X=2.195 $Y=2.75 $X2=1.98
+ $Y2=2.585
cc_170 N_A_27_115#_c_165_n N_Y_c_279_n 6.99501e-19 $X=1.765 $Y=2.675 $X2=1.98
+ $Y2=2.585
