* File: sky130_osu_sc_15T_ls__nor2_1.pex.spice
* Created: Fri Nov 12 14:58:38 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__NOR2_1%GND 1 2 21 25 27 35 41 44
r27 41 44 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r28 33 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.865
r29 27 33 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.305
r30 23 25 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r31 21 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r32 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r33 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r34 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r35 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r36 2 35 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r37 1 25 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NOR2_1%VDD 1 13 15 21 29 32
r18 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r19 26 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r20 21 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.05 $Y=3.885
+ $X2=1.05 $Y2=4.565
r21 19 26 4.25596 $w=1.7e-07 $l=2.13185e-07 $layer=LI1_cond $X=1.05 $Y=5.245
+ $X2=1.197 $Y2=5.397
r22 19 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.05 $Y=5.245
+ $X2=1.05 $Y2=4.565
r23 15 26 3.30228 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=0.965 $Y=5.397
+ $X2=1.197 $Y2=5.397
r24 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=5.397
+ $X2=0.34 $Y2=5.397
r25 13 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r26 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r27 1 24 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.825 $X2=1.05 $Y2=4.565
r28 1 21 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.825 $X2=1.05 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NOR2_1%B 3 7 10 13 19 22
r49 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.65 $Y=2.7 $X2=0.65
+ $Y2=2.7
r50 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.65 $Y=1.915
+ $X2=0.65 $Y2=2.7
r51 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=1.83
+ $X2=0.65 $Y2=1.915
r52 13 15 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.565 $Y=1.83
+ $X2=0.415 $Y2=1.83
r53 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.83 $X2=0.415 $Y2=1.83
r54 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.83
+ $X2=0.415 $Y2=1.995
r55 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.83
+ $X2=0.415 $Y2=1.665
r56 7 12 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=1.995
r57 3 11 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=1.665
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NOR2_1%A 3 7 10 14 20
r36 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=3.07
+ $X2=0.99 $Y2=3.07
r37 14 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.99 $Y=2.495
+ $X2=0.99 $Y2=3.07
r38 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.495 $X2=0.99 $Y2=2.495
r39 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.495
+ $X2=0.942 $Y2=2.66
r40 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.495
+ $X2=0.942 $Y2=2.33
r41 7 11 710.181 $w=1.5e-07 $l=1.385e-06 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=2.33
r42 3 12 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=0.835 $Y=3.825
+ $X2=0.835 $Y2=2.66
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NOR2_1%Y 1 3 10 18 23 24 28 34
r41 26 28 0.519956 $w=1.7e-07 $l=5.4e-07 $layer=MET1_cond $X=0.69 $Y=2.245
+ $X2=0.69 $Y2=1.705
r42 25 34 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.22
r43 25 28 0.356266 $w=1.7e-07 $l=3.7e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.705
r44 24 31 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=2.33
+ $X2=0.26 $Y2=2.33
r45 23 26 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=2.33
+ $X2=0.69 $Y2=2.245
r46 23 24 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=2.33
+ $X2=0.405 $Y2=2.33
r47 21 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.22
+ $X2=0.69 $Y2=1.22
r48 18 21 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.69 $Y=0.865
+ $X2=0.69 $Y2=1.22
r49 13 15 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r50 10 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.33
+ $X2=0.26 $Y2=2.33
r51 10 13 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.26 $Y=2.33
+ $X2=0.26 $Y2=3.205
r52 3 15 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r53 3 13 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r54 1 18 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

