* File: sky130_osu_sc_18T_hs__addh_1.spice
* Created: Thu Oct 29 17:05:33 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_hs__addh_1.pex.spice"
.subckt sky130_osu_sc_18T_hs__addh_1  GND VDD CON B A S CO
* 
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1005 N_GND_M1005_d N_CON_M1005_g N_S_M1005_s N_GND_M1005_b NLOWVT L=0.15 W=1
+ AD=0.17 AS=0.265 PD=1.34 PS=2.53 NRD=7.188 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1008 A_208_115# N_B_M1008_g N_GND_M1005_d N_GND_M1005_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.17 PD=1.21 PS=1.34 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1009 N_A_208_617#_M1009_d N_A_M1009_g A_208_115# N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_GND_M1001_d N_A_208_617#_M1001_g N_CO_M1001_s N_GND_M1005_b NLOWVT
+ L=0.15 W=1 AD=0.17 AS=0.265 PD=1.34 PS=2.53 NRD=7.188 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1010 N_A_570_115#_M1010_d N_A_208_617#_M1010_g N_GND_M1001_d N_GND_M1005_b
+ NLOWVT L=0.15 W=1 AD=0.14 AS=0.17 PD=1.28 PS=1.34 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.7 SB=75001 A=0.15 P=2.3 MULT=1
MM1002 N_CON_M1002_d N_B_M1002_g N_A_570_115#_M1010_d N_GND_M1005_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.1 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_570_115#_M1003_d N_A_M1003_g N_CON_M1002_d N_GND_M1005_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_VDD_M1004_d N_CON_M1004_g N_S_M1004_s N_VDD_M1004_b PSHORT L=0.15 W=3
+ AD=0.51 AS=0.795 PD=3.34 PS=6.53 NRD=3.9203 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001.6 A=0.45 P=6.3 MULT=1
MM1006 N_A_208_617#_M1006_d N_B_M1006_g N_VDD_M1004_d N_VDD_M1004_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.51 PD=3.28 PS=3.34 NRD=0 NRS=0 M=1 R=20 SA=75000.7
+ SB=75001.1 A=0.45 P=6.3 MULT=1
MM1007 N_VDD_M1007_d N_A_M1007_g N_A_208_617#_M1006_d N_VDD_M1004_b PSHORT
+ L=0.15 W=3 AD=0.51 AS=0.42 PD=3.34 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.1
+ SB=75000.7 A=0.45 P=6.3 MULT=1
MM1013 N_CO_M1013_d N_A_208_617#_M1013_g N_VDD_M1007_d N_VDD_M1004_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.51 PD=6.53 PS=3.34 NRD=0 NRS=3.9203 M=1 R=20
+ SA=75001.6 SB=75000.2 A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_A_208_617#_M1000_g N_CON_M1000_s N_VDD_M1004_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1011 A_668_617# N_B_M1011_g N_VDD_M1000_d N_VDD_M1004_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1012 N_CON_M1012_d N_A_M1012_g A_668_617# N_VDD_M1004_b PSHORT L=0.15 W=3
+ AD=0.84 AS=0.315 PD=6.56 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX14_noxref N_GND_M1005_b N_VDD_M1004_b NWDIODE A=16.074 P=16.06
pX15_noxref noxref_12 S S PROBETYPE=1
pX16_noxref noxref_13 CO CO PROBETYPE=1
pX17_noxref noxref_14 B B PROBETYPE=1
pX18_noxref noxref_15 CON CON PROBETYPE=1
pX19_noxref noxref_16 A A PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__addh_1.pxi.spice"
*
.ends
*
*
