* File: sky130_osu_sc_15T_ls__and2_4.pxi.spice
* Created: Fri Nov 12 14:53:40 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__AND2_4%GND N_GND_M1003_d N_GND_M1007_s N_GND_M1010_s
+ N_GND_M1005_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p N_GND_c_22_p N_GND_c_30_p
+ N_GND_c_36_p GND N_GND_c_3_p PM_SKY130_OSU_SC_15T_LS__AND2_4%GND
x_PM_SKY130_OSU_SC_15T_LS__AND2_4%VDD N_VDD_M1000_s N_VDD_M1006_d N_VDD_M1004_s
+ N_VDD_M1011_s N_VDD_M1000_b N_VDD_c_75_p N_VDD_c_76_p N_VDD_c_87_p
+ N_VDD_c_94_p N_VDD_c_100_p N_VDD_c_106_p N_VDD_c_111_p VDD N_VDD_c_77_p
+ PM_SKY130_OSU_SC_15T_LS__AND2_4%VDD
x_PM_SKY130_OSU_SC_15T_LS__AND2_4%A N_A_M1005_g N_A_M1000_g N_A_c_130_n
+ N_A_c_131_n A PM_SKY130_OSU_SC_15T_LS__AND2_4%A
x_PM_SKY130_OSU_SC_15T_LS__AND2_4%B N_B_M1003_g N_B_M1006_g N_B_c_164_n
+ N_B_c_165_n B PM_SKY130_OSU_SC_15T_LS__AND2_4%B
x_PM_SKY130_OSU_SC_15T_LS__AND2_4%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1000_d N_A_27_115#_M1001_g N_A_27_115#_c_237_n
+ N_A_27_115#_M1002_g N_A_27_115#_c_204_n N_A_27_115#_c_205_n
+ N_A_27_115#_M1007_g N_A_27_115#_c_242_n N_A_27_115#_M1004_g
+ N_A_27_115#_c_210_n N_A_27_115#_c_212_n N_A_27_115#_c_213_n
+ N_A_27_115#_M1009_g N_A_27_115#_c_249_n N_A_27_115#_M1008_g
+ N_A_27_115#_c_218_n N_A_27_115#_c_219_n N_A_27_115#_M1010_g
+ N_A_27_115#_c_254_n N_A_27_115#_M1011_g N_A_27_115#_c_224_n
+ N_A_27_115#_c_225_n N_A_27_115#_c_226_n N_A_27_115#_c_227_n
+ N_A_27_115#_c_228_n N_A_27_115#_c_231_n N_A_27_115#_c_232_n
+ N_A_27_115#_c_261_n N_A_27_115#_c_233_n N_A_27_115#_c_235_n
+ N_A_27_115#_c_236_n N_A_27_115#_c_277_n
+ PM_SKY130_OSU_SC_15T_LS__AND2_4%A_27_115#
x_PM_SKY130_OSU_SC_15T_LS__AND2_4%Y N_Y_M1001_d N_Y_M1009_d N_Y_M1002_d
+ N_Y_M1008_d N_Y_c_335_n N_Y_c_340_n N_Y_c_341_n N_Y_c_345_n N_Y_c_346_n
+ N_Y_c_349_n Y N_Y_c_351_n N_Y_c_353_n N_Y_c_354_n N_Y_c_357_n
+ PM_SKY130_OSU_SC_15T_LS__AND2_4%Y
cc_1 N_GND_M1005_b N_A_M1005_g 0.0806078f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1005_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_A_M1005_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1005_b N_A_c_130_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.505
cc_5 N_GND_M1005_b N_A_c_131_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.505
cc_6 N_GND_M1005_b N_B_M1003_g 0.0460664f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_7 N_GND_c_2_p N_B_M1003_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.945
cc_8 N_GND_c_8_p N_B_M1003_g 0.00319969f $X=1.05 $Y=0.74 $X2=0.835 $Y2=0.945
cc_9 N_GND_c_3_p N_B_M1003_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.835 $Y2=0.945
cc_10 N_GND_M1005_b N_B_M1006_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_11 N_GND_M1005_b N_B_c_164_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.165
cc_12 N_GND_M1005_b N_B_c_165_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.165
cc_13 N_GND_M1005_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.7
cc_14 N_GND_M1005_b N_A_27_115#_M1001_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.945
cc_15 N_GND_c_8_p N_A_27_115#_M1001_g 0.00883341f $X=1.05 $Y=0.74 $X2=1.335
+ $Y2=0.945
cc_16 N_GND_c_16_p N_A_27_115#_M1001_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.945
cc_17 N_GND_c_3_p N_A_27_115#_M1001_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.335
+ $Y2=0.945
cc_18 N_GND_M1005_b N_A_27_115#_c_204_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.55
cc_19 N_GND_M1005_b N_A_27_115#_c_205_n 0.00954592f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.625
cc_20 N_GND_M1005_b N_A_27_115#_M1007_g 0.0202142f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.945
cc_21 N_GND_c_16_p N_A_27_115#_M1007_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.945
cc_22 N_GND_c_22_p N_A_27_115#_M1007_g 0.00327323f $X=1.98 $Y=0.74 $X2=1.765
+ $Y2=0.945
cc_23 N_GND_c_3_p N_A_27_115#_M1007_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.765
+ $Y2=0.945
cc_24 N_GND_M1005_b N_A_27_115#_c_210_n 0.0179436f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_25 N_GND_c_22_p N_A_27_115#_c_210_n 0.00291042f $X=1.98 $Y=0.74 $X2=2.12
+ $Y2=1.585
cc_26 N_GND_M1005_b N_A_27_115#_c_212_n 0.0448266f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.585
cc_27 N_GND_M1005_b N_A_27_115#_c_213_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.625
cc_28 N_GND_M1005_b N_A_27_115#_M1009_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.945
cc_29 N_GND_c_22_p N_A_27_115#_M1009_g 0.00327323f $X=1.98 $Y=0.74 $X2=2.195
+ $Y2=0.945
cc_30 N_GND_c_30_p N_A_27_115#_M1009_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.945
cc_31 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.195
+ $Y2=0.945
cc_32 N_GND_M1005_b N_A_27_115#_c_218_n 0.0369419f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.585
cc_33 N_GND_M1005_b N_A_27_115#_c_219_n 0.0268552f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.625
cc_34 N_GND_M1005_b N_A_27_115#_M1010_g 0.0264941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.945
cc_35 N_GND_c_30_p N_A_27_115#_M1010_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.945
cc_36 N_GND_c_36_p N_A_27_115#_M1010_g 0.00502587f $X=2.84 $Y=0.74 $X2=2.625
+ $Y2=0.945
cc_37 N_GND_c_3_p N_A_27_115#_M1010_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.625
+ $Y2=0.945
cc_38 N_GND_M1005_b N_A_27_115#_c_224_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.625
cc_39 N_GND_M1005_b N_A_27_115#_c_225_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.625
cc_40 N_GND_M1005_b N_A_27_115#_c_226_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.585
cc_41 N_GND_M1005_b N_A_27_115#_c_227_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.625
cc_42 N_GND_M1005_b N_A_27_115#_c_228_n 0.0143389f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_43 N_GND_c_2_p N_A_27_115#_c_228_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_44 N_GND_c_3_p N_A_27_115#_c_228_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_45 N_GND_M1005_b N_A_27_115#_c_231_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.675
cc_46 N_GND_M1005_b N_A_27_115#_c_232_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.675
cc_47 N_GND_M1005_b N_A_27_115#_c_233_n 0.0227928f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_48 N_GND_c_8_p N_A_27_115#_c_233_n 0.00833003f $X=1.05 $Y=0.74 $X2=1.43
+ $Y2=1.675
cc_49 N_GND_M1005_b N_A_27_115#_c_235_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.675
cc_50 N_GND_M1005_b N_A_27_115#_c_236_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.305
cc_51 N_GND_M1005_b N_Y_c_335_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.74
cc_52 N_GND_c_8_p N_Y_c_335_n 0.0150458f $X=1.05 $Y=0.74 $X2=1.55 $Y2=0.74
cc_53 N_GND_c_16_p N_Y_c_335_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.74
cc_54 N_GND_c_22_p N_Y_c_335_n 0.0029082f $X=1.98 $Y=0.74 $X2=1.55 $Y2=0.74
cc_55 N_GND_c_3_p N_Y_c_335_n 0.00475776f $X=2.38 $Y=0.19 $X2=1.55 $Y2=0.74
cc_56 N_GND_M1005_b N_Y_c_340_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_57 N_GND_M1005_b N_Y_c_341_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.74
cc_58 N_GND_c_22_p N_Y_c_341_n 0.0029082f $X=1.98 $Y=0.74 $X2=2.41 $Y2=0.74
cc_59 N_GND_c_30_p N_Y_c_341_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.74
cc_60 N_GND_c_3_p N_Y_c_341_n 0.00475776f $X=2.38 $Y=0.19 $X2=2.41 $Y2=0.74
cc_61 N_GND_M1005_b N_Y_c_345_n 0.0152877f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.33
cc_62 N_GND_M1005_b N_Y_c_346_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.335
cc_63 N_GND_c_8_p N_Y_c_346_n 0.00377613f $X=1.05 $Y=0.74 $X2=1.55 $Y2=1.335
cc_64 N_GND_c_22_p N_Y_c_346_n 7.53951e-19 $X=1.98 $Y=0.74 $X2=1.55 $Y2=1.335
cc_65 N_GND_M1005_b N_Y_c_349_n 0.00463624f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.215
cc_66 N_GND_M1005_b Y 0.0306813f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.96
cc_67 N_GND_M1007_s N_Y_c_351_n 0.0127109f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.22
cc_68 N_GND_c_22_p N_Y_c_351_n 0.0175563f $X=1.98 $Y=0.74 $X2=2.265 $Y2=1.22
cc_69 N_GND_M1005_b N_Y_c_353_n 0.0188475f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.33
cc_70 N_GND_M1005_b N_Y_c_354_n 0.00409378f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.335
cc_71 N_GND_c_22_p N_Y_c_354_n 7.53951e-19 $X=1.98 $Y=0.74 $X2=2.41 $Y2=1.335
cc_72 N_GND_c_36_p N_Y_c_354_n 0.00399019f $X=2.84 $Y=0.74 $X2=2.41 $Y2=1.335
cc_73 N_GND_M1005_b N_Y_c_357_n 0.06145f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.215
cc_74 N_VDD_M1000_b N_A_M1000_g 0.0193382f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_75 N_VDD_c_75_p N_A_M1000_g 0.00713292f $X=0.26 $Y=3.895 $X2=0.475 $Y2=3.825
cc_76 N_VDD_c_76_p N_A_M1000_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475 $Y2=3.825
cc_77 N_VDD_c_77_p N_A_M1000_g 0.00429146f $X=2.38 $Y=5.36 $X2=0.475 $Y2=3.825
cc_78 N_VDD_M1000_b N_A_c_130_n 0.0111025f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=2.505
cc_79 N_VDD_M1000_s N_A_c_131_n 0.0127742f $X=0.135 $Y=2.825 $X2=0.27 $Y2=2.505
cc_80 N_VDD_M1000_b N_A_c_131_n 0.00612103f $X=-0.045 $Y=2.645 $X2=0.27
+ $Y2=2.505
cc_81 N_VDD_c_75_p N_A_c_131_n 0.00352433f $X=0.26 $Y=3.895 $X2=0.27 $Y2=2.505
cc_82 N_VDD_M1000_s A 0.00746694f $X=0.135 $Y=2.825 $X2=0.275 $Y2=3.07
cc_83 N_VDD_M1000_b A 0.00970321f $X=-0.045 $Y=2.645 $X2=0.275 $Y2=3.07
cc_84 N_VDD_c_75_p A 0.00428937f $X=0.26 $Y=3.895 $X2=0.275 $Y2=3.07
cc_85 N_VDD_M1000_b N_B_M1006_g 0.0191387f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_86 N_VDD_c_76_p N_B_M1006_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905 $Y2=3.825
cc_87 N_VDD_c_87_p N_B_M1006_g 0.00354579f $X=1.12 $Y=3.555 $X2=0.905 $Y2=3.825
cc_88 N_VDD_c_77_p N_B_M1006_g 0.00429146f $X=2.38 $Y=5.36 $X2=0.905 $Y2=3.825
cc_89 N_VDD_M1000_b N_B_c_165_n 0.00170274f $X=-0.045 $Y=2.645 $X2=0.95
+ $Y2=2.165
cc_90 N_VDD_M1000_b B 0.00860092f $X=-0.045 $Y=2.645 $X2=0.955 $Y2=2.7
cc_91 N_VDD_c_87_p B 0.00236322f $X=1.12 $Y=3.555 $X2=0.955 $Y2=2.7
cc_92 N_VDD_M1000_b N_A_27_115#_c_237_n 0.0174951f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.7
cc_93 N_VDD_c_87_p N_A_27_115#_c_237_n 0.00354579f $X=1.12 $Y=3.555 $X2=1.335
+ $Y2=2.7
cc_94 N_VDD_c_94_p N_A_27_115#_c_237_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335
+ $Y2=2.7
cc_95 N_VDD_c_77_p N_A_27_115#_c_237_n 0.00429146f $X=2.38 $Y=5.36 $X2=1.335
+ $Y2=2.7
cc_96 N_VDD_M1000_b N_A_27_115#_c_205_n 0.00428234f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_97 N_VDD_M1000_b N_A_27_115#_c_242_n 0.0173909f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.7
cc_98 N_VDD_c_87_p N_A_27_115#_c_242_n 3.67508e-19 $X=1.12 $Y=3.555 $X2=1.765
+ $Y2=2.7
cc_99 N_VDD_c_94_p N_A_27_115#_c_242_n 0.00500229f $X=1.895 $Y=5.397 $X2=1.765
+ $Y2=2.7
cc_100 N_VDD_c_100_p N_A_27_115#_c_242_n 0.00373985f $X=1.98 $Y=3.215 $X2=1.765
+ $Y2=2.7
cc_101 N_VDD_c_77_p N_A_27_115#_c_242_n 0.00430409f $X=2.38 $Y=5.36 $X2=1.765
+ $Y2=2.7
cc_102 N_VDD_M1000_b N_A_27_115#_c_213_n 0.00399373f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.625
cc_103 N_VDD_c_100_p N_A_27_115#_c_213_n 0.0037128f $X=1.98 $Y=3.215 $X2=2.12
+ $Y2=2.625
cc_104 N_VDD_M1000_b N_A_27_115#_c_249_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.7
cc_105 N_VDD_c_100_p N_A_27_115#_c_249_n 0.00354579f $X=1.98 $Y=3.215 $X2=2.195
+ $Y2=2.7
cc_106 N_VDD_c_106_p N_A_27_115#_c_249_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.195
+ $Y2=2.7
cc_107 N_VDD_c_77_p N_A_27_115#_c_249_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.195
+ $Y2=2.7
cc_108 N_VDD_M1000_b N_A_27_115#_c_219_n 0.00840215f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.625
cc_109 N_VDD_M1000_b N_A_27_115#_c_254_n 0.0212947f $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.7
cc_110 N_VDD_c_106_p N_A_27_115#_c_254_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.625
+ $Y2=2.7
cc_111 N_VDD_c_111_p N_A_27_115#_c_254_n 0.00713292f $X=2.84 $Y=3.215 $X2=2.625
+ $Y2=2.7
cc_112 N_VDD_c_77_p N_A_27_115#_c_254_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.625
+ $Y2=2.7
cc_113 N_VDD_M1000_b N_A_27_115#_c_224_n 0.0021704f $X=-0.045 $Y=2.645 $X2=1.352
+ $Y2=2.625
cc_114 N_VDD_M1000_b N_A_27_115#_c_225_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=1.765 $Y2=2.625
cc_115 N_VDD_M1000_b N_A_27_115#_c_227_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.195 $Y2=2.625
cc_116 N_VDD_M1000_b N_A_27_115#_c_261_n 0.00198641f $X=-0.045 $Y=2.645 $X2=0.69
+ $Y2=3.555
cc_117 N_VDD_c_76_p N_A_27_115#_c_261_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69
+ $Y2=3.555
cc_118 N_VDD_c_77_p N_A_27_115#_c_261_n 0.00434939f $X=2.38 $Y=5.36 $X2=0.69
+ $Y2=3.555
cc_119 N_VDD_M1000_b N_A_27_115#_c_236_n 8.22047e-19 $X=-0.045 $Y=2.645 $X2=0.65
+ $Y2=3.305
cc_120 N_VDD_M1000_b N_Y_c_340_n 0.00388477f $X=-0.045 $Y=2.645 $X2=1.55
+ $Y2=2.33
cc_121 N_VDD_c_94_p N_Y_c_340_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.33
cc_122 N_VDD_c_77_p N_Y_c_340_n 0.00434939f $X=2.38 $Y=5.36 $X2=1.55 $Y2=2.33
cc_123 N_VDD_M1000_b N_Y_c_345_n 0.0042387f $X=-0.045 $Y=2.645 $X2=2.41 $Y2=2.33
cc_124 N_VDD_c_106_p N_Y_c_345_n 0.0045126f $X=2.755 $Y=5.397 $X2=2.41 $Y2=2.33
cc_125 N_VDD_c_77_p N_Y_c_345_n 0.00434939f $X=2.38 $Y=5.36 $X2=2.41 $Y2=2.33
cc_126 N_VDD_c_100_p N_Y_c_353_n 0.00622932f $X=1.98 $Y=3.215 $X2=2.265 $Y2=2.33
cc_127 N_A_M1005_g N_B_M1003_g 0.113664f $X=0.475 $Y=0.945 $X2=0.835 $Y2=0.945
cc_128 N_A_M1005_g N_B_M1006_g 0.0506107f $X=0.475 $Y=0.945 $X2=0.905 $Y2=3.825
cc_129 N_A_M1005_g N_B_c_165_n 7.8234e-19 $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.165
cc_130 N_A_M1005_g N_A_27_115#_c_228_n 0.0114001f $X=0.475 $Y=0.945 $X2=0.26
+ $Y2=0.74
cc_131 N_A_M1005_g N_A_27_115#_c_231_n 0.0160984f $X=0.475 $Y=0.945 $X2=0.525
+ $Y2=1.675
cc_132 N_A_c_130_n N_A_27_115#_c_231_n 0.00117122f $X=0.475 $Y=2.505 $X2=0.525
+ $Y2=1.675
cc_133 N_A_c_131_n N_A_27_115#_c_231_n 2.65873e-19 $X=0.27 $Y=2.505 $X2=0.525
+ $Y2=1.675
cc_134 N_A_c_130_n N_A_27_115#_c_232_n 0.00133457f $X=0.475 $Y=2.505 $X2=0.345
+ $Y2=1.675
cc_135 N_A_c_131_n N_A_27_115#_c_232_n 0.0055861f $X=0.27 $Y=2.505 $X2=0.345
+ $Y2=1.675
cc_136 N_A_M1005_g N_A_27_115#_c_235_n 0.00322084f $X=0.475 $Y=0.945 $X2=0.61
+ $Y2=1.675
cc_137 N_A_M1005_g N_A_27_115#_c_236_n 0.0265302f $X=0.475 $Y=0.945 $X2=0.65
+ $Y2=3.305
cc_138 N_A_M1000_g N_A_27_115#_c_236_n 0.0149699f $X=0.475 $Y=3.825 $X2=0.65
+ $Y2=3.305
cc_139 N_A_c_130_n N_A_27_115#_c_236_n 0.00766302f $X=0.475 $Y=2.505 $X2=0.65
+ $Y2=3.305
cc_140 N_A_c_131_n N_A_27_115#_c_236_n 0.0456533f $X=0.27 $Y=2.505 $X2=0.65
+ $Y2=3.305
cc_141 A N_A_27_115#_c_236_n 0.00758489f $X=0.275 $Y=3.07 $X2=0.65 $Y2=3.305
cc_142 N_A_M1000_g N_A_27_115#_c_277_n 0.00884152f $X=0.475 $Y=3.825 $X2=0.65
+ $Y2=3.475
cc_143 N_B_M1003_g N_A_27_115#_M1001_g 0.0276217f $X=0.835 $Y=0.945 $X2=1.335
+ $Y2=0.945
cc_144 N_B_M1006_g N_A_27_115#_c_204_n 0.00773101f $X=0.905 $Y=3.825 $X2=1.37
+ $Y2=2.55
cc_145 N_B_c_164_n N_A_27_115#_c_204_n 0.0206104f $X=0.95 $Y=2.165 $X2=1.37
+ $Y2=2.55
cc_146 N_B_c_165_n N_A_27_115#_c_204_n 0.0033451f $X=0.95 $Y=2.165 $X2=1.37
+ $Y2=2.55
cc_147 N_B_M1003_g N_A_27_115#_c_212_n 0.0104742f $X=0.835 $Y=0.945 $X2=1.84
+ $Y2=1.585
cc_148 N_B_M1006_g N_A_27_115#_c_224_n 0.0410292f $X=0.905 $Y=3.825 $X2=1.352
+ $Y2=2.625
cc_149 N_B_c_165_n N_A_27_115#_c_224_n 0.00173699f $X=0.95 $Y=2.165 $X2=1.352
+ $Y2=2.625
cc_150 B N_A_27_115#_c_224_n 0.00389258f $X=0.955 $Y=2.7 $X2=1.352 $Y2=2.625
cc_151 N_B_M1003_g N_A_27_115#_c_233_n 0.0182215f $X=0.835 $Y=0.945 $X2=1.43
+ $Y2=1.675
cc_152 N_B_c_164_n N_A_27_115#_c_233_n 0.00258465f $X=0.95 $Y=2.165 $X2=1.43
+ $Y2=1.675
cc_153 N_B_c_165_n N_A_27_115#_c_233_n 0.0101796f $X=0.95 $Y=2.165 $X2=1.43
+ $Y2=1.675
cc_154 N_B_M1003_g N_A_27_115#_c_236_n 0.00755919f $X=0.835 $Y=0.945 $X2=0.65
+ $Y2=3.305
cc_155 N_B_M1006_g N_A_27_115#_c_236_n 0.0137515f $X=0.905 $Y=3.825 $X2=0.65
+ $Y2=3.305
cc_156 N_B_c_165_n N_A_27_115#_c_236_n 0.0541375f $X=0.95 $Y=2.165 $X2=0.65
+ $Y2=3.305
cc_157 B N_A_27_115#_c_236_n 0.00866797f $X=0.955 $Y=2.7 $X2=0.65 $Y2=3.305
cc_158 B N_A_27_115#_c_277_n 0.00281588f $X=0.955 $Y=2.7 $X2=0.65 $Y2=3.475
cc_159 N_B_c_165_n N_Y_c_340_n 0.0149875f $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.33
cc_160 B N_Y_c_340_n 0.00649253f $X=0.955 $Y=2.7 $X2=1.55 $Y2=2.33
cc_161 N_B_M1003_g N_Y_c_346_n 3.57178e-19 $X=0.835 $Y=0.945 $X2=1.55 $Y2=1.335
cc_162 N_B_c_164_n N_Y_c_349_n 5.85867e-19 $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.215
cc_163 N_B_c_165_n N_Y_c_349_n 0.00592261f $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.215
cc_164 N_B_M1003_g Y 6.71108e-19 $X=0.835 $Y=0.945 $X2=1.555 $Y2=1.96
cc_165 N_B_c_165_n Y 0.00695761f $X=0.95 $Y=2.165 $X2=1.555 $Y2=1.96
cc_166 N_A_27_115#_M1001_g N_Y_c_335_n 9.07985e-19 $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=0.74
cc_167 N_A_27_115#_M1007_g N_Y_c_335_n 8.52215e-19 $X=1.765 $Y=0.945 $X2=1.55
+ $Y2=0.74
cc_168 N_A_27_115#_c_212_n N_Y_c_335_n 0.00171364f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=0.74
cc_169 N_A_27_115#_c_233_n N_Y_c_335_n 0.00500271f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.74
cc_170 N_A_27_115#_c_237_n N_Y_c_340_n 0.00287202f $X=1.335 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_171 N_A_27_115#_c_204_n N_Y_c_340_n 0.00744772f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_172 N_A_27_115#_c_205_n N_Y_c_340_n 0.0167599f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_173 N_A_27_115#_c_242_n N_Y_c_340_n 0.00401146f $X=1.765 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_174 N_A_27_115#_c_212_n N_Y_c_340_n 0.0013767f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.33
cc_175 N_A_27_115#_c_233_n N_Y_c_340_n 0.00273485f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_176 N_A_27_115#_M1009_g N_Y_c_341_n 8.52215e-19 $X=2.195 $Y=0.945 $X2=2.41
+ $Y2=0.74
cc_177 N_A_27_115#_c_218_n N_Y_c_341_n 0.00280419f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=0.74
cc_178 N_A_27_115#_M1010_g N_Y_c_341_n 8.52215e-19 $X=2.625 $Y=0.945 $X2=2.41
+ $Y2=0.74
cc_179 N_A_27_115#_c_249_n N_Y_c_345_n 0.00401146f $X=2.195 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_180 N_A_27_115#_c_218_n N_Y_c_345_n 0.00250559f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.33
cc_181 N_A_27_115#_c_219_n N_Y_c_345_n 0.0206674f $X=2.55 $Y=2.625 $X2=2.41
+ $Y2=2.33
cc_182 N_A_27_115#_c_254_n N_Y_c_345_n 0.00401146f $X=2.625 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_183 N_A_27_115#_M1001_g N_Y_c_346_n 0.00345902f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=1.335
cc_184 N_A_27_115#_M1007_g N_Y_c_346_n 0.00134358f $X=1.765 $Y=0.945 $X2=1.55
+ $Y2=1.335
cc_185 N_A_27_115#_c_233_n N_Y_c_346_n 0.00238892f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=1.335
cc_186 N_A_27_115#_c_204_n N_Y_c_349_n 0.00821104f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.215
cc_187 N_A_27_115#_c_205_n N_Y_c_349_n 0.00229755f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.215
cc_188 N_A_27_115#_c_212_n N_Y_c_349_n 0.00174847f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.215
cc_189 N_A_27_115#_c_233_n N_Y_c_349_n 0.00181779f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.215
cc_190 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=0.945 $X2=1.555 $Y2=1.96
cc_191 N_A_27_115#_c_204_n Y 0.00892438f $X=1.37 $Y=2.55 $X2=1.555 $Y2=1.96
cc_192 N_A_27_115#_M1007_g Y 0.00251111f $X=1.765 $Y=0.945 $X2=1.555 $Y2=1.96
cc_193 N_A_27_115#_c_212_n Y 0.0128645f $X=1.84 $Y=1.585 $X2=1.555 $Y2=1.96
cc_194 N_A_27_115#_c_233_n Y 0.0148238f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_195 N_A_27_115#_M1007_g N_Y_c_351_n 0.0120124f $X=1.765 $Y=0.945 $X2=2.265
+ $Y2=1.22
cc_196 N_A_27_115#_c_210_n N_Y_c_351_n 0.00213861f $X=2.12 $Y=1.585 $X2=2.265
+ $Y2=1.22
cc_197 N_A_27_115#_M1009_g N_Y_c_351_n 0.0120124f $X=2.195 $Y=0.945 $X2=2.265
+ $Y2=1.22
cc_198 N_A_27_115#_c_212_n N_Y_c_353_n 0.0121767f $X=1.84 $Y=1.585 $X2=2.265
+ $Y2=2.33
cc_199 N_A_27_115#_c_225_n N_Y_c_353_n 0.0158479f $X=1.765 $Y=2.625 $X2=2.265
+ $Y2=2.33
cc_200 N_A_27_115#_M1009_g N_Y_c_354_n 0.00134358f $X=2.195 $Y=0.945 $X2=2.41
+ $Y2=1.335
cc_201 N_A_27_115#_M1010_g N_Y_c_354_n 0.00534683f $X=2.625 $Y=0.945 $X2=2.41
+ $Y2=1.335
cc_202 N_A_27_115#_M1009_g N_Y_c_357_n 0.00251111f $X=2.195 $Y=0.945 $X2=2.41
+ $Y2=2.215
cc_203 N_A_27_115#_c_218_n N_Y_c_357_n 0.0184054f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_204 N_A_27_115#_M1010_g N_Y_c_357_n 0.00251111f $X=2.625 $Y=0.945 $X2=2.41
+ $Y2=2.215
cc_205 N_A_27_115#_c_226_n N_Y_c_357_n 0.00140336f $X=2.195 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_206 N_A_27_115#_c_227_n N_Y_c_357_n 0.00372651f $X=2.195 $Y=2.625 $X2=2.41
+ $Y2=2.215
