* File: sky130_osu_sc_18T_ls__addh_l.pex.spice
* Created: Thu Oct 29 17:33:30 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%GND 1 2 31 35 37 50 52 60 62
r96 60 62 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r97 54 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r98 52 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r99 48 55 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r100 48 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.825
r101 38 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r102 37 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r103 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r104 33 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.825
r105 31 54 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r106 31 52 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r107 31 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.17
+ $X2=3.74 $Y2=0.17
r108 31 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r109 31 37 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r110 31 38 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r111 2 50 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.825
r112 1 35 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%VDD 1 2 3 28 32 36 42 46 54 58 65 70 77
r58 70 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=6.49
+ $X2=3.74 $Y2=6.49
r59 65 70 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.74 $Y2=6.507
r60 65 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r61 61 77 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.74 $Y2=6.507
r62 61 63 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.05 $Y2=6.507
r63 58 74 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.34 $Y2=6.507
r64 58 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.75 $Y2=6.507
r65 54 57 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.05 $Y=3.455
+ $X2=3.05 $Y2=5.835
r66 52 63 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=6.507
r67 52 57 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=5.835
r68 49 51 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=6.507
+ $X2=2.38 $Y2=6.507
r69 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.61 $Y2=6.507
r70 47 49 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.7 $Y2=6.507
r71 46 63 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=3.05 $Y2=6.507
r72 46 51 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=2.38 $Y2=6.507
r73 42 45 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.61 $Y=3.795
+ $X2=1.61 $Y2=5.835
r74 40 60 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=6.507
r75 40 45 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=5.835
r76 37 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=0.75 $Y2=6.507
r77 37 39 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=1.02 $Y2=6.507
r78 36 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.61 $Y2=6.507
r79 36 39 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.02 $Y2=6.507
r80 32 35 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.75 $Y=3.455
+ $X2=0.75 $Y2=5.835
r81 30 59 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=6.507
r82 30 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=5.835
r83 28 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r84 28 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r85 28 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r86 28 51 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r87 28 49 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r88 28 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r89 3 57 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=5.835
r90 3 54 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=3.455
r91 2 45 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=5.835
r92 2 42 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=3.795
r93 1 35 150 $w=1.7e-07 $l=1.49666e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=4.435 $X2=0.75 $Y2=5.835
r94 1 32 150 $w=1.7e-07 $l=1.07536e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=4.435 $X2=0.75 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%CON 1 2 3 12 16 18 19 22 26 28 30 32 36
+ 40 41 42 45 48 52 58
c128 52 0 2.7119e-19 $X=3.42 $Y=1.85
c129 42 0 1.57622e-19 $X=0.78 $Y=1.85
c130 30 0 1.92558e-19 $X=3.42 $Y=1.765
r131 58 60 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=2.015
r132 58 59 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=1.685
r133 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.85 $X2=0.35 $Y2=1.85
r134 52 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.85
+ $X2=3.42 $Y2=1.85
r135 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.85
+ $X2=2.62 $Y2=1.85
r136 45 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.635 $Y=1.85
+ $X2=0.35 $Y2=1.85
r137 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.85
+ $X2=0.635 $Y2=1.85
r138 42 44 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.85
+ $X2=0.635 $Y2=1.85
r139 41 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=2.62 $Y2=1.85
r140 41 42 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=0.78 $Y2=1.85
r141 36 38 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.84 $Y=3.455
+ $X2=3.84 $Y2=5.835
r142 34 36 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.84 $Y=3.035
+ $X2=3.84 $Y2=3.455
r143 30 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.85
r144 30 32 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.165
r145 29 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.95
+ $X2=2.62 $Y2=2.95
r146 28 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=3.84 $Y2=3.035
r147 28 29 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=2.705 $Y2=2.95
r148 27 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.85
+ $X2=2.62 $Y2=1.85
r149 26 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=3.42 $Y2=1.85
r150 26 27 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=2.705 $Y2=1.85
r151 22 24 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.62 $Y=3.455
+ $X2=2.62 $Y2=5.835
r152 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=2.95
r153 20 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=3.455
r154 19 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.865
+ $X2=2.62 $Y2=2.95
r155 18 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=1.85
r156 18 19 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=2.865
r157 16 60 1663.93 $w=1.5e-07 $l=3.245e-06 $layer=POLY_cond $X=0.475 $Y=5.26
+ $X2=0.475 $Y2=2.015
r158 12 59 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=1.685
r159 3 38 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=5.835
r160 3 36 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=3.455
r161 2 24 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=5.835
r162 2 22 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=3.455
r163 1 32 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=1.165
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%B 3 7 11 15 21 23 26 27 28 33 38
c101 38 0 1.42567e-19 $X=3.205 $Y=2.22
c102 33 0 1.57622e-19 $X=0.905 $Y=2.22
c103 28 0 4.99902e-20 $X=3.21 $Y=2.22
r104 38 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.385
r105 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.385
r106 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.055
r107 27 28 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.06 $Y=2.22
+ $X2=3.205 $Y2=2.22
r108 26 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=2.22 $X2=3.205 $Y2=2.22
r109 26 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.22
r110 23 27 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=2.222
+ $X2=3.06 $Y2=2.222
r111 21 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=2.22 $X2=0.905 $Y2=2.22
r112 20 23 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=2.22
+ $X2=1.05 $Y2=2.22
r113 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.22
r114 15 39 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=3.265 $Y=4.585
+ $X2=3.265 $Y2=2.385
r115 9 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=2.22
r116 9 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=1.075
r117 7 35 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.965 $Y=4.585
+ $X2=0.965 $Y2=2.385
r118 3 34 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.965 $Y=1.075
+ $X2=0.965 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%A 3 7 11 15 21 23 25 26 28 33 38
c87 38 0 1.74252e-19 $X=3.685 $Y=2.59
r88 38 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.755
r89 38 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.425
r90 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.755
r91 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.425
r92 28 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.59 $X2=3.685 $Y2=2.59
r93 25 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.59
r94 25 26 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.59
+ $X2=3.54 $Y2=2.59
r95 23 26 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.587
+ $X2=3.54 $Y2=2.587
r96 21 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.59 $X2=1.385 $Y2=2.59
r97 20 23 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.59
+ $X2=1.53 $Y2=2.59
r98 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.59
r99 15 39 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=3.635 $Y=1.075
+ $X2=3.635 $Y2=2.425
r100 11 40 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.625 $Y=4.585
+ $X2=3.625 $Y2=2.755
r101 7 35 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=1.395 $Y=4.585
+ $X2=1.395 $Y2=2.755
r102 3 34 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=1.325 $Y=1.075
+ $X2=1.325 $Y2=2.425
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%A_208_617# 1 2 8 11 13 15 19 21 25 29 31
+ 32 35 39 40 43 46 48 52
c114 29 0 2.52869e-20 $X=2.835 $Y=4.585
c115 21 0 9.69384e-20 $X=2.7 $Y=1.8
r116 51 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.955
+ $X2=1.825 $Y2=2.12
r117 51 52 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.955
+ $X2=1.825 $Y2=1.8
r118 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.955 $X2=1.825 $Y2=1.955
r119 48 50 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.955
+ $X2=1.825 $Y2=1.955
r120 47 48 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.955
+ $X2=1.725 $Y2=1.955
r121 45 48 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=1.955
r122 45 46 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=2.925
r123 41 47 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=1.955
r124 41 43 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=0.825
r125 39 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.725 $Y2=2.925
r126 39 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.265 $Y2=3.01
r127 35 37 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.18 $Y=3.795
+ $X2=1.18 $Y2=5.835
r128 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.265 $Y2=3.01
r129 33 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.18 $Y2=3.795
r130 27 29 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=2.835 $Y=2.745
+ $X2=2.835 $Y2=4.585
r131 23 25 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=1.075
r132 22 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.8
+ $X2=2.285 $Y2=1.8
r133 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.8
+ $X2=2.775 $Y2=1.725
r134 21 22 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.8 $X2=2.36
+ $Y2=1.8
r135 17 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=1.8
r136 17 19 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=0.895
r137 16 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.67
+ $X2=1.885 $Y2=2.67
r138 15 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.67
+ $X2=2.835 $Y2=2.745
r139 15 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.67 $X2=1.96
+ $Y2=2.67
r140 14 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.8
+ $X2=1.825 $Y2=1.8
r141 13 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=2.285 $Y2=1.8
r142 13 14 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=1.96 $Y2=1.8
r143 9 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=2.67
r144 9 11 1289.61 $w=1.5e-07 $l=2.515e-06 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=5.26
r145 8 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.67
r146 8 55 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.12
r147 2 37 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=5.835
r148 2 35 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=3.795
r149 1 43 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%S 1 2 10 13 17 18 21
r32 28 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=4.815
+ $X2=0.26 $Y2=5.835
r33 18 28 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=4.815
r34 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=3.33
r35 14 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.26 $Y=1.475
+ $X2=0.26 $Y2=0.825
r36 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.475
+ $X2=0.26 $Y2=1.475
r37 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=3.33
r38 8 10 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=2.385
r39 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=1.475
r40 7 10 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=2.385
r41 2 30 300 $w=1.7e-07 $l=1.46116e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.435 $X2=0.26 $Y2=5.835
r42 2 28 300 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.435 $X2=0.26 $Y2=4.815
r43 1 21 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%CO 1 2 9 13 21 24 26 29
c55 26 0 2.52869e-20 $X=2.175 $Y=2.96
r56 26 30 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=3.045
r57 26 29 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=2.875
r58 24 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.96
+ $X2=2.175 $Y2=2.96
r59 17 21 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=1.472
r60 17 29 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=2.875
r61 13 15 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.1 $Y=4.815
+ $X2=2.1 $Y2=5.835
r62 13 30 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=2.1 $Y=4.815
+ $X2=2.1 $Y2=3.045
r63 7 21 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.472
+ $X2=2.175 $Y2=1.472
r64 7 9 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.07 $Y=1.385 $X2=2.07
+ $Y2=0.825
r65 2 15 300 $w=1.7e-07 $l=1.46833e-06 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=4.435 $X2=2.1 $Y2=5.835
r66 2 13 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=4.435 $X2=2.1 $Y2=4.815
r67 1 9 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%A_570_115# 1 2 9 11 12
r11 13 15 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.85 $Y=0.72
+ $X2=3.85 $Y2=0.825
r12 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.85 $Y2=0.72
r13 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.075 $Y2=0.635
r14 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.72
+ $X2=3.075 $Y2=0.635
r15 7 9 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.72 $X2=2.99
+ $Y2=0.825
r16 2 15 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.825
r17 1 9 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.825
.ends

