* File: sky130_osu_sc_12T_hs__and2_8.spice
* Created: Fri Nov 12 15:07:17 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__and2_8.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_8  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1008 A_110_115# N_A_M1008_g N_A_27_115#_M1008_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1004_d N_B_M1004_g A_110_115# N_GND_M1008_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_GND_M1004_d N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.09625 PD=0.83 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1003_d N_A_27_115#_M1009_g N_GND_M1009_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1012 N_Y_M1012_d N_A_27_115#_M1012_g N_GND_M1009_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1015 N_Y_M1012_d N_A_27_115#_M1015_g N_GND_M1015_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1016 N_Y_M1016_d N_A_27_115#_M1016_g N_GND_M1015_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1017 N_Y_M1016_d N_A_27_115#_M1017_g N_GND_M1017_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1018 N_Y_M1018_d N_A_27_115#_M1018_g N_GND_M1017_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1019 N_Y_M1018_d N_A_27_115#_M1019_g N_GND_M1019_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75004.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1013 N_VDD_M1013_d N_B_M1013_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_VDD_M1013_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1001_d N_A_27_115#_M1002_g N_VDD_M1002_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_VDD_M1002_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1005_d N_A_27_115#_M1006_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A_27_115#_M1007_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1007_d N_A_27_115#_M1010_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_A_27_115#_M1011_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1011_d N_A_27_115#_M1014_g N_VDD_M1014_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref N_GND_M1008_b N_VDD_M1000_b NWDIODE A=10.2897 P=14.11
pX21_noxref noxref_8 A A PROBETYPE=1
pX22_noxref noxref_9 B B PROBETYPE=1
pX23_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_8.pxi.spice"
*
.ends
*
*
