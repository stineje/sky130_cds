magic
tech sky130A
magscale 1 2
timestamp 1606864603
<< checkpaint >>
rect -1210 -1243 3112 2575
<< nwell >>
rect -10 581 1917 1341
<< nmos >>
rect 80 115 110 315
rect 270 115 300 263
rect 356 115 386 263
rect 546 115 576 315
rect 618 115 648 315
rect 738 115 768 315
rect 810 115 840 315
rect 896 115 926 315
rect 968 115 998 315
rect 1088 115 1118 315
rect 1160 115 1190 315
rect 1246 115 1276 315
rect 1436 115 1466 263
rect 1522 115 1552 263
rect 1712 115 1742 315
rect 1798 115 1828 315
<< pmos >>
rect 80 617 110 1217
rect 270 817 300 1217
rect 342 817 372 1217
rect 546 617 576 1217
rect 618 617 648 1217
rect 738 617 768 1217
rect 810 617 840 1217
rect 896 617 926 1217
rect 968 617 998 1217
rect 1088 617 1118 1217
rect 1160 617 1190 1217
rect 1246 617 1276 1217
rect 1436 817 1466 1217
rect 1508 817 1538 1217
rect 1712 617 1742 1217
rect 1798 617 1828 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 163 315
rect 110 131 121 267
rect 155 131 163 267
rect 493 267 546 315
rect 110 115 163 131
rect 217 199 270 263
rect 217 131 225 199
rect 259 131 270 199
rect 217 115 270 131
rect 300 199 356 263
rect 300 131 311 199
rect 345 131 356 199
rect 300 115 356 131
rect 386 199 439 263
rect 386 131 397 199
rect 431 131 439 199
rect 386 115 439 131
rect 493 131 501 267
rect 535 131 546 267
rect 493 115 546 131
rect 576 115 618 315
rect 648 267 738 315
rect 648 131 659 267
rect 727 131 738 267
rect 648 115 738 131
rect 768 115 810 315
rect 840 199 896 315
rect 840 131 851 199
rect 885 131 896 199
rect 840 115 896 131
rect 926 115 968 315
rect 998 267 1088 315
rect 998 131 1009 267
rect 1077 131 1088 267
rect 998 115 1088 131
rect 1118 115 1160 315
rect 1190 267 1246 315
rect 1190 131 1201 267
rect 1235 131 1246 267
rect 1190 115 1246 131
rect 1276 267 1329 315
rect 1276 131 1287 267
rect 1321 131 1329 267
rect 1276 115 1329 131
rect 1383 199 1436 263
rect 1383 131 1391 199
rect 1425 131 1436 199
rect 1383 115 1436 131
rect 1466 199 1522 263
rect 1466 131 1477 199
rect 1511 131 1522 199
rect 1466 115 1522 131
rect 1552 199 1605 263
rect 1552 131 1563 199
rect 1597 131 1605 199
rect 1552 115 1605 131
rect 1659 199 1712 315
rect 1659 131 1667 199
rect 1701 131 1712 199
rect 1659 115 1712 131
rect 1742 199 1798 315
rect 1742 131 1753 199
rect 1787 131 1798 199
rect 1742 115 1798 131
rect 1828 199 1881 315
rect 1828 131 1839 199
rect 1873 131 1881 199
rect 1828 115 1881 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 163 1217
rect 110 657 121 1201
rect 155 657 163 1201
rect 217 1201 270 1217
rect 217 861 225 1201
rect 259 861 270 1201
rect 217 817 270 861
rect 300 817 342 1217
rect 372 1201 425 1217
rect 372 861 383 1201
rect 417 861 425 1201
rect 372 817 425 861
rect 493 1201 546 1217
rect 110 617 163 657
rect 493 725 501 1201
rect 535 725 546 1201
rect 493 617 546 725
rect 576 617 618 1217
rect 648 1201 738 1217
rect 648 657 659 1201
rect 727 657 738 1201
rect 648 617 738 657
rect 768 617 810 1217
rect 840 1201 896 1217
rect 840 725 851 1201
rect 885 725 896 1201
rect 840 617 896 725
rect 926 617 968 1217
rect 998 1201 1088 1217
rect 998 725 1009 1201
rect 1077 725 1088 1201
rect 998 617 1088 725
rect 1118 617 1160 1217
rect 1190 1201 1246 1217
rect 1190 657 1201 1201
rect 1235 657 1246 1201
rect 1190 617 1246 657
rect 1276 1201 1329 1217
rect 1276 657 1287 1201
rect 1321 657 1329 1201
rect 1383 1201 1436 1217
rect 1383 861 1391 1201
rect 1425 861 1436 1201
rect 1383 817 1436 861
rect 1466 817 1508 1217
rect 1538 1201 1591 1217
rect 1538 861 1549 1201
rect 1583 861 1591 1201
rect 1538 817 1591 861
rect 1659 1201 1712 1217
rect 1659 861 1667 1201
rect 1701 861 1712 1201
rect 1276 617 1329 657
rect 1659 617 1712 861
rect 1742 1201 1798 1217
rect 1742 861 1753 1201
rect 1787 861 1798 1201
rect 1742 617 1798 861
rect 1828 1201 1881 1217
rect 1828 861 1839 1201
rect 1873 861 1881 1201
rect 1828 617 1881 861
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 225 131 259 199
rect 311 131 345 199
rect 397 131 431 199
rect 501 131 535 267
rect 659 131 727 267
rect 851 131 885 199
rect 1009 131 1077 267
rect 1201 131 1235 267
rect 1287 131 1321 267
rect 1391 131 1425 199
rect 1477 131 1511 199
rect 1563 131 1597 199
rect 1667 131 1701 199
rect 1753 131 1787 199
rect 1839 131 1873 199
<< pdiffc >>
rect 35 793 69 1201
rect 121 657 155 1201
rect 225 861 259 1201
rect 383 861 417 1201
rect 501 725 535 1201
rect 659 657 727 1201
rect 851 725 885 1201
rect 1009 725 1077 1201
rect 1201 657 1235 1201
rect 1287 657 1321 1201
rect 1391 861 1425 1201
rect 1549 861 1583 1201
rect 1667 861 1701 1201
rect 1753 861 1787 1201
rect 1839 861 1873 1201
<< psubdiff >>
rect 26 27 50 61
rect 84 27 108 61
rect 162 27 186 61
rect 220 27 244 61
rect 298 27 322 61
rect 356 27 380 61
rect 434 27 458 61
rect 492 27 516 61
rect 570 27 594 61
rect 628 27 652 61
rect 706 27 730 61
rect 764 27 788 61
rect 842 27 866 61
rect 900 27 924 61
rect 978 27 1002 61
rect 1036 27 1060 61
rect 1114 27 1138 61
rect 1172 27 1196 61
rect 1250 27 1274 61
rect 1308 27 1332 61
rect 1386 27 1410 61
rect 1444 27 1468 61
rect 1522 27 1546 61
rect 1580 27 1604 61
rect 1658 27 1682 61
rect 1716 27 1740 61
rect 1794 27 1818 61
rect 1852 27 1876 61
<< nsubdiff >>
rect 26 1271 50 1305
rect 84 1271 108 1305
rect 162 1271 186 1305
rect 220 1271 244 1305
rect 298 1271 322 1305
rect 356 1271 380 1305
rect 434 1271 458 1305
rect 492 1271 516 1305
rect 570 1271 594 1305
rect 628 1271 652 1305
rect 706 1271 730 1305
rect 764 1271 788 1305
rect 842 1271 866 1305
rect 900 1271 924 1305
rect 978 1271 1002 1305
rect 1036 1271 1060 1305
rect 1114 1271 1138 1305
rect 1172 1271 1196 1305
rect 1250 1271 1274 1305
rect 1308 1271 1332 1305
rect 1386 1271 1410 1305
rect 1444 1271 1468 1305
rect 1522 1271 1546 1305
rect 1580 1271 1604 1305
rect 1658 1271 1682 1305
rect 1716 1271 1740 1305
rect 1794 1271 1818 1305
rect 1852 1271 1876 1305
<< psubdiffcont >>
rect 50 27 84 61
rect 186 27 220 61
rect 322 27 356 61
rect 458 27 492 61
rect 594 27 628 61
rect 730 27 764 61
rect 866 27 900 61
rect 1002 27 1036 61
rect 1138 27 1172 61
rect 1274 27 1308 61
rect 1410 27 1444 61
rect 1546 27 1580 61
rect 1682 27 1716 61
rect 1818 27 1852 61
<< nsubdiffcont >>
rect 50 1271 84 1305
rect 186 1271 220 1305
rect 322 1271 356 1305
rect 458 1271 492 1305
rect 594 1271 628 1305
rect 730 1271 764 1305
rect 866 1271 900 1305
rect 1002 1271 1036 1305
rect 1138 1271 1172 1305
rect 1274 1271 1308 1305
rect 1410 1271 1444 1305
rect 1546 1271 1580 1305
rect 1682 1271 1716 1305
rect 1818 1271 1852 1305
<< poly >>
rect 80 1217 110 1243
rect 270 1217 300 1243
rect 342 1217 372 1243
rect 546 1217 576 1243
rect 618 1217 648 1243
rect 738 1217 768 1243
rect 810 1217 840 1243
rect 896 1217 926 1243
rect 968 1217 998 1243
rect 1088 1217 1118 1243
rect 1160 1217 1190 1243
rect 1246 1217 1276 1243
rect 1436 1217 1466 1243
rect 1508 1217 1538 1243
rect 1712 1217 1742 1243
rect 1798 1217 1828 1243
rect 80 494 110 617
rect 79 478 133 494
rect 79 444 89 478
rect 123 444 133 478
rect 79 428 133 444
rect 79 427 110 428
rect 80 315 110 427
rect 270 351 300 817
rect 342 584 372 817
rect 342 568 415 584
rect 342 534 371 568
rect 405 534 415 568
rect 342 518 415 534
rect 219 335 300 351
rect 219 301 229 335
rect 263 301 300 335
rect 219 285 300 301
rect 270 263 300 285
rect 356 263 386 518
rect 546 477 576 617
rect 618 586 648 617
rect 618 570 672 586
rect 618 536 628 570
rect 662 536 672 570
rect 618 520 672 536
rect 546 461 600 477
rect 738 475 768 617
rect 810 580 840 617
rect 896 580 926 617
rect 810 570 926 580
rect 810 536 842 570
rect 876 536 926 570
rect 810 526 926 536
rect 968 475 998 617
rect 1088 586 1118 617
rect 1064 570 1118 586
rect 1064 536 1074 570
rect 1108 536 1118 570
rect 1064 520 1118 536
rect 546 427 556 461
rect 590 427 600 461
rect 546 411 600 427
rect 642 445 1094 475
rect 546 315 576 411
rect 642 367 672 445
rect 1064 403 1094 445
rect 1160 471 1190 617
rect 1246 586 1276 617
rect 1246 570 1317 586
rect 1246 556 1273 570
rect 1257 536 1273 556
rect 1307 536 1317 570
rect 1257 520 1317 536
rect 1160 455 1214 471
rect 1160 421 1170 455
rect 1204 421 1214 455
rect 1160 405 1214 421
rect 618 337 672 367
rect 714 387 768 403
rect 714 353 724 387
rect 758 353 768 387
rect 714 337 768 353
rect 618 315 648 337
rect 738 315 768 337
rect 810 387 926 397
rect 810 353 842 387
rect 876 353 926 387
rect 810 343 926 353
rect 810 315 840 343
rect 896 315 926 343
rect 968 387 1022 403
rect 968 353 978 387
rect 1012 353 1022 387
rect 968 337 1022 353
rect 1064 387 1118 403
rect 1064 353 1074 387
rect 1108 353 1118 387
rect 1064 337 1118 353
rect 968 315 998 337
rect 1088 315 1118 337
rect 1160 315 1190 405
rect 1257 367 1287 520
rect 1436 403 1466 817
rect 1246 337 1287 367
rect 1399 387 1466 403
rect 1399 353 1409 387
rect 1443 353 1466 387
rect 1399 337 1466 353
rect 1246 315 1276 337
rect 1423 336 1466 337
rect 1436 263 1466 336
rect 1508 351 1538 817
rect 1712 601 1742 617
rect 1702 571 1742 601
rect 1702 471 1732 571
rect 1798 512 1828 617
rect 1677 455 1732 471
rect 1677 421 1687 455
rect 1721 421 1732 455
rect 1774 496 1828 512
rect 1774 462 1784 496
rect 1818 462 1828 496
rect 1774 446 1828 462
rect 1677 405 1732 421
rect 1702 360 1732 405
rect 1508 335 1589 351
rect 1508 301 1545 335
rect 1579 301 1589 335
rect 1702 330 1742 360
rect 1712 315 1742 330
rect 1798 315 1828 446
rect 1508 285 1589 301
rect 1522 263 1552 285
rect 80 89 110 115
rect 270 89 300 115
rect 356 89 386 115
rect 546 89 576 115
rect 618 89 648 115
rect 738 89 768 115
rect 810 89 840 115
rect 896 89 926 115
rect 968 89 998 115
rect 1088 89 1118 115
rect 1160 89 1190 115
rect 1246 89 1276 115
rect 1436 89 1466 115
rect 1522 89 1552 115
rect 1712 89 1742 115
rect 1798 89 1828 115
<< polycont >>
rect 89 444 123 478
rect 371 534 405 568
rect 229 301 263 335
rect 628 536 662 570
rect 842 536 876 570
rect 1074 536 1108 570
rect 556 427 590 461
rect 1273 536 1307 570
rect 1170 421 1204 455
rect 724 353 758 387
rect 842 353 876 387
rect 978 353 1012 387
rect 1074 353 1108 387
rect 1409 353 1443 387
rect 1687 421 1721 455
rect 1784 462 1818 496
rect 1545 301 1579 335
<< locali >>
rect 0 1311 1914 1332
rect 0 1271 50 1311
rect 84 1271 186 1311
rect 220 1271 322 1311
rect 356 1271 458 1311
rect 492 1271 594 1311
rect 628 1271 730 1311
rect 764 1271 866 1311
rect 900 1271 1002 1311
rect 1036 1271 1138 1311
rect 1172 1271 1274 1311
rect 1308 1271 1410 1311
rect 1444 1271 1546 1311
rect 1580 1271 1682 1311
rect 1716 1271 1818 1311
rect 1852 1271 1914 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 47 494 81 649
rect 121 565 155 657
rect 225 1201 259 1217
rect 121 531 191 565
rect 47 478 123 494
rect 47 444 89 478
rect 89 428 123 444
rect 157 335 191 531
rect 225 421 259 861
rect 383 1201 417 1271
rect 383 845 417 861
rect 501 1201 535 1271
rect 501 709 535 725
rect 659 1201 727 1217
rect 851 1201 885 1271
rect 851 709 885 725
rect 1009 1201 1077 1217
rect 659 654 727 657
rect 1009 654 1077 725
rect 405 620 727 654
rect 910 620 1077 654
rect 1201 1201 1235 1271
rect 1201 641 1235 657
rect 1287 1201 1321 1217
rect 1391 1201 1425 1217
rect 1391 773 1425 861
rect 1549 1201 1583 1271
rect 1549 845 1583 861
rect 1667 1201 1701 1217
rect 1391 739 1511 773
rect 1287 654 1321 657
rect 1287 620 1377 654
rect 405 584 439 620
rect 371 568 439 584
rect 405 534 439 568
rect 371 518 439 534
rect 225 387 345 421
rect 229 335 263 351
rect 121 301 229 335
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 301
rect 121 115 155 131
rect 225 199 259 215
rect 225 61 259 131
rect 311 199 345 353
rect 405 370 439 518
rect 628 570 662 586
rect 628 535 662 536
rect 842 570 876 586
rect 662 501 758 535
rect 556 461 590 477
rect 556 411 590 427
rect 724 387 758 501
rect 842 387 876 536
rect 405 336 690 370
rect 724 337 758 353
rect 842 337 876 353
rect 910 387 944 620
rect 1074 570 1108 586
rect 1074 535 1108 536
rect 656 283 690 336
rect 910 303 944 353
rect 978 501 1074 535
rect 1273 570 1307 586
rect 1273 535 1307 536
rect 978 387 1012 501
rect 1341 455 1377 620
rect 1154 421 1170 455
rect 1204 421 1220 455
rect 1287 421 1377 455
rect 1477 455 1511 739
rect 1667 609 1701 861
rect 1753 1201 1787 1271
rect 1753 845 1787 861
rect 1839 1201 1873 1217
rect 1839 683 1873 861
rect 1872 666 1873 683
rect 1872 649 1896 666
rect 1839 632 1896 649
rect 1667 570 1701 575
rect 1667 536 1818 570
rect 1784 496 1818 536
rect 1477 421 1687 455
rect 1721 421 1737 455
rect 1287 387 1321 421
rect 1058 353 1074 387
rect 1108 353 1321 387
rect 978 337 1012 353
rect 501 267 535 283
rect 311 115 345 131
rect 397 199 431 215
rect 397 61 431 131
rect 656 267 727 283
rect 910 269 1077 303
rect 656 249 659 267
rect 501 61 535 131
rect 1009 267 1077 269
rect 659 115 727 131
rect 851 199 885 215
rect 851 61 885 131
rect 1009 115 1077 131
rect 1201 267 1235 283
rect 1201 61 1235 131
rect 1287 267 1321 353
rect 1409 387 1443 403
rect 1409 337 1443 353
rect 1287 115 1321 131
rect 1391 199 1425 215
rect 1391 61 1425 131
rect 1477 199 1511 421
rect 1784 387 1818 462
rect 1667 353 1818 387
rect 1545 335 1579 351
rect 1477 115 1511 131
rect 1563 199 1597 215
rect 1563 61 1597 131
rect 1667 199 1701 353
rect 1862 320 1896 632
rect 1839 286 1896 320
rect 1667 115 1701 131
rect 1753 199 1787 215
rect 1753 61 1787 131
rect 1839 199 1873 286
rect 1839 115 1873 131
rect 0 21 50 61
rect 84 21 186 61
rect 220 21 322 61
rect 356 21 458 61
rect 492 21 594 61
rect 628 21 730 61
rect 764 21 866 61
rect 900 21 1002 61
rect 1036 21 1138 61
rect 1172 21 1274 61
rect 1308 21 1410 61
rect 1444 21 1546 61
rect 1580 21 1682 61
rect 1716 21 1818 61
rect 1852 21 1914 61
rect 0 0 1914 21
<< viali >>
rect 50 1305 84 1311
rect 50 1277 84 1305
rect 186 1305 220 1311
rect 186 1277 220 1305
rect 322 1305 356 1311
rect 322 1277 356 1305
rect 458 1305 492 1311
rect 458 1277 492 1305
rect 594 1305 628 1311
rect 594 1277 628 1305
rect 730 1305 764 1311
rect 730 1277 764 1305
rect 866 1305 900 1311
rect 866 1277 900 1305
rect 1002 1305 1036 1311
rect 1002 1277 1036 1305
rect 1138 1305 1172 1311
rect 1138 1277 1172 1305
rect 1274 1305 1308 1311
rect 1274 1277 1308 1305
rect 1410 1305 1444 1311
rect 1410 1277 1444 1305
rect 1546 1305 1580 1311
rect 1546 1277 1580 1305
rect 1682 1305 1716 1311
rect 1682 1277 1716 1305
rect 1818 1305 1852 1311
rect 1818 1277 1852 1305
rect 47 649 81 683
rect 311 353 345 387
rect 229 301 263 313
rect 229 279 263 301
rect 628 501 662 535
rect 556 427 590 461
rect 824 353 842 387
rect 842 353 858 387
rect 910 353 944 387
rect 1074 501 1108 535
rect 1273 501 1307 535
rect 1170 421 1204 455
rect 1838 649 1872 683
rect 1667 575 1701 609
rect 1687 421 1721 455
rect 1409 353 1443 387
rect 1545 301 1579 313
rect 1545 279 1579 301
rect 50 27 84 55
rect 50 21 84 27
rect 186 27 220 55
rect 186 21 220 27
rect 322 27 356 55
rect 322 21 356 27
rect 458 27 492 55
rect 458 21 492 27
rect 594 27 628 55
rect 594 21 628 27
rect 730 27 764 55
rect 730 21 764 27
rect 866 27 900 55
rect 866 21 900 27
rect 1002 27 1036 55
rect 1002 21 1036 27
rect 1138 27 1172 55
rect 1138 21 1172 27
rect 1274 27 1308 55
rect 1274 21 1308 27
rect 1410 27 1444 55
rect 1410 21 1444 27
rect 1546 27 1580 55
rect 1546 21 1580 27
rect 1682 27 1716 55
rect 1682 21 1716 27
rect 1818 27 1852 55
rect 1818 21 1852 27
<< metal1 >>
rect 0 1311 1914 1332
rect 0 1277 50 1311
rect 84 1277 186 1311
rect 220 1277 322 1311
rect 356 1277 458 1311
rect 492 1277 594 1311
rect 628 1277 730 1311
rect 764 1277 866 1311
rect 900 1277 1002 1311
rect 1036 1277 1138 1311
rect 1172 1277 1274 1311
rect 1308 1277 1410 1311
rect 1444 1277 1546 1311
rect 1580 1277 1682 1311
rect 1716 1277 1818 1311
rect 1852 1277 1914 1311
rect 0 1271 1914 1277
rect 35 683 93 689
rect 1826 683 1884 689
rect 35 649 47 683
rect 81 649 127 683
rect 1804 649 1838 683
rect 1872 649 1884 683
rect 35 643 93 649
rect 1826 643 1884 649
rect 1655 609 1713 615
rect 1632 575 1667 609
rect 1701 575 1713 609
rect 1655 569 1713 575
rect 616 535 674 541
rect 1062 535 1120 541
rect 1261 535 1319 541
rect 616 501 628 535
rect 662 501 1074 535
rect 1108 501 1273 535
rect 1307 501 1319 535
rect 616 495 674 501
rect 1062 495 1120 501
rect 1261 495 1319 501
rect 544 461 602 467
rect 544 427 556 461
rect 590 427 624 461
rect 1158 455 1216 461
rect 1675 455 1733 461
rect 544 421 602 427
rect 1158 421 1170 455
rect 1204 421 1687 455
rect 1721 421 1733 455
rect 1158 415 1216 421
rect 1675 415 1733 421
rect 299 387 357 393
rect 812 387 870 393
rect 299 353 311 387
rect 345 353 824 387
rect 858 353 870 387
rect 299 347 357 353
rect 812 347 870 353
rect 898 387 956 393
rect 1397 387 1455 393
rect 898 353 910 387
rect 944 353 1409 387
rect 1443 353 1455 387
rect 898 347 956 353
rect 1397 347 1455 353
rect 217 313 275 319
rect 1533 313 1591 319
rect 217 279 229 313
rect 263 279 1545 313
rect 1579 279 1591 313
rect 217 273 275 279
rect 1533 273 1591 279
rect 0 55 1914 61
rect 0 21 50 55
rect 84 21 186 55
rect 220 21 322 55
rect 356 21 458 55
rect 492 21 594 55
rect 628 21 730 55
rect 764 21 866 55
rect 900 21 1002 55
rect 1036 21 1138 55
rect 1172 21 1274 55
rect 1308 21 1410 55
rect 1444 21 1546 55
rect 1580 21 1682 55
rect 1716 21 1818 55
rect 1852 21 1914 55
rect 0 0 1914 21
<< labels >>
rlabel metal1 65 666 65 666 1 RN
port 1 n
rlabel metal1 573 444 573 444 1 D
port 2 n
rlabel metal1 1290 518 1290 518 1 CK
port 3 n
rlabel metal1 1855 666 1855 666 1 Q
port 4 n
rlabel metal1 1685 592 1685 592 1 QN
port 5 n
rlabel viali 67 48 67 48 1 gnd
rlabel viali 67 1284 67 1284 1 vdd
<< end >>
