* File: sky130_osu_sc_18T_ms__dffsr_l.pxi.spice
* Created: Fri Nov 12 14:03:24 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%GND N_GND_M1017_s N_GND_M1032_s N_GND_M1001_d
+ N_GND_M1005_s N_GND_M1021_d N_GND_M1006_d N_GND_M1013_s N_GND_M1023_d
+ N_GND_M1007_d N_GND_M1017_b N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_14_p
+ N_GND_c_47_p N_GND_c_48_p N_GND_c_88_p N_GND_c_49_p N_GND_c_107_p N_GND_c_50_p
+ N_GND_c_112_p N_GND_c_51_p N_GND_c_17_p N_GND_c_18_p N_GND_c_189_p
+ N_GND_c_190_p GND N_GND_c_5_p PM_SKY130_OSU_SC_18T_MS__DFFSR_L%GND
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%VDD N_VDD_M1019_s N_VDD_M1000_d N_VDD_M1008_s
+ N_VDD_M1024_d N_VDD_M1009_d N_VDD_M1014_d N_VDD_M1028_d N_VDD_M1019_b
+ N_VDD_c_249_p N_VDD_c_250_p N_VDD_c_268_p N_VDD_c_283_p N_VDD_c_284_p
+ N_VDD_c_292_p N_VDD_c_277_p N_VDD_c_302_p N_VDD_c_278_p N_VDD_c_307_p
+ N_VDD_c_271_p N_VDD_c_261_p N_VDD_c_345_p N_VDD_c_362_p VDD N_VDD_c_251_p
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%VDD
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%RN N_RN_M1017_g N_RN_c_397_n N_RN_M1019_g
+ N_RN_c_399_n N_RN_c_400_n RN PM_SKY130_OSU_SC_18T_MS__DFFSR_L%RN
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_110_115# N_A_110_115#_M1017_d
+ N_A_110_115#_M1019_d N_A_110_115#_c_432_n N_A_110_115#_M1016_g
+ N_A_110_115#_c_434_n N_A_110_115#_M1032_g N_A_110_115#_c_438_n
+ N_A_110_115#_M1023_g N_A_110_115#_M1004_g N_A_110_115#_c_443_n
+ N_A_110_115#_c_444_n N_A_110_115#_c_445_n N_A_110_115#_c_447_n
+ N_A_110_115#_c_448_n N_A_110_115#_c_450_n N_A_110_115#_c_454_n
+ N_A_110_115#_c_455_n N_A_110_115#_c_456_n N_A_110_115#_c_457_n
+ N_A_110_115#_c_458_n N_A_110_115#_c_459_n N_A_110_115#_c_461_n
+ N_A_110_115#_c_463_n N_A_110_115#_c_475_n N_A_110_115#_c_477_n
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_110_115#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%SN N_SN_M1000_g N_SN_M1015_g N_SN_M1002_g
+ N_SN_M1035_g N_SN_c_649_n N_SN_c_650_n N_SN_c_651_n N_SN_c_652_n N_SN_c_653_n
+ N_SN_c_654_n N_SN_c_655_n N_SN_c_656_n N_SN_c_657_n N_SN_c_658_n SN
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%SN
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_432_520# N_A_432_520#_M1033_d
+ N_A_432_520#_M1034_d N_A_432_520#_M1001_g N_A_432_520#_M1003_g
+ N_A_432_520#_c_816_n N_A_432_520#_c_817_n N_A_432_520#_c_818_n
+ N_A_432_520#_c_821_n N_A_432_520#_c_833_n N_A_432_520#_c_863_n
+ N_A_432_520#_c_822_n N_A_432_520#_c_823_n N_A_432_520#_c_836_n
+ N_A_432_520#_c_844_n PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_432_520#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%D N_D_M1005_g N_D_M1008_g N_D_c_907_n
+ N_D_c_908_n D PM_SKY130_OSU_SC_18T_MS__DFFSR_L%D
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%CK N_CK_M1034_g N_CK_M1030_g N_CK_M1022_g
+ N_CK_M1020_g N_CK_M1011_g N_CK_c_941_n N_CK_M1012_g N_CK_c_942_n N_CK_c_943_n
+ N_CK_c_944_n N_CK_c_945_n N_CK_c_948_n N_CK_c_949_n N_CK_c_952_n N_CK_c_953_n
+ N_CK_c_958_n N_CK_c_959_n N_CK_c_960_n N_CK_c_961_n N_CK_c_962_n N_CK_c_963_n
+ N_CK_c_964_n N_CK_c_965_n N_CK_c_966_n N_CK_c_967_n N_CK_c_968_n N_CK_c_969_n
+ N_CK_c_970_n CK PM_SKY130_OSU_SC_18T_MS__DFFSR_L%CK
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_217_617# N_A_217_617#_M1032_d
+ N_A_217_617#_M1016_s N_A_217_617#_M1021_g N_A_217_617#_M1024_g
+ N_A_217_617#_c_1178_n N_A_217_617#_c_1180_n N_A_217_617#_c_1181_n
+ N_A_217_617#_c_1182_n N_A_217_617#_M1026_g N_A_217_617#_M1027_g
+ N_A_217_617#_c_1187_n N_A_217_617#_c_1188_n N_A_217_617#_c_1189_n
+ N_A_217_617#_c_1190_n N_A_217_617#_c_1193_n N_A_217_617#_c_1194_n
+ N_A_217_617#_c_1196_n N_A_217_617#_c_1197_n N_A_217_617#_c_1247_n
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_217_617#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_704_89# N_A_704_89#_M1011_d
+ N_A_704_89#_M1012_d N_A_704_89#_c_1338_n N_A_704_89#_M1033_g
+ N_A_704_89#_c_1341_n N_A_704_89#_c_1342_n N_A_704_89#_c_1343_n
+ N_A_704_89#_M1031_g N_A_704_89#_c_1345_n N_A_704_89#_M1025_g
+ N_A_704_89#_c_1347_n N_A_704_89#_c_1348_n N_A_704_89#_M1018_g
+ N_A_704_89#_c_1349_n N_A_704_89#_c_1350_n N_A_704_89#_c_1351_n
+ N_A_704_89#_c_1352_n N_A_704_89#_c_1353_n N_A_704_89#_c_1356_n
+ N_A_704_89#_c_1358_n N_A_704_89#_c_1363_n N_A_704_89#_c_1373_n
+ N_A_704_89#_c_1364_n N_A_704_89#_c_1365_n N_A_704_89#_c_1366_n
+ N_A_704_89#_c_1377_n PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_704_89#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_1246_89# N_A_1246_89#_M1002_d
+ N_A_1246_89#_M1004_d N_A_1246_89#_M1006_g N_A_1246_89#_M1009_g
+ N_A_1246_89#_M1007_g N_A_1246_89#_M1028_g N_A_1246_89#_c_1539_n
+ N_A_1246_89#_c_1540_n N_A_1246_89#_c_1541_n N_A_1246_89#_c_1542_n
+ N_A_1246_89#_c_1543_n N_A_1246_89#_c_1544_n N_A_1246_89#_c_1545_n
+ N_A_1246_89#_c_1546_n N_A_1246_89#_c_1549_n N_A_1246_89#_c_1550_n
+ N_A_1246_89#_c_1551_n N_A_1246_89#_c_1552_n N_A_1246_89#_c_1553_n
+ N_A_1246_89#_c_1554_n PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_1246_89#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_1084_115# N_A_1084_115#_M1022_d
+ N_A_1084_115#_M1025_d N_A_1084_115#_c_1705_n N_A_1084_115#_c_1706_n
+ N_A_1084_115#_M1013_g N_A_1084_115#_M1014_g N_A_1084_115#_c_1710_n
+ N_A_1084_115#_c_1712_n N_A_1084_115#_c_1713_n N_A_1084_115#_c_1738_n
+ N_A_1084_115#_c_1739_n N_A_1084_115#_c_1757_n N_A_1084_115#_c_1805_n
+ N_A_1084_115#_c_1714_n N_A_1084_115#_c_1730_n N_A_1084_115#_c_1717_n
+ N_A_1084_115#_c_1719_n N_A_1084_115#_c_1722_n N_A_1084_115#_c_1723_n
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_1084_115#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%QN N_QN_M1007_s N_QN_M1028_s N_QN_M1010_g
+ N_QN_M1029_g N_QN_c_1866_n N_QN_c_1867_n N_QN_c_1871_n N_QN_c_1872_n
+ N_QN_c_1873_n N_QN_c_1874_n N_QN_c_1875_n N_QN_c_1876_n QN
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%QN
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_300_617# N_A_300_617#_M1016_d
+ N_A_300_617#_M1003_d N_A_300_617#_c_1946_n N_A_300_617#_c_1949_n
+ N_A_300_617#_c_1960_n N_A_300_617#_c_1952_n
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_300_617#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_1469_617# N_A_1469_617#_M1014_s
+ N_A_1469_617#_M1035_d N_A_1469_617#_c_1970_n N_A_1469_617#_c_1973_n
+ N_A_1469_617#_c_1982_n N_A_1469_617#_c_1975_n
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%A_1469_617#
x_PM_SKY130_OSU_SC_18T_MS__DFFSR_L%Q N_Q_M1010_d N_Q_M1029_d N_Q_c_1989_n
+ N_Q_c_1993_n N_Q_c_1991_n N_Q_c_1992_n N_Q_c_1997_n Q
+ PM_SKY130_OSU_SC_18T_MS__DFFSR_L%Q
cc_1 N_GND_M1017_b N_RN_M1017_g 0.0636982f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_RN_M1017_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_RN_M1017_g 0.00606474f $X=1.135 $Y=0.152 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_RN_M1017_g 0.00392369f $X=1.22 $Y=0.825 $X2=0.475 $Y2=1.075
cc_5 N_GND_c_5_p N_RN_M1017_g 0.00468827f $X=9.855 $Y=0.19 $X2=0.475 $Y2=1.075
cc_6 N_GND_M1017_b N_RN_c_397_n 0.0367952f $X=-0.05 $Y=0 $X2=0.475 $Y2=2.47
cc_7 N_GND_M1017_b N_RN_M1019_g 0.0318003f $X=-0.05 $Y=0 $X2=0.475 $Y2=4.585
cc_8 N_GND_M1017_b N_RN_c_399_n 0.0149094f $X=-0.05 $Y=0 $X2=0.32 $Y2=3.33
cc_9 N_GND_M1017_b N_RN_c_400_n 0.020318f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.305
cc_10 N_GND_M1017_b N_A_110_115#_c_432_n 0.0591015f $X=-0.05 $Y=0 $X2=1.29
+ $Y2=2.745
cc_11 N_GND_M1017_b N_A_110_115#_M1016_g 5.04534e-19 $X=-0.05 $Y=0 $X2=1.425
+ $Y2=4.585
cc_12 N_GND_M1017_b N_A_110_115#_c_434_n 0.0188414f $X=-0.05 $Y=0 $X2=1.435
+ $Y2=1.425
cc_13 N_GND_c_4_p N_A_110_115#_c_434_n 0.00713292f $X=1.22 $Y=0.825 $X2=1.435
+ $Y2=1.425
cc_14 N_GND_c_14_p N_A_110_115#_c_434_n 0.00606474f $X=2.415 $Y=0.152 $X2=1.435
+ $Y2=1.425
cc_15 N_GND_c_5_p N_A_110_115#_c_434_n 0.00468827f $X=9.855 $Y=0.19 $X2=1.435
+ $Y2=1.425
cc_16 N_GND_M1017_b N_A_110_115#_c_438_n 0.0187247f $X=-0.05 $Y=0 $X2=8.535
+ $Y2=1.425
cc_17 N_GND_c_17_p N_A_110_115#_c_438_n 0.00606474f $X=8.665 $Y=0.152 $X2=8.535
+ $Y2=1.425
cc_18 N_GND_c_18_p N_A_110_115#_c_438_n 0.00713292f $X=8.75 $Y=0.825 $X2=8.535
+ $Y2=1.425
cc_19 N_GND_c_5_p N_A_110_115#_c_438_n 0.00468827f $X=9.855 $Y=0.19 $X2=8.535
+ $Y2=1.425
cc_20 N_GND_M1017_b N_A_110_115#_M1004_g 5.06723e-19 $X=-0.05 $Y=0 $X2=8.545
+ $Y2=4.585
cc_21 N_GND_M1017_b N_A_110_115#_c_443_n 0.060764f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=2.745
cc_22 N_GND_M1017_b N_A_110_115#_c_444_n 0.0211399f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=2.82
cc_23 N_GND_M1017_b N_A_110_115#_c_445_n 0.0420101f $X=-0.05 $Y=0 $X2=1.29
+ $Y2=1.59
cc_24 N_GND_c_4_p N_A_110_115#_c_445_n 0.00122958f $X=1.22 $Y=0.825 $X2=1.29
+ $Y2=1.59
cc_25 N_GND_M1017_b N_A_110_115#_c_447_n 0.0303251f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=2.82
cc_26 N_GND_M1017_b N_A_110_115#_c_448_n 0.0484075f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=1.59
cc_27 N_GND_c_18_p N_A_110_115#_c_448_n 0.00254087f $X=8.75 $Y=0.825 $X2=8.8
+ $Y2=1.59
cc_28 N_GND_M1017_b N_A_110_115#_c_450_n 0.00156053f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=0.825
cc_29 N_GND_c_3_p N_A_110_115#_c_450_n 0.00757793f $X=1.135 $Y=0.152 $X2=0.69
+ $Y2=0.825
cc_30 N_GND_c_4_p N_A_110_115#_c_450_n 0.0209197f $X=1.22 $Y=0.825 $X2=0.69
+ $Y2=0.825
cc_31 N_GND_c_5_p N_A_110_115#_c_450_n 0.00476261f $X=9.855 $Y=0.19 $X2=0.69
+ $Y2=0.825
cc_32 N_GND_M1017_b N_A_110_115#_c_454_n 0.00214428f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=3.455
cc_33 N_GND_M1017_b N_A_110_115#_c_455_n 0.021684f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.655
cc_34 N_GND_M1017_b N_A_110_115#_c_456_n 0.0093348f $X=-0.05 $Y=0 $X2=1.145
+ $Y2=1.59
cc_35 N_GND_M1017_b N_A_110_115#_c_457_n 0.0126143f $X=-0.05 $Y=0 $X2=0.955
+ $Y2=1.59
cc_36 N_GND_M1017_b N_A_110_115#_c_458_n 0.0161505f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.74
cc_37 N_GND_M1017_b N_A_110_115#_c_459_n 0.00245576f $X=-0.05 $Y=0 $X2=1.23
+ $Y2=1.59
cc_38 N_GND_c_4_p N_A_110_115#_c_459_n 0.00596498f $X=1.22 $Y=0.825 $X2=1.23
+ $Y2=1.59
cc_39 N_GND_M1017_b N_A_110_115#_c_461_n 0.00578126f $X=-0.05 $Y=0 $X2=8.86
+ $Y2=1.48
cc_40 N_GND_c_18_p N_A_110_115#_c_461_n 0.00402542f $X=8.75 $Y=0.825 $X2=8.86
+ $Y2=1.48
cc_41 N_GND_M1001_d N_A_110_115#_c_463_n 0.00506015f $X=2.36 $Y=0.575 $X2=8.715
+ $Y2=1.48
cc_42 N_GND_M1005_s N_A_110_115#_c_463_n 0.00506021f $X=2.895 $Y=0.575 $X2=8.715
+ $Y2=1.48
cc_43 N_GND_M1021_d N_A_110_115#_c_463_n 0.0109039f $X=4.63 $Y=0.575 $X2=8.715
+ $Y2=1.48
cc_44 N_GND_M1006_d N_A_110_115#_c_463_n 0.00557645f $X=6.38 $Y=0.575 $X2=8.715
+ $Y2=1.48
cc_45 N_GND_M1013_s N_A_110_115#_c_463_n 0.00564702f $X=7.345 $Y=0.575 $X2=8.715
+ $Y2=1.48
cc_46 N_GND_M1017_b N_A_110_115#_c_463_n 0.0324773f $X=-0.05 $Y=0 $X2=8.715
+ $Y2=1.48
cc_47 N_GND_c_47_p N_A_110_115#_c_463_n 0.0118179f $X=2.5 $Y=0.825 $X2=8.715
+ $Y2=1.48
cc_48 N_GND_c_48_p N_A_110_115#_c_463_n 0.0118117f $X=3.02 $Y=0.825 $X2=8.715
+ $Y2=1.48
cc_49 N_GND_c_49_p N_A_110_115#_c_463_n 0.00558854f $X=4.77 $Y=0.825 $X2=8.715
+ $Y2=1.48
cc_50 N_GND_c_50_p N_A_110_115#_c_463_n 0.0119903f $X=6.52 $Y=0.825 $X2=8.715
+ $Y2=1.48
cc_51 N_GND_c_51_p N_A_110_115#_c_463_n 0.0139059f $X=7.47 $Y=0.825 $X2=8.715
+ $Y2=1.48
cc_52 N_GND_c_18_p N_A_110_115#_c_463_n 0.00182727f $X=8.75 $Y=0.825 $X2=8.715
+ $Y2=1.48
cc_53 N_GND_M1017_b N_A_110_115#_c_475_n 0.00666043f $X=-0.05 $Y=0 $X2=1.375
+ $Y2=1.48
cc_54 N_GND_c_4_p N_A_110_115#_c_475_n 0.00459186f $X=1.22 $Y=0.825 $X2=1.375
+ $Y2=1.48
cc_55 N_GND_M1017_b N_A_110_115#_c_477_n 0.00874177f $X=-0.05 $Y=0 $X2=8.86
+ $Y2=1.48
cc_56 N_GND_c_18_p N_A_110_115#_c_477_n 0.00334239f $X=8.75 $Y=0.825 $X2=8.86
+ $Y2=1.48
cc_57 N_GND_M1017_b N_SN_M1000_g 0.0180465f $X=-0.05 $Y=0 $X2=1.855 $Y2=4.585
cc_58 N_GND_M1017_b N_SN_M1015_g 0.0219538f $X=-0.05 $Y=0 $X2=1.925 $Y2=1.075
cc_59 N_GND_c_14_p N_SN_M1015_g 0.00606474f $X=2.415 $Y=0.152 $X2=1.925
+ $Y2=1.075
cc_60 N_GND_c_5_p N_SN_M1015_g 0.00468827f $X=9.855 $Y=0.19 $X2=1.925 $Y2=1.075
cc_61 N_GND_M1017_b N_SN_M1002_g 0.0426369f $X=-0.05 $Y=0 $X2=8.045 $Y2=1.075
cc_62 N_GND_c_17_p N_SN_M1002_g 0.00606474f $X=8.665 $Y=0.152 $X2=8.045
+ $Y2=1.075
cc_63 N_GND_c_5_p N_SN_M1002_g 0.00468827f $X=9.855 $Y=0.19 $X2=8.045 $Y2=1.075
cc_64 N_GND_M1017_b N_SN_M1035_g 0.0296048f $X=-0.05 $Y=0 $X2=8.115 $Y2=4.585
cc_65 N_GND_M1017_b N_SN_c_649_n 0.0343303f $X=-0.05 $Y=0 $X2=1.71 $Y2=2.37
cc_66 N_GND_M1017_b N_SN_c_650_n 0.0152246f $X=-0.05 $Y=0 $X2=1.752 $Y2=2.205
cc_67 N_GND_M1017_b N_SN_c_651_n 0.0125147f $X=-0.05 $Y=0 $X2=1.89 $Y2=1.925
cc_68 N_GND_M1017_b N_SN_c_652_n 0.0336181f $X=-0.05 $Y=0 $X2=8.025 $Y2=2.255
cc_69 N_GND_M1017_b N_SN_c_653_n 0.00274437f $X=-0.05 $Y=0 $X2=1.71 $Y2=2.96
cc_70 N_GND_M1017_b N_SN_c_654_n 0.00920532f $X=-0.05 $Y=0 $X2=7.935 $Y2=2.96
cc_71 N_GND_M1017_b N_SN_c_655_n 0.00222947f $X=-0.05 $Y=0 $X2=1.71 $Y2=2.37
cc_72 N_GND_M1017_b N_SN_c_656_n 0.00365816f $X=-0.05 $Y=0 $X2=8.025 $Y2=2.255
cc_73 N_GND_M1017_b N_SN_c_657_n 0.0543271f $X=-0.05 $Y=0 $X2=7.79 $Y2=2.96
cc_74 N_GND_M1017_b N_SN_c_658_n 0.00107924f $X=-0.05 $Y=0 $X2=1.855 $Y2=2.96
cc_75 N_GND_M1017_b SN 0.00268604f $X=-0.05 $Y=0 $X2=7.935 $Y2=2.96
cc_76 N_GND_M1017_b N_A_432_520#_M1001_g 0.0754451f $X=-0.05 $Y=0 $X2=2.285
+ $Y2=1.075
cc_77 N_GND_c_14_p N_A_432_520#_M1001_g 0.00606474f $X=2.415 $Y=0.152 $X2=2.285
+ $Y2=1.075
cc_78 N_GND_c_47_p N_A_432_520#_M1001_g 0.00715019f $X=2.5 $Y=0.825 $X2=2.285
+ $Y2=1.075
cc_79 N_GND_c_5_p N_A_432_520#_M1001_g 0.00468827f $X=9.855 $Y=0.19 $X2=2.285
+ $Y2=1.075
cc_80 N_GND_M1017_b N_A_432_520#_c_816_n 0.0343446f $X=-0.05 $Y=0 $X2=2.295
+ $Y2=2.765
cc_81 N_GND_M1017_b N_A_432_520#_c_817_n 0.0239207f $X=-0.05 $Y=0 $X2=2.295
+ $Y2=2.765
cc_82 N_GND_M1017_b N_A_432_520#_c_818_n 0.0278215f $X=-0.05 $Y=0 $X2=3.71
+ $Y2=1.765
cc_83 N_GND_c_47_p N_A_432_520#_c_818_n 0.00673409f $X=2.5 $Y=0.825 $X2=3.71
+ $Y2=1.765
cc_84 N_GND_c_48_p N_A_432_520#_c_818_n 0.00673409f $X=3.02 $Y=0.825 $X2=3.71
+ $Y2=1.765
cc_85 N_GND_M1017_b N_A_432_520#_c_821_n 0.00154034f $X=-0.05 $Y=0 $X2=2.38
+ $Y2=1.765
cc_86 N_GND_M1017_b N_A_432_520#_c_822_n 0.00198494f $X=-0.05 $Y=0 $X2=3.795
+ $Y2=1.68
cc_87 N_GND_M1017_b N_A_432_520#_c_823_n 0.00313975f $X=-0.05 $Y=0 $X2=3.895
+ $Y2=0.825
cc_88 N_GND_c_88_p N_A_432_520#_c_823_n 0.0149718f $X=4.685 $Y=0.152 $X2=3.895
+ $Y2=0.825
cc_89 N_GND_c_5_p N_A_432_520#_c_823_n 0.00958198f $X=9.855 $Y=0.19 $X2=3.895
+ $Y2=0.825
cc_90 N_GND_M1017_b N_D_M1005_g 0.0440753f $X=-0.05 $Y=0 $X2=3.235 $Y2=1.075
cc_91 N_GND_c_48_p N_D_M1005_g 0.0071489f $X=3.02 $Y=0.825 $X2=3.235 $Y2=1.075
cc_92 N_GND_c_88_p N_D_M1005_g 0.00606474f $X=4.685 $Y=0.152 $X2=3.235 $Y2=1.075
cc_93 N_GND_c_5_p N_D_M1005_g 0.00468827f $X=9.855 $Y=0.19 $X2=3.235 $Y2=1.075
cc_94 N_GND_M1017_b N_D_M1008_g 0.0445147f $X=-0.05 $Y=0 $X2=3.235 $Y2=4.585
cc_95 N_GND_M1017_b N_D_c_907_n 0.0337053f $X=-0.05 $Y=0 $X2=3.295 $Y2=2.22
cc_96 N_GND_M1017_b N_D_c_908_n 0.00170741f $X=-0.05 $Y=0 $X2=3.295 $Y2=2.22
cc_97 N_GND_M1017_b D 0.0155354f $X=-0.05 $Y=0 $X2=3.295 $Y2=2.22
cc_98 N_GND_M1017_b N_CK_c_941_n 0.0294225f $X=-0.05 $Y=0 $X2=6.735 $Y2=2.93
cc_99 N_GND_M1017_b N_CK_c_942_n 0.0432725f $X=-0.05 $Y=0 $X2=6.79 $Y2=2.6
cc_100 N_GND_M1017_b N_CK_c_943_n 0.0240652f $X=-0.05 $Y=0 $X2=3.655 $Y2=2.765
cc_101 N_GND_M1017_b N_CK_c_944_n 0.0254608f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.85
cc_102 N_GND_M1017_b N_CK_c_945_n 0.0173906f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.685
cc_103 N_GND_c_88_p N_CK_c_945_n 0.00606474f $X=4.685 $Y=0.152 $X2=4.135
+ $Y2=1.685
cc_104 N_GND_c_5_p N_CK_c_945_n 0.00468827f $X=9.855 $Y=0.19 $X2=4.135 $Y2=1.685
cc_105 N_GND_M1017_b N_CK_c_948_n 0.0252285f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.85
cc_106 N_GND_M1017_b N_CK_c_949_n 0.0175305f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.685
cc_107 N_GND_c_107_p N_CK_c_949_n 0.00606474f $X=6.435 $Y=0.152 $X2=5.405
+ $Y2=1.685
cc_108 N_GND_c_5_p N_CK_c_949_n 0.00468827f $X=9.855 $Y=0.19 $X2=5.405 $Y2=1.685
cc_109 N_GND_M1017_b N_CK_c_952_n 0.0230394f $X=-0.05 $Y=0 $X2=5.885 $Y2=2.765
cc_110 N_GND_M1017_b N_CK_c_953_n 0.0183851f $X=-0.05 $Y=0 $X2=6.762 $Y2=1.685
cc_111 N_GND_c_50_p N_CK_c_953_n 0.00356864f $X=6.52 $Y=0.825 $X2=6.762
+ $Y2=1.685
cc_112 N_GND_c_112_p N_CK_c_953_n 0.00606474f $X=7.385 $Y=0.152 $X2=6.762
+ $Y2=1.685
cc_113 N_GND_c_51_p N_CK_c_953_n 0.00462235f $X=7.47 $Y=0.825 $X2=6.762
+ $Y2=1.685
cc_114 N_GND_c_5_p N_CK_c_953_n 0.00468827f $X=9.855 $Y=0.19 $X2=6.762 $Y2=1.685
cc_115 N_GND_M1017_b N_CK_c_958_n 0.0130903f $X=-0.05 $Y=0 $X2=6.762 $Y2=1.835
cc_116 N_GND_M1017_b N_CK_c_959_n 0.00600607f $X=-0.05 $Y=0 $X2=4.05 $Y2=2.59
cc_117 N_GND_M1017_b N_CK_c_960_n 0.00921066f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.85
cc_118 N_GND_M1017_b N_CK_c_961_n 0.00838835f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.85
cc_119 N_GND_M1017_b N_CK_c_962_n 0.00543853f $X=-0.05 $Y=0 $X2=5.8 $Y2=2.59
cc_120 N_GND_M1017_b N_CK_c_963_n 5.00459e-19 $X=-0.05 $Y=0 $X2=5.49 $Y2=2.59
cc_121 N_GND_M1017_b N_CK_c_964_n 7.61111e-19 $X=-0.05 $Y=0 $X2=6.88 $Y2=2.59
cc_122 N_GND_M1017_b N_CK_c_965_n 0.00276905f $X=-0.05 $Y=0 $X2=3.655 $Y2=2.59
cc_123 N_GND_M1017_b N_CK_c_966_n 0.00265612f $X=-0.05 $Y=0 $X2=5.885 $Y2=2.59
cc_124 N_GND_M1017_b N_CK_c_967_n 0.0238264f $X=-0.05 $Y=0 $X2=5.74 $Y2=2.59
cc_125 N_GND_M1017_b N_CK_c_968_n 0.00704113f $X=-0.05 $Y=0 $X2=3.8 $Y2=2.59
cc_126 N_GND_M1017_b N_CK_c_969_n 0.00818551f $X=-0.05 $Y=0 $X2=6.735 $Y2=2.59
cc_127 N_GND_M1017_b N_CK_c_970_n 0.0038305f $X=-0.05 $Y=0 $X2=6.03 $Y2=2.59
cc_128 N_GND_M1017_b CK 0.00234237f $X=-0.05 $Y=0 $X2=6.88 $Y2=2.59
cc_129 N_GND_M1017_b N_A_217_617#_M1021_g 0.0171814f $X=-0.05 $Y=0 $X2=4.555
+ $Y2=1.075
cc_130 N_GND_c_88_p N_A_217_617#_M1021_g 0.00606474f $X=4.685 $Y=0.152 $X2=4.555
+ $Y2=1.075
cc_131 N_GND_c_49_p N_A_217_617#_M1021_g 0.00354579f $X=4.77 $Y=0.825 $X2=4.555
+ $Y2=1.075
cc_132 N_GND_c_5_p N_A_217_617#_M1021_g 0.00468827f $X=9.855 $Y=0.19 $X2=4.555
+ $Y2=1.075
cc_133 N_GND_M1017_b N_A_217_617#_c_1178_n 0.0240953f $X=-0.05 $Y=0 $X2=4.91
+ $Y2=1.85
cc_134 N_GND_c_49_p N_A_217_617#_c_1178_n 8.07204e-19 $X=4.77 $Y=0.825 $X2=4.91
+ $Y2=1.85
cc_135 N_GND_M1017_b N_A_217_617#_c_1180_n 0.0105855f $X=-0.05 $Y=0 $X2=4.63
+ $Y2=1.85
cc_136 N_GND_M1017_b N_A_217_617#_c_1181_n 0.023252f $X=-0.05 $Y=0 $X2=4.91
+ $Y2=2.765
cc_137 N_GND_M1017_b N_A_217_617#_c_1182_n 0.0103717f $X=-0.05 $Y=0 $X2=4.63
+ $Y2=2.765
cc_138 N_GND_M1017_b N_A_217_617#_M1026_g 0.0163216f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=1.075
cc_139 N_GND_c_49_p N_A_217_617#_M1026_g 0.00354579f $X=4.77 $Y=0.825 $X2=4.985
+ $Y2=1.075
cc_140 N_GND_c_107_p N_A_217_617#_M1026_g 0.00606474f $X=6.435 $Y=0.152
+ $X2=4.985 $Y2=1.075
cc_141 N_GND_c_5_p N_A_217_617#_M1026_g 0.00468827f $X=9.855 $Y=0.19 $X2=4.985
+ $Y2=1.075
cc_142 N_GND_M1017_b N_A_217_617#_c_1187_n 0.00601555f $X=-0.05 $Y=0 $X2=1.21
+ $Y2=3.795
cc_143 N_GND_M1017_b N_A_217_617#_c_1188_n 0.00760261f $X=-0.05 $Y=0 $X2=1.625
+ $Y2=2.02
cc_144 N_GND_M1017_b N_A_217_617#_c_1189_n 0.00184107f $X=-0.05 $Y=0 $X2=1.295
+ $Y2=2.02
cc_145 N_GND_M1017_b N_A_217_617#_c_1190_n 0.00648484f $X=-0.05 $Y=0 $X2=1.71
+ $Y2=0.825
cc_146 N_GND_c_14_p N_A_217_617#_c_1190_n 0.00736239f $X=2.415 $Y=0.152 $X2=1.71
+ $Y2=0.825
cc_147 N_GND_c_5_p N_A_217_617#_c_1190_n 0.00476261f $X=9.855 $Y=0.19 $X2=1.71
+ $Y2=0.825
cc_148 N_GND_M1017_b N_A_217_617#_c_1193_n 0.0087185f $X=-0.05 $Y=0 $X2=4.725
+ $Y2=2.765
cc_149 N_GND_M1017_b N_A_217_617#_c_1194_n 0.00245573f $X=-0.05 $Y=0 $X2=4.725
+ $Y2=1.85
cc_150 N_GND_c_49_p N_A_217_617#_c_1194_n 0.00177942f $X=4.77 $Y=0.825 $X2=4.725
+ $Y2=1.85
cc_151 N_GND_M1017_b N_A_217_617#_c_1196_n 0.0504449f $X=-0.05 $Y=0 $X2=4.49
+ $Y2=1.85
cc_152 N_GND_M1017_b N_A_217_617#_c_1197_n 0.00355505f $X=-0.05 $Y=0 $X2=1.855
+ $Y2=1.85
cc_153 N_GND_M1017_b N_A_704_89#_c_1338_n 0.0173059f $X=-0.05 $Y=0 $X2=3.595
+ $Y2=1.685
cc_154 N_GND_c_88_p N_A_704_89#_c_1338_n 0.00606474f $X=4.685 $Y=0.152 $X2=3.595
+ $Y2=1.685
cc_155 N_GND_c_5_p N_A_704_89#_c_1338_n 0.00468827f $X=9.855 $Y=0.19 $X2=3.595
+ $Y2=1.685
cc_156 N_GND_M1017_b N_A_704_89#_c_1341_n 0.0203057f $X=-0.05 $Y=0 $X2=3.715
+ $Y2=2.225
cc_157 N_GND_M1017_b N_A_704_89#_c_1342_n 0.0187566f $X=-0.05 $Y=0 $X2=4.12
+ $Y2=2.3
cc_158 N_GND_M1017_b N_A_704_89#_c_1343_n 0.00755029f $X=-0.05 $Y=0 $X2=3.79
+ $Y2=2.3
cc_159 N_GND_M1017_b N_A_704_89#_M1031_g 0.0321382f $X=-0.05 $Y=0 $X2=4.195
+ $Y2=4.585
cc_160 N_GND_M1017_b N_A_704_89#_c_1345_n 0.0559794f $X=-0.05 $Y=0 $X2=5.27
+ $Y2=2.3
cc_161 N_GND_M1017_b N_A_704_89#_M1025_g 0.0316517f $X=-0.05 $Y=0 $X2=5.345
+ $Y2=4.585
cc_162 N_GND_M1017_b N_A_704_89#_c_1347_n 0.0270462f $X=-0.05 $Y=0 $X2=5.75
+ $Y2=2.3
cc_163 N_GND_M1017_b N_A_704_89#_c_1348_n 0.0125754f $X=-0.05 $Y=0 $X2=5.825
+ $Y2=2.225
cc_164 N_GND_M1017_b N_A_704_89#_c_1349_n 0.0141451f $X=-0.05 $Y=0 $X2=3.715
+ $Y2=1.76
cc_165 N_GND_M1017_b N_A_704_89#_c_1350_n 0.00426512f $X=-0.05 $Y=0 $X2=4.195
+ $Y2=2.3
cc_166 N_GND_M1017_b N_A_704_89#_c_1351_n 0.00426512f $X=-0.05 $Y=0 $X2=5.345
+ $Y2=2.3
cc_167 N_GND_M1017_b N_A_704_89#_c_1352_n 0.0256431f $X=-0.05 $Y=0 $X2=5.885
+ $Y2=1.85
cc_168 N_GND_M1017_b N_A_704_89#_c_1353_n 0.01755f $X=-0.05 $Y=0 $X2=5.885
+ $Y2=1.685
cc_169 N_GND_c_107_p N_A_704_89#_c_1353_n 0.00606474f $X=6.435 $Y=0.152
+ $X2=5.885 $Y2=1.685
cc_170 N_GND_c_5_p N_A_704_89#_c_1353_n 0.00468827f $X=9.855 $Y=0.19 $X2=5.885
+ $Y2=1.685
cc_171 N_GND_M1017_b N_A_704_89#_c_1356_n 0.0116005f $X=-0.05 $Y=0 $X2=6.865
+ $Y2=1.85
cc_172 N_GND_c_50_p N_A_704_89#_c_1356_n 0.00564434f $X=6.52 $Y=0.825 $X2=6.865
+ $Y2=1.85
cc_173 N_GND_M1017_b N_A_704_89#_c_1358_n 0.00557295f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=0.825
cc_174 N_GND_c_50_p N_A_704_89#_c_1358_n 4.65312e-19 $X=6.52 $Y=0.825 $X2=6.95
+ $Y2=0.825
cc_175 N_GND_c_112_p N_A_704_89#_c_1358_n 0.0074445f $X=7.385 $Y=0.152 $X2=6.95
+ $Y2=0.825
cc_176 N_GND_c_51_p N_A_704_89#_c_1358_n 0.0356656f $X=7.47 $Y=0.825 $X2=6.95
+ $Y2=0.825
cc_177 N_GND_c_5_p N_A_704_89#_c_1358_n 0.00476261f $X=9.855 $Y=0.19 $X2=6.95
+ $Y2=0.825
cc_178 N_GND_M1017_b N_A_704_89#_c_1363_n 0.00299027f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=2.105
cc_179 N_GND_M1017_b N_A_704_89#_c_1364_n 0.011861f $X=-0.05 $Y=0 $X2=7.22
+ $Y2=3.1
cc_180 N_GND_M1017_b N_A_704_89#_c_1365_n 0.001308f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=1.85
cc_181 N_GND_M1017_b N_A_704_89#_c_1366_n 0.00945336f $X=-0.05 $Y=0 $X2=7.22
+ $Y2=2.19
cc_182 N_GND_M1017_b N_A_1246_89#_M1006_g 0.0319752f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=1.075
cc_183 N_GND_c_107_p N_A_1246_89#_M1006_g 0.00606474f $X=6.435 $Y=0.152
+ $X2=6.305 $Y2=1.075
cc_184 N_GND_c_50_p N_A_1246_89#_M1006_g 0.00360474f $X=6.52 $Y=0.825 $X2=6.305
+ $Y2=1.075
cc_185 N_GND_c_5_p N_A_1246_89#_M1006_g 0.00468827f $X=9.855 $Y=0.19 $X2=6.305
+ $Y2=1.075
cc_186 N_GND_M1017_b N_A_1246_89#_M1009_g 0.0327124f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=4.585
cc_187 N_GND_M1017_b N_A_1246_89#_M1007_g 0.0315215f $X=-0.05 $Y=0 $X2=9.495
+ $Y2=0.945
cc_188 N_GND_c_18_p N_A_1246_89#_M1007_g 0.00392369f $X=8.75 $Y=0.825 $X2=9.495
+ $Y2=0.945
cc_189 N_GND_c_189_p N_A_1246_89#_M1007_g 0.00606474f $X=9.625 $Y=0.152
+ $X2=9.495 $Y2=0.945
cc_190 N_GND_c_190_p N_A_1246_89#_M1007_g 0.00354579f $X=9.71 $Y=0.825 $X2=9.495
+ $Y2=0.945
cc_191 N_GND_c_5_p N_A_1246_89#_M1007_g 0.00468827f $X=9.855 $Y=0.19 $X2=9.495
+ $Y2=0.945
cc_192 N_GND_M1017_b N_A_1246_89#_c_1539_n 0.0263478f $X=-0.05 $Y=0 $X2=6.365
+ $Y2=2.19
cc_193 N_GND_M1017_b N_A_1246_89#_c_1540_n 0.0270403f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=2.19
cc_194 N_GND_M1017_b N_A_1246_89#_c_1541_n 0.0124759f $X=-0.05 $Y=0 $X2=9.382
+ $Y2=2.025
cc_195 N_GND_M1017_b N_A_1246_89#_c_1542_n 0.0133302f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=1.8
cc_196 N_GND_M1017_b N_A_1246_89#_c_1543_n 0.0282913f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=2.855
cc_197 N_GND_M1017_b N_A_1246_89#_c_1544_n 0.00443937f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=3.005
cc_198 N_GND_M1017_b N_A_1246_89#_c_1545_n 0.0039674f $X=-0.05 $Y=0 $X2=6.365
+ $Y2=2.19
cc_199 N_GND_M1017_b N_A_1246_89#_c_1546_n 0.00796703f $X=-0.05 $Y=0 $X2=8.26
+ $Y2=0.825
cc_200 N_GND_c_17_p N_A_1246_89#_c_1546_n 0.00750865f $X=8.665 $Y=0.152 $X2=8.26
+ $Y2=0.825
cc_201 N_GND_c_5_p N_A_1246_89#_c_1546_n 0.00476261f $X=9.855 $Y=0.19 $X2=8.26
+ $Y2=0.825
cc_202 N_GND_M1017_b N_A_1246_89#_c_1549_n 0.00551501f $X=-0.05 $Y=0 $X2=8.76
+ $Y2=3.795
cc_203 N_GND_M1017_b N_A_1246_89#_c_1550_n 0.0207701f $X=-0.05 $Y=0 $X2=8.845
+ $Y2=2.19
cc_204 N_GND_M1017_b N_A_1246_89#_c_1551_n 0.00950815f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=2.19
cc_205 N_GND_M1017_b N_A_1246_89#_c_1552_n 0.0568381f $X=-0.05 $Y=0 $X2=9.235
+ $Y2=2.19
cc_206 N_GND_M1017_b N_A_1246_89#_c_1553_n 0.00189525f $X=-0.05 $Y=0 $X2=6.51
+ $Y2=2.19
cc_207 N_GND_M1017_b N_A_1246_89#_c_1554_n 0.0014645f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=2.19
cc_208 N_GND_M1017_b N_A_1084_115#_c_1705_n 0.0450481f $X=-0.05 $Y=0 $X2=7.505
+ $Y2=2.63
cc_209 N_GND_M1017_b N_A_1084_115#_c_1706_n 0.0178887f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.69
cc_210 N_GND_c_51_p N_A_1084_115#_c_1706_n 0.00715019f $X=7.47 $Y=0.825
+ $X2=7.685 $Y2=1.69
cc_211 N_GND_c_17_p N_A_1084_115#_c_1706_n 0.00606474f $X=8.665 $Y=0.152
+ $X2=7.685 $Y2=1.69
cc_212 N_GND_c_5_p N_A_1084_115#_c_1706_n 0.00468827f $X=9.855 $Y=0.19 $X2=7.685
+ $Y2=1.69
cc_213 N_GND_M1017_b N_A_1084_115#_c_1710_n 0.0235095f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.77
cc_214 N_GND_c_51_p N_A_1084_115#_c_1710_n 0.00391038f $X=7.47 $Y=0.825
+ $X2=7.685 $Y2=1.77
cc_215 N_GND_M1017_b N_A_1084_115#_c_1712_n 0.0324837f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=2.765
cc_216 N_GND_M1017_b N_A_1084_115#_c_1713_n 0.011286f $X=-0.05 $Y=0 $X2=5.065
+ $Y2=1.85
cc_217 N_GND_M1017_b N_A_1084_115#_c_1714_n 0.00313975f $X=-0.05 $Y=0 $X2=5.645
+ $Y2=0.825
cc_218 N_GND_c_107_p N_A_1084_115#_c_1714_n 0.0149333f $X=6.435 $Y=0.152
+ $X2=5.645 $Y2=0.825
cc_219 N_GND_c_5_p N_A_1084_115#_c_1714_n 0.00958198f $X=9.855 $Y=0.19 $X2=5.645
+ $Y2=0.825
cc_220 N_GND_M1017_b N_A_1084_115#_c_1717_n 0.00582616f $X=-0.05 $Y=0 $X2=7.595
+ $Y2=1.85
cc_221 N_GND_c_51_p N_A_1084_115#_c_1717_n 0.00131024f $X=7.47 $Y=0.825
+ $X2=7.595 $Y2=1.85
cc_222 N_GND_M1017_b N_A_1084_115#_c_1719_n 0.022645f $X=-0.05 $Y=0 $X2=7.45
+ $Y2=1.85
cc_223 N_GND_c_50_p N_A_1084_115#_c_1719_n 5.03331e-19 $X=6.52 $Y=0.825 $X2=7.45
+ $Y2=1.85
cc_224 N_GND_c_51_p N_A_1084_115#_c_1719_n 3.1624e-19 $X=7.47 $Y=0.825 $X2=7.45
+ $Y2=1.85
cc_225 N_GND_M1017_b N_A_1084_115#_c_1722_n 0.00120467f $X=-0.05 $Y=0 $X2=5.21
+ $Y2=1.85
cc_226 N_GND_M1017_b N_A_1084_115#_c_1723_n 0.00169121f $X=-0.05 $Y=0 $X2=7.595
+ $Y2=1.85
cc_227 N_GND_c_51_p N_A_1084_115#_c_1723_n 4.00959e-19 $X=7.47 $Y=0.825
+ $X2=7.595 $Y2=1.85
cc_228 N_GND_M1017_b N_QN_M1010_g 0.0707753f $X=-0.05 $Y=0 $X2=9.925 $Y2=0.945
cc_229 N_GND_c_190_p N_QN_M1010_g 0.00354579f $X=9.71 $Y=0.825 $X2=9.925
+ $Y2=0.945
cc_230 N_GND_c_5_p N_QN_M1010_g 0.00468827f $X=9.855 $Y=0.19 $X2=9.925 $Y2=0.945
cc_231 N_GND_M1017_b N_QN_M1029_g 0.0186095f $X=-0.05 $Y=0 $X2=9.925 $Y2=5.085
cc_232 N_GND_M1017_b N_QN_c_1866_n 0.0291912f $X=-0.05 $Y=0 $X2=9.865 $Y2=2.395
cc_233 N_GND_M1017_b N_QN_c_1867_n 0.0105985f $X=-0.05 $Y=0 $X2=9.28 $Y2=0.825
cc_234 N_GND_c_18_p N_QN_c_1867_n 0.0209197f $X=8.75 $Y=0.825 $X2=9.28 $Y2=0.825
cc_235 N_GND_c_189_p N_QN_c_1867_n 0.00736239f $X=9.625 $Y=0.152 $X2=9.28
+ $Y2=0.825
cc_236 N_GND_c_5_p N_QN_c_1867_n 0.00476261f $X=9.855 $Y=0.19 $X2=9.28 $Y2=0.825
cc_237 N_GND_M1017_b N_QN_c_1871_n 0.00102655f $X=-0.05 $Y=0 $X2=9.28 $Y2=2.96
cc_238 N_GND_M1017_b N_QN_c_1872_n 0.0171269f $X=-0.05 $Y=0 $X2=9.78 $Y2=1.85
cc_239 N_GND_M1017_b N_QN_c_1873_n 0.00294844f $X=-0.05 $Y=0 $X2=9.365 $Y2=1.85
cc_240 N_GND_M1017_b N_QN_c_1874_n 0.0176115f $X=-0.05 $Y=0 $X2=9.78 $Y2=2.765
cc_241 N_GND_M1017_b N_QN_c_1875_n 0.00297015f $X=-0.05 $Y=0 $X2=9.365 $Y2=2.765
cc_242 N_GND_M1017_b N_QN_c_1876_n 0.0034889f $X=-0.05 $Y=0 $X2=9.865 $Y2=2.395
cc_243 N_GND_M1017_b QN 0.00258296f $X=-0.05 $Y=0 $X2=9.285 $Y2=2.96
cc_244 N_GND_M1017_b N_Q_c_1989_n 0.0153135f $X=-0.05 $Y=0 $X2=10.14 $Y2=0.825
cc_245 N_GND_c_5_p N_Q_c_1989_n 0.00476261f $X=9.855 $Y=0.19 $X2=10.14 $Y2=0.825
cc_246 N_GND_M1017_b N_Q_c_1991_n 0.0625704f $X=-0.05 $Y=0 $X2=10.255 $Y2=3.16
cc_247 N_GND_M1017_b N_Q_c_1992_n 0.0184431f $X=-0.05 $Y=0 $X2=10.255 $Y2=1.515
cc_248 N_VDD_M1019_b N_RN_M1019_g 0.0266406f $X=-0.05 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_249 N_VDD_c_249_p N_RN_M1019_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_250 N_VDD_c_250_p N_RN_M1019_g 0.00606474f $X=1.985 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_251 N_VDD_c_251_p N_RN_M1019_g 0.00468827f $X=9.855 $Y=6.47 $X2=0.475
+ $Y2=4.585
cc_252 N_VDD_M1019_s N_RN_c_399_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32
+ $Y2=3.33
cc_253 N_VDD_M1019_b N_RN_c_399_n 0.00618364f $X=-0.05 $Y=2.905 $X2=0.32
+ $Y2=3.33
cc_254 N_VDD_c_249_p N_RN_c_399_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_255 N_VDD_M1019_s RN 0.0162774f $X=0.135 $Y=3.085 $X2=0.325 $Y2=3.33
cc_256 N_VDD_c_249_p RN 0.00522047f $X=0.26 $Y=4.135 $X2=0.325 $Y2=3.33
cc_257 N_VDD_M1019_b N_A_110_115#_M1016_g 0.0246426f $X=-0.05 $Y=2.905 $X2=1.425
+ $Y2=4.585
cc_258 N_VDD_c_250_p N_A_110_115#_M1016_g 0.00606474f $X=1.985 $Y=6.507
+ $X2=1.425 $Y2=4.585
cc_259 N_VDD_c_251_p N_A_110_115#_M1016_g 0.00468827f $X=9.855 $Y=6.47 $X2=1.425
+ $Y2=4.585
cc_260 N_VDD_M1019_b N_A_110_115#_M1004_g 0.0246768f $X=-0.05 $Y=2.905 $X2=8.545
+ $Y2=4.585
cc_261 N_VDD_c_261_p N_A_110_115#_M1004_g 0.00606474f $X=9.625 $Y=6.507
+ $X2=8.545 $Y2=4.585
cc_262 N_VDD_c_251_p N_A_110_115#_M1004_g 0.00468827f $X=9.855 $Y=6.47 $X2=8.545
+ $Y2=4.585
cc_263 N_VDD_M1019_b N_A_110_115#_c_454_n 0.00549797f $X=-0.05 $Y=2.905 $X2=0.69
+ $Y2=3.455
cc_264 N_VDD_c_250_p N_A_110_115#_c_454_n 0.00757793f $X=1.985 $Y=6.507 $X2=0.69
+ $Y2=3.455
cc_265 N_VDD_c_251_p N_A_110_115#_c_454_n 0.00476261f $X=9.855 $Y=6.47 $X2=0.69
+ $Y2=3.455
cc_266 N_VDD_M1019_b N_SN_M1000_g 0.0188578f $X=-0.05 $Y=2.905 $X2=1.855
+ $Y2=4.585
cc_267 N_VDD_c_250_p N_SN_M1000_g 0.00606474f $X=1.985 $Y=6.507 $X2=1.855
+ $Y2=4.585
cc_268 N_VDD_c_268_p N_SN_M1000_g 0.00354579f $X=2.07 $Y=4.135 $X2=1.855
+ $Y2=4.585
cc_269 N_VDD_c_251_p N_SN_M1000_g 0.00468827f $X=9.855 $Y=6.47 $X2=1.855
+ $Y2=4.585
cc_270 N_VDD_M1019_b N_SN_M1035_g 0.019722f $X=-0.05 $Y=2.905 $X2=8.115
+ $Y2=4.585
cc_271 N_VDD_c_271_p N_SN_M1035_g 0.00354579f $X=7.9 $Y=4.135 $X2=8.115
+ $Y2=4.585
cc_272 N_VDD_c_261_p N_SN_M1035_g 0.00606474f $X=9.625 $Y=6.507 $X2=8.115
+ $Y2=4.585
cc_273 N_VDD_c_251_p N_SN_M1035_g 0.00468827f $X=9.855 $Y=6.47 $X2=8.115
+ $Y2=4.585
cc_274 N_VDD_M1019_b N_SN_c_653_n 0.00205457f $X=-0.05 $Y=2.905 $X2=1.71
+ $Y2=2.96
cc_275 N_VDD_M1019_b N_SN_c_654_n 0.00449283f $X=-0.05 $Y=2.905 $X2=7.935
+ $Y2=2.96
cc_276 N_VDD_M1019_b N_SN_c_657_n 0.0566252f $X=-0.05 $Y=2.905 $X2=7.79 $Y2=2.96
cc_277 N_VDD_c_277_p N_SN_c_657_n 0.00464215f $X=4.77 $Y=3.795 $X2=7.79 $Y2=2.96
cc_278 N_VDD_c_278_p N_SN_c_657_n 0.0090257f $X=6.52 $Y=3.455 $X2=7.79 $Y2=2.96
cc_279 N_VDD_M1019_b N_SN_c_658_n 0.00372061f $X=-0.05 $Y=2.905 $X2=1.855
+ $Y2=2.96
cc_280 N_VDD_M1019_b SN 0.00292685f $X=-0.05 $Y=2.905 $X2=7.935 $Y2=2.96
cc_281 N_VDD_M1019_b N_A_432_520#_M1003_g 0.0213832f $X=-0.05 $Y=2.905 $X2=2.285
+ $Y2=4.585
cc_282 N_VDD_c_268_p N_A_432_520#_M1003_g 0.00354579f $X=2.07 $Y=4.135 $X2=2.285
+ $Y2=4.585
cc_283 N_VDD_c_283_p N_A_432_520#_M1003_g 0.00606474f $X=2.935 $Y=6.507
+ $X2=2.285 $Y2=4.585
cc_284 N_VDD_c_284_p N_A_432_520#_M1003_g 0.00822619f $X=3.02 $Y=3.795 $X2=2.285
+ $Y2=4.585
cc_285 N_VDD_c_251_p N_A_432_520#_M1003_g 0.00468827f $X=9.855 $Y=6.47 $X2=2.285
+ $Y2=4.585
cc_286 N_VDD_M1019_b N_A_432_520#_c_816_n 0.0057899f $X=-0.05 $Y=2.905 $X2=2.295
+ $Y2=2.765
cc_287 N_VDD_M1019_b N_A_432_520#_c_817_n 0.00281226f $X=-0.05 $Y=2.905
+ $X2=2.295 $Y2=2.765
cc_288 N_VDD_M1008_s N_A_432_520#_c_833_n 0.00705065f $X=2.895 $Y=3.085
+ $X2=3.725 $Y2=3.185
cc_289 N_VDD_M1019_b N_A_432_520#_c_833_n 0.013691f $X=-0.05 $Y=2.905 $X2=3.725
+ $Y2=3.185
cc_290 N_VDD_c_284_p N_A_432_520#_c_833_n 0.00850976f $X=3.02 $Y=3.795 $X2=3.725
+ $Y2=3.185
cc_291 N_VDD_M1019_b N_A_432_520#_c_836_n 0.00313975f $X=-0.05 $Y=2.905
+ $X2=3.895 $Y2=3.455
cc_292 N_VDD_c_292_p N_A_432_520#_c_836_n 0.0149718f $X=4.685 $Y=6.507 $X2=3.895
+ $Y2=3.455
cc_293 N_VDD_c_251_p N_A_432_520#_c_836_n 0.00958198f $X=9.855 $Y=6.47 $X2=3.895
+ $Y2=3.455
cc_294 N_VDD_M1019_b N_D_M1008_g 0.0224773f $X=-0.05 $Y=2.905 $X2=3.235
+ $Y2=4.585
cc_295 N_VDD_c_284_p N_D_M1008_g 0.00713292f $X=3.02 $Y=3.795 $X2=3.235
+ $Y2=4.585
cc_296 N_VDD_c_292_p N_D_M1008_g 0.00606474f $X=4.685 $Y=6.507 $X2=3.235
+ $Y2=4.585
cc_297 N_VDD_c_251_p N_D_M1008_g 0.00468827f $X=9.855 $Y=6.47 $X2=3.235
+ $Y2=4.585
cc_298 N_VDD_M1019_b N_CK_M1034_g 0.0188823f $X=-0.05 $Y=2.905 $X2=3.595
+ $Y2=4.585
cc_299 N_VDD_c_292_p N_CK_M1034_g 0.00606474f $X=4.685 $Y=6.507 $X2=3.595
+ $Y2=4.585
cc_300 N_VDD_c_251_p N_CK_M1034_g 0.00468827f $X=9.855 $Y=6.47 $X2=3.595
+ $Y2=4.585
cc_301 N_VDD_M1019_b N_CK_M1020_g 0.0188823f $X=-0.05 $Y=2.905 $X2=5.945
+ $Y2=4.585
cc_302 N_VDD_c_302_p N_CK_M1020_g 0.00606474f $X=6.435 $Y=6.507 $X2=5.945
+ $Y2=4.585
cc_303 N_VDD_c_251_p N_CK_M1020_g 0.00468827f $X=9.855 $Y=6.47 $X2=5.945
+ $Y2=4.585
cc_304 N_VDD_M1019_b N_CK_c_941_n 0.007968f $X=-0.05 $Y=2.905 $X2=6.735 $Y2=2.93
cc_305 N_VDD_M1019_b N_CK_M1012_g 0.0241401f $X=-0.05 $Y=2.905 $X2=6.735
+ $Y2=4.585
cc_306 N_VDD_c_278_p N_CK_M1012_g 0.00354579f $X=6.52 $Y=3.455 $X2=6.735
+ $Y2=4.585
cc_307 N_VDD_c_307_p N_CK_M1012_g 0.00606474f $X=7.815 $Y=6.507 $X2=6.735
+ $Y2=4.585
cc_308 N_VDD_c_251_p N_CK_M1012_g 0.00468827f $X=9.855 $Y=6.47 $X2=6.735
+ $Y2=4.585
cc_309 N_VDD_M1019_b N_CK_c_943_n 0.00508175f $X=-0.05 $Y=2.905 $X2=3.655
+ $Y2=2.765
cc_310 N_VDD_M1019_b N_CK_c_952_n 0.00508175f $X=-0.05 $Y=2.905 $X2=5.885
+ $Y2=2.765
cc_311 N_VDD_M1019_b N_CK_c_964_n 0.0010436f $X=-0.05 $Y=2.905 $X2=6.88 $Y2=2.59
cc_312 N_VDD_M1019_b N_CK_c_965_n 2.35021e-19 $X=-0.05 $Y=2.905 $X2=3.655
+ $Y2=2.59
cc_313 N_VDD_M1019_b N_CK_c_966_n 7.56914e-19 $X=-0.05 $Y=2.905 $X2=5.885
+ $Y2=2.59
cc_314 N_VDD_M1019_b N_A_217_617#_M1024_g 0.0179013f $X=-0.05 $Y=2.905 $X2=4.555
+ $Y2=4.585
cc_315 N_VDD_c_292_p N_A_217_617#_M1024_g 0.00606474f $X=4.685 $Y=6.507
+ $X2=4.555 $Y2=4.585
cc_316 N_VDD_c_277_p N_A_217_617#_M1024_g 0.00354579f $X=4.77 $Y=3.795 $X2=4.555
+ $Y2=4.585
cc_317 N_VDD_c_251_p N_A_217_617#_M1024_g 0.00468827f $X=9.855 $Y=6.47 $X2=4.555
+ $Y2=4.585
cc_318 N_VDD_c_277_p N_A_217_617#_c_1181_n 7.6376e-19 $X=4.77 $Y=3.795 $X2=4.91
+ $Y2=2.765
cc_319 N_VDD_M1019_b N_A_217_617#_M1027_g 0.0175507f $X=-0.05 $Y=2.905 $X2=4.985
+ $Y2=4.585
cc_320 N_VDD_c_277_p N_A_217_617#_M1027_g 0.00354579f $X=4.77 $Y=3.795 $X2=4.985
+ $Y2=4.585
cc_321 N_VDD_c_302_p N_A_217_617#_M1027_g 0.00606474f $X=6.435 $Y=6.507
+ $X2=4.985 $Y2=4.585
cc_322 N_VDD_c_251_p N_A_217_617#_M1027_g 0.00468827f $X=9.855 $Y=6.47 $X2=4.985
+ $Y2=4.585
cc_323 N_VDD_M1019_b N_A_217_617#_c_1187_n 0.00436897f $X=-0.05 $Y=2.905
+ $X2=1.21 $Y2=3.795
cc_324 N_VDD_c_250_p N_A_217_617#_c_1187_n 0.00745733f $X=1.985 $Y=6.507
+ $X2=1.21 $Y2=3.795
cc_325 N_VDD_c_251_p N_A_217_617#_c_1187_n 0.00476261f $X=9.855 $Y=6.47 $X2=1.21
+ $Y2=3.795
cc_326 N_VDD_M1019_b N_A_217_617#_c_1193_n 0.00208967f $X=-0.05 $Y=2.905
+ $X2=4.725 $Y2=2.765
cc_327 N_VDD_c_277_p N_A_217_617#_c_1193_n 0.00215846f $X=4.77 $Y=3.795
+ $X2=4.725 $Y2=2.765
cc_328 N_VDD_M1019_b N_A_704_89#_M1031_g 0.0199908f $X=-0.05 $Y=2.905 $X2=4.195
+ $Y2=4.585
cc_329 N_VDD_c_292_p N_A_704_89#_M1031_g 0.00606474f $X=4.685 $Y=6.507 $X2=4.195
+ $Y2=4.585
cc_330 N_VDD_c_251_p N_A_704_89#_M1031_g 0.00468827f $X=9.855 $Y=6.47 $X2=4.195
+ $Y2=4.585
cc_331 N_VDD_M1019_b N_A_704_89#_M1025_g 0.0199837f $X=-0.05 $Y=2.905 $X2=5.345
+ $Y2=4.585
cc_332 N_VDD_c_302_p N_A_704_89#_M1025_g 0.00606474f $X=6.435 $Y=6.507 $X2=5.345
+ $Y2=4.585
cc_333 N_VDD_c_251_p N_A_704_89#_M1025_g 0.00468827f $X=9.855 $Y=6.47 $X2=5.345
+ $Y2=4.585
cc_334 N_VDD_M1019_b N_A_704_89#_c_1373_n 0.00156053f $X=-0.05 $Y=2.905 $X2=6.95
+ $Y2=3.455
cc_335 N_VDD_c_307_p N_A_704_89#_c_1373_n 0.0074445f $X=7.815 $Y=6.507 $X2=6.95
+ $Y2=3.455
cc_336 N_VDD_c_251_p N_A_704_89#_c_1373_n 0.00476261f $X=9.855 $Y=6.47 $X2=6.95
+ $Y2=3.455
cc_337 N_VDD_M1019_b N_A_704_89#_c_1364_n 0.00526199f $X=-0.05 $Y=2.905 $X2=7.22
+ $Y2=3.1
cc_338 N_VDD_M1019_b N_A_704_89#_c_1377_n 0.012303f $X=-0.05 $Y=2.905 $X2=7.22
+ $Y2=3.185
cc_339 N_VDD_M1019_b N_A_1246_89#_M1009_g 0.0182476f $X=-0.05 $Y=2.905 $X2=6.305
+ $Y2=4.585
cc_340 N_VDD_c_302_p N_A_1246_89#_M1009_g 0.00606474f $X=6.435 $Y=6.507
+ $X2=6.305 $Y2=4.585
cc_341 N_VDD_c_278_p N_A_1246_89#_M1009_g 0.00354579f $X=6.52 $Y=3.455 $X2=6.305
+ $Y2=4.585
cc_342 N_VDD_c_251_p N_A_1246_89#_M1009_g 0.00468827f $X=9.855 $Y=6.47 $X2=6.305
+ $Y2=4.585
cc_343 N_VDD_M1019_b N_A_1246_89#_M1028_g 0.0761326f $X=-0.05 $Y=2.905 $X2=9.495
+ $Y2=5.085
cc_344 N_VDD_c_261_p N_A_1246_89#_M1028_g 0.00606474f $X=9.625 $Y=6.507
+ $X2=9.495 $Y2=5.085
cc_345 N_VDD_c_345_p N_A_1246_89#_M1028_g 0.00354579f $X=9.71 $Y=4.475 $X2=9.495
+ $Y2=5.085
cc_346 N_VDD_c_251_p N_A_1246_89#_M1028_g 0.00468827f $X=9.855 $Y=6.47 $X2=9.495
+ $Y2=5.085
cc_347 N_VDD_M1019_b N_A_1246_89#_c_1544_n 0.00913729f $X=-0.05 $Y=2.905
+ $X2=9.47 $Y2=3.005
cc_348 N_VDD_M1019_b N_A_1246_89#_c_1549_n 0.00440545f $X=-0.05 $Y=2.905
+ $X2=8.76 $Y2=3.795
cc_349 N_VDD_c_261_p N_A_1246_89#_c_1549_n 0.00754714f $X=9.625 $Y=6.507
+ $X2=8.76 $Y2=3.795
cc_350 N_VDD_c_251_p N_A_1246_89#_c_1549_n 0.00476261f $X=9.855 $Y=6.47 $X2=8.76
+ $Y2=3.795
cc_351 N_VDD_M1019_b N_A_1084_115#_M1014_g 0.0254863f $X=-0.05 $Y=2.905
+ $X2=7.685 $Y2=4.585
cc_352 N_VDD_c_307_p N_A_1084_115#_M1014_g 0.00606474f $X=7.815 $Y=6.507
+ $X2=7.685 $Y2=4.585
cc_353 N_VDD_c_271_p N_A_1084_115#_M1014_g 0.00354579f $X=7.9 $Y=4.135 $X2=7.685
+ $Y2=4.585
cc_354 N_VDD_c_251_p N_A_1084_115#_M1014_g 0.00468827f $X=9.855 $Y=6.47
+ $X2=7.685 $Y2=4.585
cc_355 N_VDD_M1019_b N_A_1084_115#_c_1713_n 0.00207418f $X=-0.05 $Y=2.905
+ $X2=5.065 $Y2=1.85
cc_356 N_VDD_M1019_b N_A_1084_115#_c_1730_n 0.00313975f $X=-0.05 $Y=2.905
+ $X2=5.645 $Y2=3.795
cc_357 N_VDD_c_302_p N_A_1084_115#_c_1730_n 0.0149333f $X=6.435 $Y=6.507
+ $X2=5.645 $Y2=3.795
cc_358 N_VDD_c_251_p N_A_1084_115#_c_1730_n 0.00958198f $X=9.855 $Y=6.47
+ $X2=5.645 $Y2=3.795
cc_359 N_VDD_M1019_b N_A_1084_115#_c_1717_n 9.87966e-19 $X=-0.05 $Y=2.905
+ $X2=7.595 $Y2=1.85
cc_360 N_VDD_M1019_b N_QN_M1029_g 0.0840918f $X=-0.05 $Y=2.905 $X2=9.925
+ $Y2=5.085
cc_361 N_VDD_c_345_p N_QN_M1029_g 0.00354579f $X=9.71 $Y=4.475 $X2=9.925
+ $Y2=5.085
cc_362 N_VDD_c_362_p N_QN_M1029_g 0.00606474f $X=9.855 $Y=6.44 $X2=9.925
+ $Y2=5.085
cc_363 N_VDD_c_251_p N_QN_M1029_g 0.00468827f $X=9.855 $Y=6.47 $X2=9.925
+ $Y2=5.085
cc_364 N_VDD_M1019_b N_QN_c_1871_n 0.029401f $X=-0.05 $Y=2.905 $X2=9.28 $Y2=2.96
cc_365 N_VDD_c_261_p N_QN_c_1871_n 0.00736239f $X=9.625 $Y=6.507 $X2=9.28
+ $Y2=2.96
cc_366 N_VDD_c_251_p N_QN_c_1871_n 0.00476261f $X=9.855 $Y=6.47 $X2=9.28
+ $Y2=2.96
cc_367 N_VDD_M1019_b QN 0.0101088f $X=-0.05 $Y=2.905 $X2=9.285 $Y2=2.96
cc_368 N_VDD_M1019_b N_A_300_617#_c_1946_n 0.00155118f $X=-0.05 $Y=2.905
+ $X2=1.64 $Y2=3.795
cc_369 N_VDD_c_250_p N_A_300_617#_c_1946_n 0.00734006f $X=1.985 $Y=6.507
+ $X2=1.64 $Y2=3.795
cc_370 N_VDD_c_251_p N_A_300_617#_c_1946_n 0.00475776f $X=9.855 $Y=6.47 $X2=1.64
+ $Y2=3.795
cc_371 N_VDD_M1000_d N_A_300_617#_c_1949_n 0.00482635f $X=1.93 $Y=3.085
+ $X2=2.415 $Y2=3.63
cc_372 N_VDD_c_268_p N_A_300_617#_c_1949_n 0.0135055f $X=2.07 $Y=4.135 $X2=2.415
+ $Y2=3.63
cc_373 N_VDD_c_284_p N_A_300_617#_c_1949_n 0.00811594f $X=3.02 $Y=3.795
+ $X2=2.415 $Y2=3.63
cc_374 N_VDD_M1019_b N_A_300_617#_c_1952_n 0.00156053f $X=-0.05 $Y=2.905 $X2=2.5
+ $Y2=3.795
cc_375 N_VDD_c_283_p N_A_300_617#_c_1952_n 0.00736752f $X=2.935 $Y=6.507 $X2=2.5
+ $Y2=3.795
cc_376 N_VDD_c_284_p N_A_300_617#_c_1952_n 0.101221f $X=3.02 $Y=3.795 $X2=2.5
+ $Y2=3.795
cc_377 N_VDD_c_251_p N_A_300_617#_c_1952_n 0.00476261f $X=9.855 $Y=6.47 $X2=2.5
+ $Y2=3.795
cc_378 N_VDD_M1019_b N_A_1469_617#_c_1970_n 0.00156053f $X=-0.05 $Y=2.905
+ $X2=7.47 $Y2=3.795
cc_379 N_VDD_c_307_p N_A_1469_617#_c_1970_n 0.00757793f $X=7.815 $Y=6.507
+ $X2=7.47 $Y2=3.795
cc_380 N_VDD_c_251_p N_A_1469_617#_c_1970_n 0.00476261f $X=9.855 $Y=6.47
+ $X2=7.47 $Y2=3.795
cc_381 N_VDD_M1014_d N_A_1469_617#_c_1973_n 0.00462014f $X=7.76 $Y=3.085
+ $X2=8.245 $Y2=3.63
cc_382 N_VDD_c_271_p N_A_1469_617#_c_1973_n 0.0135055f $X=7.9 $Y=4.135 $X2=8.245
+ $Y2=3.63
cc_383 N_VDD_M1019_b N_A_1469_617#_c_1975_n 0.00155118f $X=-0.05 $Y=2.905
+ $X2=8.33 $Y2=3.795
cc_384 N_VDD_c_261_p N_A_1469_617#_c_1975_n 0.00739652f $X=9.625 $Y=6.507
+ $X2=8.33 $Y2=3.795
cc_385 N_VDD_c_251_p N_A_1469_617#_c_1975_n 0.00475776f $X=9.855 $Y=6.47
+ $X2=8.33 $Y2=3.795
cc_386 N_VDD_M1019_b N_Q_c_1993_n 0.0342497f $X=-0.05 $Y=2.905 $X2=10.14
+ $Y2=4.475
cc_387 N_VDD_c_362_p N_Q_c_1993_n 0.0075728f $X=9.855 $Y=6.44 $X2=10.14
+ $Y2=4.475
cc_388 N_VDD_c_251_p N_Q_c_1993_n 0.00476261f $X=9.855 $Y=6.47 $X2=10.14
+ $Y2=4.475
cc_389 N_VDD_M1019_b N_Q_c_1991_n 0.0127419f $X=-0.05 $Y=2.905 $X2=10.255
+ $Y2=3.16
cc_390 N_VDD_M1019_b N_Q_c_1997_n 0.0207082f $X=-0.05 $Y=2.905 $X2=10.14
+ $Y2=3.287
cc_391 N_VDD_M1019_b Q 0.0106945f $X=-0.05 $Y=2.905 $X2=10.135 $Y2=3.33
cc_392 RN N_A_110_115#_M1019_d 0.00414531f $X=0.325 $Y=3.33 $X2=0.55 $Y2=3.085
cc_393 N_RN_M1017_g N_A_110_115#_c_432_n 0.00386334f $X=0.475 $Y=1.075 $X2=1.29
+ $Y2=2.745
cc_394 N_RN_c_397_n N_A_110_115#_c_432_n 0.00491728f $X=0.475 $Y=2.47 $X2=1.29
+ $Y2=2.745
cc_395 N_RN_M1019_g N_A_110_115#_c_432_n 0.00426455f $X=0.475 $Y=4.585 $X2=1.29
+ $Y2=2.745
cc_396 N_RN_M1017_g N_A_110_115#_c_445_n 0.00500507f $X=0.475 $Y=1.075 $X2=1.29
+ $Y2=1.59
cc_397 N_RN_M1019_g N_A_110_115#_c_454_n 0.00966906f $X=0.475 $Y=4.585 $X2=0.69
+ $Y2=3.455
cc_398 N_RN_c_399_n N_A_110_115#_c_454_n 0.0282684f $X=0.32 $Y=3.33 $X2=0.69
+ $Y2=3.455
cc_399 RN N_A_110_115#_c_454_n 0.00974028f $X=0.325 $Y=3.33 $X2=0.69 $Y2=3.455
cc_400 N_RN_M1017_g N_A_110_115#_c_455_n 0.0102878f $X=0.475 $Y=1.075 $X2=0.87
+ $Y2=2.655
cc_401 N_RN_c_397_n N_A_110_115#_c_455_n 0.00325637f $X=0.475 $Y=2.47 $X2=0.87
+ $Y2=2.655
cc_402 N_RN_M1019_g N_A_110_115#_c_455_n 0.00186244f $X=0.475 $Y=4.585 $X2=0.87
+ $Y2=2.655
cc_403 N_RN_c_399_n N_A_110_115#_c_455_n 0.0072511f $X=0.32 $Y=3.33 $X2=0.87
+ $Y2=2.655
cc_404 N_RN_c_400_n N_A_110_115#_c_455_n 0.0248372f $X=0.32 $Y=2.305 $X2=0.87
+ $Y2=2.655
cc_405 N_RN_M1017_g N_A_110_115#_c_457_n 0.00392272f $X=0.475 $Y=1.075 $X2=0.955
+ $Y2=1.59
cc_406 N_RN_c_397_n N_A_110_115#_c_457_n 0.00143285f $X=0.475 $Y=2.47 $X2=0.955
+ $Y2=1.59
cc_407 N_RN_c_400_n N_A_110_115#_c_457_n 3.54179e-19 $X=0.32 $Y=2.305 $X2=0.955
+ $Y2=1.59
cc_408 N_RN_c_397_n N_A_110_115#_c_458_n 0.00191737f $X=0.475 $Y=2.47 $X2=0.87
+ $Y2=2.74
cc_409 N_RN_M1019_g N_A_110_115#_c_458_n 0.00207383f $X=0.475 $Y=4.585 $X2=0.87
+ $Y2=2.74
cc_410 N_RN_c_399_n N_A_110_115#_c_458_n 0.0113366f $X=0.32 $Y=3.33 $X2=0.87
+ $Y2=2.74
cc_411 N_RN_c_400_n N_A_110_115#_c_458_n 7.08415e-19 $X=0.32 $Y=2.305 $X2=0.87
+ $Y2=2.74
cc_412 N_RN_M1019_g N_A_217_617#_c_1187_n 0.00707175f $X=0.475 $Y=4.585 $X2=1.21
+ $Y2=3.795
cc_413 RN N_A_217_617#_c_1187_n 9.10636e-19 $X=0.325 $Y=3.33 $X2=1.21 $Y2=3.795
cc_414 N_A_110_115#_c_432_n N_SN_M1000_g 0.00495566f $X=1.29 $Y=2.745 $X2=1.855
+ $Y2=4.585
cc_415 N_A_110_115#_c_444_n N_SN_M1000_g 0.0457188f $X=1.425 $Y=2.82 $X2=1.855
+ $Y2=4.585
cc_416 N_A_110_115#_c_434_n N_SN_M1015_g 0.024613f $X=1.435 $Y=1.425 $X2=1.925
+ $Y2=1.075
cc_417 N_A_110_115#_c_445_n N_SN_M1015_g 0.00344794f $X=1.29 $Y=1.59 $X2=1.925
+ $Y2=1.075
cc_418 N_A_110_115#_c_463_n N_SN_M1015_g 0.0106787f $X=8.715 $Y=1.48 $X2=1.925
+ $Y2=1.075
cc_419 N_A_110_115#_c_438_n N_SN_M1002_g 0.0243548f $X=8.535 $Y=1.425 $X2=8.045
+ $Y2=1.075
cc_420 N_A_110_115#_c_448_n N_SN_M1002_g 0.00479479f $X=8.8 $Y=1.59 $X2=8.045
+ $Y2=1.075
cc_421 N_A_110_115#_c_463_n N_SN_M1002_g 0.0110943f $X=8.715 $Y=1.48 $X2=8.045
+ $Y2=1.075
cc_422 N_A_110_115#_c_447_n N_SN_M1035_g 0.0462268f $X=8.8 $Y=2.82 $X2=8.115
+ $Y2=4.585
cc_423 N_A_110_115#_c_432_n N_SN_c_649_n 0.0199681f $X=1.29 $Y=2.745 $X2=1.71
+ $Y2=2.37
cc_424 N_A_110_115#_c_432_n N_SN_c_651_n 0.0112402f $X=1.29 $Y=2.745 $X2=1.89
+ $Y2=1.925
cc_425 N_A_110_115#_c_463_n N_SN_c_651_n 2.91248e-19 $X=8.715 $Y=1.48 $X2=1.89
+ $Y2=1.925
cc_426 N_A_110_115#_c_443_n N_SN_c_652_n 0.00975715f $X=8.8 $Y=2.745 $X2=8.025
+ $Y2=2.255
cc_427 N_A_110_115#_c_463_n N_SN_c_652_n 0.00212668f $X=8.715 $Y=1.48 $X2=8.025
+ $Y2=2.255
cc_428 N_A_110_115#_c_432_n N_SN_c_653_n 0.00177359f $X=1.29 $Y=2.745 $X2=1.71
+ $Y2=2.96
cc_429 N_A_110_115#_c_444_n N_SN_c_653_n 0.00231894f $X=1.425 $Y=2.82 $X2=1.71
+ $Y2=2.96
cc_430 N_A_110_115#_c_432_n N_SN_c_655_n 0.00103414f $X=1.29 $Y=2.745 $X2=1.71
+ $Y2=2.37
cc_431 N_A_110_115#_c_443_n N_SN_c_656_n 2.72295e-19 $X=8.8 $Y=2.745 $X2=8.025
+ $Y2=2.255
cc_432 N_A_110_115#_c_463_n N_SN_c_656_n 0.00342638f $X=8.715 $Y=1.48 $X2=8.025
+ $Y2=2.255
cc_433 N_A_110_115#_c_444_n N_SN_c_658_n 0.00457686f $X=1.425 $Y=2.82 $X2=1.855
+ $Y2=2.96
cc_434 N_A_110_115#_c_447_n SN 0.00111722f $X=8.8 $Y=2.82 $X2=7.935 $Y2=2.96
cc_435 N_A_110_115#_c_463_n N_A_432_520#_M1033_d 0.00558831f $X=8.715 $Y=1.48
+ $X2=3.67 $Y2=0.575
cc_436 N_A_110_115#_c_463_n N_A_432_520#_M1001_g 0.0116352f $X=8.715 $Y=1.48
+ $X2=2.285 $Y2=1.075
cc_437 N_A_110_115#_c_463_n N_A_432_520#_c_818_n 0.0295499f $X=8.715 $Y=1.48
+ $X2=3.71 $Y2=1.765
cc_438 N_A_110_115#_c_463_n N_A_432_520#_c_821_n 0.00540043f $X=8.715 $Y=1.48
+ $X2=2.38 $Y2=1.765
cc_439 N_A_110_115#_c_463_n N_A_432_520#_c_822_n 0.0151351f $X=8.715 $Y=1.48
+ $X2=3.795 $Y2=1.68
cc_440 N_A_110_115#_c_463_n N_A_432_520#_c_844_n 0.0254135f $X=8.715 $Y=1.48
+ $X2=3.887 $Y2=1.415
cc_441 N_A_110_115#_c_463_n N_D_M1005_g 0.0116357f $X=8.715 $Y=1.48 $X2=3.235
+ $Y2=1.075
cc_442 N_A_110_115#_c_463_n N_CK_c_944_n 8.06574e-19 $X=8.715 $Y=1.48 $X2=4.135
+ $Y2=1.85
cc_443 N_A_110_115#_c_463_n N_CK_c_945_n 0.0106495f $X=8.715 $Y=1.48 $X2=4.135
+ $Y2=1.685
cc_444 N_A_110_115#_c_463_n N_CK_c_948_n 8.06574e-19 $X=8.715 $Y=1.48 $X2=5.405
+ $Y2=1.85
cc_445 N_A_110_115#_c_463_n N_CK_c_949_n 0.00177838f $X=8.715 $Y=1.48 $X2=5.405
+ $Y2=1.685
cc_446 N_A_110_115#_c_463_n N_CK_c_953_n 0.01159f $X=8.715 $Y=1.48 $X2=6.762
+ $Y2=1.685
cc_447 N_A_110_115#_c_463_n N_CK_c_958_n 0.00107886f $X=8.715 $Y=1.48 $X2=6.762
+ $Y2=1.835
cc_448 N_A_110_115#_c_463_n N_CK_c_960_n 0.00496158f $X=8.715 $Y=1.48 $X2=4.135
+ $Y2=1.85
cc_449 N_A_110_115#_c_463_n N_CK_c_961_n 0.00118606f $X=8.715 $Y=1.48 $X2=5.405
+ $Y2=1.85
cc_450 N_A_110_115#_c_463_n N_A_217_617#_M1032_d 0.00428739f $X=8.715 $Y=1.48
+ $X2=1.51 $Y2=0.575
cc_451 N_A_110_115#_c_463_n N_A_217_617#_M1021_g 0.0104272f $X=8.715 $Y=1.48
+ $X2=4.555 $Y2=1.075
cc_452 N_A_110_115#_c_463_n N_A_217_617#_c_1178_n 2.42482e-19 $X=8.715 $Y=1.48
+ $X2=4.91 $Y2=1.85
cc_453 N_A_110_115#_c_463_n N_A_217_617#_M1026_g 0.00491871f $X=8.715 $Y=1.48
+ $X2=4.985 $Y2=1.075
cc_454 N_A_110_115#_c_432_n N_A_217_617#_c_1187_n 0.0189043f $X=1.29 $Y=2.745
+ $X2=1.21 $Y2=3.795
cc_455 N_A_110_115#_M1016_g N_A_217_617#_c_1187_n 0.0160567f $X=1.425 $Y=4.585
+ $X2=1.21 $Y2=3.795
cc_456 N_A_110_115#_c_444_n N_A_217_617#_c_1187_n 0.00689282f $X=1.425 $Y=2.82
+ $X2=1.21 $Y2=3.795
cc_457 N_A_110_115#_c_454_n N_A_217_617#_c_1187_n 0.139023f $X=0.69 $Y=3.455
+ $X2=1.21 $Y2=3.795
cc_458 N_A_110_115#_c_455_n N_A_217_617#_c_1187_n 0.041373f $X=0.87 $Y=2.655
+ $X2=1.21 $Y2=3.795
cc_459 N_A_110_115#_c_458_n N_A_217_617#_c_1187_n 0.0134429f $X=0.87 $Y=2.74
+ $X2=1.21 $Y2=3.795
cc_460 N_A_110_115#_c_432_n N_A_217_617#_c_1188_n 0.00793321f $X=1.29 $Y=2.745
+ $X2=1.625 $Y2=2.02
cc_461 N_A_110_115#_c_444_n N_A_217_617#_c_1188_n 0.00344703f $X=1.425 $Y=2.82
+ $X2=1.625 $Y2=2.02
cc_462 N_A_110_115#_c_445_n N_A_217_617#_c_1188_n 0.00409968f $X=1.29 $Y=1.59
+ $X2=1.625 $Y2=2.02
cc_463 N_A_110_115#_c_459_n N_A_217_617#_c_1188_n 0.00447433f $X=1.23 $Y=1.59
+ $X2=1.625 $Y2=2.02
cc_464 N_A_110_115#_c_463_n N_A_217_617#_c_1188_n 0.00645871f $X=8.715 $Y=1.48
+ $X2=1.625 $Y2=2.02
cc_465 N_A_110_115#_c_475_n N_A_217_617#_c_1188_n 4.44945e-19 $X=1.375 $Y=1.48
+ $X2=1.625 $Y2=2.02
cc_466 N_A_110_115#_c_432_n N_A_217_617#_c_1189_n 0.00476027f $X=1.29 $Y=2.745
+ $X2=1.295 $Y2=2.02
cc_467 N_A_110_115#_c_445_n N_A_217_617#_c_1189_n 0.00219831f $X=1.29 $Y=1.59
+ $X2=1.295 $Y2=2.02
cc_468 N_A_110_115#_c_455_n N_A_217_617#_c_1189_n 0.0142869f $X=0.87 $Y=2.655
+ $X2=1.295 $Y2=2.02
cc_469 N_A_110_115#_c_456_n N_A_217_617#_c_1189_n 9.79192e-19 $X=1.145 $Y=1.59
+ $X2=1.295 $Y2=2.02
cc_470 N_A_110_115#_c_459_n N_A_217_617#_c_1189_n 0.00756801f $X=1.23 $Y=1.59
+ $X2=1.295 $Y2=2.02
cc_471 N_A_110_115#_c_475_n N_A_217_617#_c_1189_n 0.00115029f $X=1.375 $Y=1.48
+ $X2=1.295 $Y2=2.02
cc_472 N_A_110_115#_c_434_n N_A_217_617#_c_1190_n 0.0130665f $X=1.435 $Y=1.425
+ $X2=1.71 $Y2=0.825
cc_473 N_A_110_115#_c_445_n N_A_217_617#_c_1190_n 0.00271061f $X=1.29 $Y=1.59
+ $X2=1.71 $Y2=0.825
cc_474 N_A_110_115#_c_455_n N_A_217_617#_c_1190_n 0.00468672f $X=0.87 $Y=2.655
+ $X2=1.71 $Y2=0.825
cc_475 N_A_110_115#_c_459_n N_A_217_617#_c_1190_n 0.0140184f $X=1.23 $Y=1.59
+ $X2=1.71 $Y2=0.825
cc_476 N_A_110_115#_c_463_n N_A_217_617#_c_1190_n 0.0227909f $X=8.715 $Y=1.48
+ $X2=1.71 $Y2=0.825
cc_477 N_A_110_115#_c_475_n N_A_217_617#_c_1190_n 0.00144419f $X=1.375 $Y=1.48
+ $X2=1.71 $Y2=0.825
cc_478 N_A_110_115#_c_463_n N_A_217_617#_c_1194_n 0.00546464f $X=8.715 $Y=1.48
+ $X2=4.725 $Y2=1.85
cc_479 N_A_110_115#_c_463_n N_A_217_617#_c_1196_n 0.212985f $X=8.715 $Y=1.48
+ $X2=4.49 $Y2=1.85
cc_480 N_A_110_115#_c_445_n N_A_217_617#_c_1197_n 0.00390253f $X=1.29 $Y=1.59
+ $X2=1.855 $Y2=1.85
cc_481 N_A_110_115#_c_455_n N_A_217_617#_c_1197_n 0.0049761f $X=0.87 $Y=2.655
+ $X2=1.855 $Y2=1.85
cc_482 N_A_110_115#_c_463_n N_A_217_617#_c_1197_n 0.0252928f $X=8.715 $Y=1.48
+ $X2=1.855 $Y2=1.85
cc_483 N_A_110_115#_c_463_n N_A_217_617#_c_1247_n 0.0259207f $X=8.715 $Y=1.48
+ $X2=4.635 $Y2=1.85
cc_484 N_A_110_115#_c_463_n N_A_704_89#_M1011_d 0.00421798f $X=8.715 $Y=1.48
+ $X2=6.81 $Y2=0.575
cc_485 N_A_110_115#_c_463_n N_A_704_89#_c_1338_n 0.0102209f $X=8.715 $Y=1.48
+ $X2=3.595 $Y2=1.685
cc_486 N_A_110_115#_c_463_n N_A_704_89#_c_1352_n 0.00232964f $X=8.715 $Y=1.48
+ $X2=5.885 $Y2=1.85
cc_487 N_A_110_115#_c_463_n N_A_704_89#_c_1353_n 0.0103799f $X=8.715 $Y=1.48
+ $X2=5.885 $Y2=1.685
cc_488 N_A_110_115#_c_463_n N_A_704_89#_c_1356_n 0.0115848f $X=8.715 $Y=1.48
+ $X2=6.865 $Y2=1.85
cc_489 N_A_110_115#_c_463_n N_A_704_89#_c_1358_n 0.0252668f $X=8.715 $Y=1.48
+ $X2=6.95 $Y2=0.825
cc_490 N_A_110_115#_c_463_n N_A_704_89#_c_1366_n 4.8388e-19 $X=8.715 $Y=1.48
+ $X2=7.22 $Y2=2.19
cc_491 N_A_110_115#_c_463_n N_A_1246_89#_M1002_d 0.00453588f $X=8.715 $Y=1.48
+ $X2=8.12 $Y2=0.575
cc_492 N_A_110_115#_c_463_n N_A_1246_89#_M1006_g 0.0100216f $X=8.715 $Y=1.48
+ $X2=6.305 $Y2=1.075
cc_493 N_A_110_115#_c_448_n N_A_1246_89#_M1007_g 0.00523483f $X=8.8 $Y=1.59
+ $X2=9.495 $Y2=0.945
cc_494 N_A_110_115#_c_443_n N_A_1246_89#_c_1540_n 0.0112463f $X=8.8 $Y=2.745
+ $X2=9.38 $Y2=2.19
cc_495 N_A_110_115#_c_443_n N_A_1246_89#_c_1542_n 0.0059544f $X=8.8 $Y=2.745
+ $X2=9.47 $Y2=1.8
cc_496 N_A_110_115#_c_448_n N_A_1246_89#_c_1542_n 0.0026679f $X=8.8 $Y=1.59
+ $X2=9.47 $Y2=1.8
cc_497 N_A_110_115#_c_443_n N_A_1246_89#_c_1543_n 0.00627484f $X=8.8 $Y=2.745
+ $X2=9.47 $Y2=2.855
cc_498 N_A_110_115#_c_447_n N_A_1246_89#_c_1544_n 0.00627484f $X=8.8 $Y=2.82
+ $X2=9.47 $Y2=3.005
cc_499 N_A_110_115#_c_438_n N_A_1246_89#_c_1546_n 0.0132066f $X=8.535 $Y=1.425
+ $X2=8.26 $Y2=0.825
cc_500 N_A_110_115#_c_448_n N_A_1246_89#_c_1546_n 0.00281336f $X=8.8 $Y=1.59
+ $X2=8.26 $Y2=0.825
cc_501 N_A_110_115#_c_461_n N_A_1246_89#_c_1546_n 0.00937374f $X=8.86 $Y=1.48
+ $X2=8.26 $Y2=0.825
cc_502 N_A_110_115#_c_463_n N_A_1246_89#_c_1546_n 0.0255246f $X=8.715 $Y=1.48
+ $X2=8.26 $Y2=0.825
cc_503 N_A_110_115#_c_477_n N_A_1246_89#_c_1546_n 0.0014036f $X=8.86 $Y=1.48
+ $X2=8.26 $Y2=0.825
cc_504 N_A_110_115#_M1004_g N_A_1246_89#_c_1549_n 0.0166065f $X=8.545 $Y=4.585
+ $X2=8.76 $Y2=3.795
cc_505 N_A_110_115#_c_443_n N_A_1246_89#_c_1549_n 0.0154628f $X=8.8 $Y=2.745
+ $X2=8.76 $Y2=3.795
cc_506 N_A_110_115#_c_447_n N_A_1246_89#_c_1549_n 0.0119447f $X=8.8 $Y=2.82
+ $X2=8.76 $Y2=3.795
cc_507 N_A_110_115#_c_443_n N_A_1246_89#_c_1550_n 0.0122218f $X=8.8 $Y=2.745
+ $X2=8.845 $Y2=2.19
cc_508 N_A_110_115#_c_447_n N_A_1246_89#_c_1550_n 0.00504106f $X=8.8 $Y=2.82
+ $X2=8.845 $Y2=2.19
cc_509 N_A_110_115#_c_448_n N_A_1246_89#_c_1550_n 0.00661521f $X=8.8 $Y=1.59
+ $X2=8.845 $Y2=2.19
cc_510 N_A_110_115#_c_461_n N_A_1246_89#_c_1550_n 0.00327223f $X=8.86 $Y=1.48
+ $X2=8.845 $Y2=2.19
cc_511 N_A_110_115#_c_463_n N_A_1246_89#_c_1550_n 0.00679136f $X=8.715 $Y=1.48
+ $X2=8.845 $Y2=2.19
cc_512 N_A_110_115#_c_477_n N_A_1246_89#_c_1550_n 3.46405e-19 $X=8.86 $Y=1.48
+ $X2=8.845 $Y2=2.19
cc_513 N_A_110_115#_c_443_n N_A_1246_89#_c_1551_n 0.00404253f $X=8.8 $Y=2.745
+ $X2=9.38 $Y2=2.19
cc_514 N_A_110_115#_c_448_n N_A_1246_89#_c_1551_n 0.0023029f $X=8.8 $Y=1.59
+ $X2=9.38 $Y2=2.19
cc_515 N_A_110_115#_c_461_n N_A_1246_89#_c_1551_n 0.00426127f $X=8.86 $Y=1.48
+ $X2=9.38 $Y2=2.19
cc_516 N_A_110_115#_c_477_n N_A_1246_89#_c_1551_n 2.04613e-19 $X=8.86 $Y=1.48
+ $X2=9.38 $Y2=2.19
cc_517 N_A_110_115#_c_443_n N_A_1246_89#_c_1552_n 0.0029248f $X=8.8 $Y=2.745
+ $X2=9.235 $Y2=2.19
cc_518 N_A_110_115#_c_448_n N_A_1246_89#_c_1552_n 0.00182149f $X=8.8 $Y=1.59
+ $X2=9.235 $Y2=2.19
cc_519 N_A_110_115#_c_461_n N_A_1246_89#_c_1552_n 0.00247528f $X=8.86 $Y=1.48
+ $X2=9.235 $Y2=2.19
cc_520 N_A_110_115#_c_463_n N_A_1246_89#_c_1552_n 0.0442421f $X=8.715 $Y=1.48
+ $X2=9.235 $Y2=2.19
cc_521 N_A_110_115#_c_477_n N_A_1246_89#_c_1552_n 0.0129171f $X=8.86 $Y=1.48
+ $X2=9.235 $Y2=2.19
cc_522 N_A_110_115#_c_443_n N_A_1246_89#_c_1554_n 8.29185e-19 $X=8.8 $Y=2.745
+ $X2=9.38 $Y2=2.19
cc_523 N_A_110_115#_c_463_n N_A_1084_115#_M1022_d 0.0051762f $X=8.715 $Y=1.48
+ $X2=5.42 $Y2=0.575
cc_524 N_A_110_115#_c_463_n N_A_1084_115#_c_1706_n 0.0119742f $X=8.715 $Y=1.48
+ $X2=7.685 $Y2=1.69
cc_525 N_A_110_115#_c_463_n N_A_1084_115#_c_1710_n 0.00328689f $X=8.715 $Y=1.48
+ $X2=7.685 $Y2=1.77
cc_526 N_A_110_115#_c_463_n N_A_1084_115#_c_1713_n 0.00616681f $X=8.715 $Y=1.48
+ $X2=5.065 $Y2=1.85
cc_527 N_A_110_115#_c_463_n N_A_1084_115#_c_1738_n 0.0537388f $X=8.715 $Y=1.48
+ $X2=5.475 $Y2=1.43
cc_528 N_A_110_115#_c_463_n N_A_1084_115#_c_1739_n 0.0129425f $X=8.715 $Y=1.48
+ $X2=5.15 $Y2=1.43
cc_529 N_A_110_115#_c_463_n N_A_1084_115#_c_1717_n 0.00241187f $X=8.715 $Y=1.48
+ $X2=7.595 $Y2=1.85
cc_530 N_A_110_115#_c_463_n N_A_1084_115#_c_1719_n 0.186671f $X=8.715 $Y=1.48
+ $X2=7.45 $Y2=1.85
cc_531 N_A_110_115#_c_463_n N_A_1084_115#_c_1722_n 0.0252354f $X=8.715 $Y=1.48
+ $X2=5.21 $Y2=1.85
cc_532 N_A_110_115#_c_463_n N_A_1084_115#_c_1723_n 0.0265552f $X=8.715 $Y=1.48
+ $X2=7.595 $Y2=1.85
cc_533 N_A_110_115#_c_438_n N_QN_c_1867_n 0.00819338f $X=8.535 $Y=1.425 $X2=9.28
+ $Y2=0.825
cc_534 N_A_110_115#_c_448_n N_QN_c_1867_n 0.0028329f $X=8.8 $Y=1.59 $X2=9.28
+ $Y2=0.825
cc_535 N_A_110_115#_c_461_n N_QN_c_1867_n 0.0175339f $X=8.86 $Y=1.48 $X2=9.28
+ $Y2=0.825
cc_536 N_A_110_115#_c_477_n N_QN_c_1867_n 0.0057712f $X=8.86 $Y=1.48 $X2=9.28
+ $Y2=0.825
cc_537 N_A_110_115#_c_447_n N_QN_c_1871_n 3.3286e-19 $X=8.8 $Y=2.82 $X2=9.28
+ $Y2=2.96
cc_538 N_A_110_115#_c_443_n N_QN_c_1873_n 0.00277409f $X=8.8 $Y=2.745 $X2=9.365
+ $Y2=1.85
cc_539 N_A_110_115#_c_443_n N_QN_c_1875_n 0.00166888f $X=8.8 $Y=2.745 $X2=9.365
+ $Y2=2.765
cc_540 N_A_110_115#_c_447_n QN 8.90472e-19 $X=8.8 $Y=2.82 $X2=9.285 $Y2=2.96
cc_541 N_A_110_115#_c_463_n A_400_115# 0.0100396f $X=8.715 $Y=1.48 $X2=2
+ $Y2=0.575
cc_542 N_A_110_115#_c_463_n A_662_115# 0.00911585f $X=8.715 $Y=1.48 $X2=3.31
+ $Y2=0.575
cc_543 N_A_110_115#_c_463_n A_854_115# 0.0100396f $X=8.715 $Y=1.48 $X2=4.27
+ $Y2=0.575
cc_544 N_A_110_115#_c_463_n A_1012_115# 0.00106636f $X=8.715 $Y=1.48 $X2=5.06
+ $Y2=0.575
cc_545 N_A_110_115#_c_463_n A_1204_115# 0.00917995f $X=8.715 $Y=1.48 $X2=6.02
+ $Y2=0.575
cc_546 N_A_110_115#_c_463_n A_1552_115# 0.0106361f $X=8.715 $Y=1.48 $X2=7.76
+ $Y2=0.575
cc_547 N_SN_M1015_g N_A_432_520#_M1001_g 0.0906459f $X=1.925 $Y=1.075 $X2=2.285
+ $Y2=1.075
cc_548 N_SN_c_650_n N_A_432_520#_M1001_g 0.0282237f $X=1.752 $Y=2.205 $X2=2.285
+ $Y2=1.075
cc_549 N_SN_c_653_n N_A_432_520#_M1001_g 3.95753e-19 $X=1.71 $Y=2.96 $X2=2.285
+ $Y2=1.075
cc_550 N_SN_c_655_n N_A_432_520#_M1001_g 5.25039e-19 $X=1.71 $Y=2.37 $X2=2.285
+ $Y2=1.075
cc_551 N_SN_M1000_g N_A_432_520#_M1003_g 0.0523493f $X=1.855 $Y=4.585 $X2=2.285
+ $Y2=4.585
cc_552 N_SN_c_653_n N_A_432_520#_M1003_g 3.16831e-19 $X=1.71 $Y=2.96 $X2=2.285
+ $Y2=4.585
cc_553 N_SN_c_657_n N_A_432_520#_M1003_g 7.19848e-19 $X=7.79 $Y=2.96 $X2=2.285
+ $Y2=4.585
cc_554 N_SN_M1000_g N_A_432_520#_c_816_n 0.0179454f $X=1.855 $Y=4.585 $X2=2.295
+ $Y2=2.765
cc_555 N_SN_c_653_n N_A_432_520#_c_816_n 9.94587e-19 $X=1.71 $Y=2.96 $X2=2.295
+ $Y2=2.765
cc_556 N_SN_c_657_n N_A_432_520#_c_816_n 0.00593089f $X=7.79 $Y=2.96 $X2=2.295
+ $Y2=2.765
cc_557 N_SN_c_650_n N_A_432_520#_c_817_n 0.00496844f $X=1.752 $Y=2.205 $X2=2.295
+ $Y2=2.765
cc_558 N_SN_c_651_n N_A_432_520#_c_817_n 3.15898e-19 $X=1.89 $Y=1.925 $X2=2.295
+ $Y2=2.765
cc_559 N_SN_c_653_n N_A_432_520#_c_817_n 0.0170473f $X=1.71 $Y=2.96 $X2=2.295
+ $Y2=2.765
cc_560 N_SN_c_655_n N_A_432_520#_c_817_n 0.00704947f $X=1.71 $Y=2.37 $X2=2.295
+ $Y2=2.765
cc_561 N_SN_c_657_n N_A_432_520#_c_817_n 0.0236889f $X=7.79 $Y=2.96 $X2=2.295
+ $Y2=2.765
cc_562 N_SN_c_658_n N_A_432_520#_c_817_n 0.00164393f $X=1.855 $Y=2.96 $X2=2.295
+ $Y2=2.765
cc_563 N_SN_M1015_g N_A_432_520#_c_821_n 6.84827e-19 $X=1.925 $Y=1.075 $X2=2.38
+ $Y2=1.765
cc_564 N_SN_c_657_n N_A_432_520#_c_833_n 0.0775662f $X=7.79 $Y=2.96 $X2=3.725
+ $Y2=3.185
cc_565 N_SN_M1000_g N_A_432_520#_c_863_n 0.00105594f $X=1.855 $Y=4.585 $X2=2.38
+ $Y2=3.185
cc_566 N_SN_c_657_n N_D_M1008_g 0.00799543f $X=7.79 $Y=2.96 $X2=3.235 $Y2=4.585
cc_567 N_SN_c_657_n N_D_c_907_n 7.07415e-19 $X=7.79 $Y=2.96 $X2=3.295 $Y2=2.22
cc_568 N_SN_c_657_n N_D_c_908_n 0.00333216f $X=7.79 $Y=2.96 $X2=3.295 $Y2=2.22
cc_569 N_SN_c_657_n D 0.0134431f $X=7.79 $Y=2.96 $X2=3.295 $Y2=2.22
cc_570 N_SN_c_657_n N_CK_M1034_g 0.00294331f $X=7.79 $Y=2.96 $X2=3.595 $Y2=4.585
cc_571 N_SN_c_657_n N_CK_M1020_g 0.00796817f $X=7.79 $Y=2.96 $X2=5.945 $Y2=4.585
cc_572 N_SN_c_657_n N_CK_c_941_n 0.00448328f $X=7.79 $Y=2.96 $X2=6.735 $Y2=2.93
cc_573 N_SN_c_657_n N_CK_M1012_g 0.00909285f $X=7.79 $Y=2.96 $X2=6.735 $Y2=4.585
cc_574 N_SN_c_657_n N_CK_c_943_n 0.00264508f $X=7.79 $Y=2.96 $X2=3.655 $Y2=2.765
cc_575 N_SN_c_657_n N_CK_c_952_n 0.00264508f $X=7.79 $Y=2.96 $X2=5.885 $Y2=2.765
cc_576 N_SN_c_657_n N_CK_c_959_n 0.003555f $X=7.79 $Y=2.96 $X2=4.05 $Y2=2.59
cc_577 N_SN_c_657_n N_CK_c_962_n 0.00141703f $X=7.79 $Y=2.96 $X2=5.8 $Y2=2.59
cc_578 N_SN_c_657_n N_CK_c_963_n 9.71861e-19 $X=7.79 $Y=2.96 $X2=5.49 $Y2=2.59
cc_579 N_SN_c_657_n N_CK_c_964_n 0.00700078f $X=7.79 $Y=2.96 $X2=6.88 $Y2=2.59
cc_580 N_SN_c_657_n N_CK_c_965_n 0.00732128f $X=7.79 $Y=2.96 $X2=3.655 $Y2=2.59
cc_581 N_SN_c_657_n N_CK_c_966_n 0.00860578f $X=7.79 $Y=2.96 $X2=5.885 $Y2=2.59
cc_582 N_SN_c_657_n N_CK_c_967_n 0.15926f $X=7.79 $Y=2.96 $X2=5.74 $Y2=2.59
cc_583 N_SN_c_657_n N_CK_c_968_n 0.0251654f $X=7.79 $Y=2.96 $X2=3.8 $Y2=2.59
cc_584 N_SN_c_657_n N_CK_c_969_n 0.0598286f $X=7.79 $Y=2.96 $X2=6.735 $Y2=2.59
cc_585 N_SN_c_657_n N_CK_c_970_n 0.0251663f $X=7.79 $Y=2.96 $X2=6.03 $Y2=2.59
cc_586 N_SN_c_657_n CK 0.025144f $X=7.79 $Y=2.96 $X2=6.88 $Y2=2.59
cc_587 N_SN_c_657_n N_A_217_617#_M1024_g 0.00827407f $X=7.79 $Y=2.96 $X2=4.555
+ $Y2=4.585
cc_588 N_SN_c_657_n N_A_217_617#_c_1181_n 0.00177706f $X=7.79 $Y=2.96 $X2=4.91
+ $Y2=2.765
cc_589 N_SN_c_657_n N_A_217_617#_c_1182_n 0.00157006f $X=7.79 $Y=2.96 $X2=4.63
+ $Y2=2.765
cc_590 N_SN_c_657_n N_A_217_617#_M1027_g 0.00382698f $X=7.79 $Y=2.96 $X2=4.985
+ $Y2=4.585
cc_591 N_SN_M1000_g N_A_217_617#_c_1187_n 3.2027e-19 $X=1.855 $Y=4.585 $X2=1.21
+ $Y2=3.795
cc_592 N_SN_c_649_n N_A_217_617#_c_1187_n 9.40033e-19 $X=1.71 $Y=2.37 $X2=1.21
+ $Y2=3.795
cc_593 N_SN_c_650_n N_A_217_617#_c_1187_n 5.0101e-19 $X=1.752 $Y=2.205 $X2=1.21
+ $Y2=3.795
cc_594 N_SN_c_653_n N_A_217_617#_c_1187_n 0.0231905f $X=1.71 $Y=2.96 $X2=1.21
+ $Y2=3.795
cc_595 N_SN_c_655_n N_A_217_617#_c_1187_n 0.00963813f $X=1.71 $Y=2.37 $X2=1.21
+ $Y2=3.795
cc_596 N_SN_c_658_n N_A_217_617#_c_1187_n 0.00754015f $X=1.855 $Y=2.96 $X2=1.21
+ $Y2=3.795
cc_597 N_SN_c_649_n N_A_217_617#_c_1188_n 0.00517882f $X=1.71 $Y=2.37 $X2=1.625
+ $Y2=2.02
cc_598 N_SN_c_650_n N_A_217_617#_c_1188_n 0.00527195f $X=1.752 $Y=2.205
+ $X2=1.625 $Y2=2.02
cc_599 N_SN_c_655_n N_A_217_617#_c_1188_n 0.0186534f $X=1.71 $Y=2.37 $X2=1.625
+ $Y2=2.02
cc_600 N_SN_M1015_g N_A_217_617#_c_1190_n 0.00641257f $X=1.925 $Y=1.075 $X2=1.71
+ $Y2=0.825
cc_601 N_SN_c_651_n N_A_217_617#_c_1190_n 0.00374345f $X=1.89 $Y=1.925 $X2=1.71
+ $Y2=0.825
cc_602 N_SN_c_657_n N_A_217_617#_c_1193_n 0.00880485f $X=7.79 $Y=2.96 $X2=4.725
+ $Y2=2.765
cc_603 N_SN_M1015_g N_A_217_617#_c_1196_n 0.00153565f $X=1.925 $Y=1.075 $X2=4.49
+ $Y2=1.85
cc_604 N_SN_c_650_n N_A_217_617#_c_1196_n 0.00261695f $X=1.752 $Y=2.205 $X2=4.49
+ $Y2=1.85
cc_605 N_SN_c_651_n N_A_217_617#_c_1196_n 0.00200303f $X=1.89 $Y=1.925 $X2=4.49
+ $Y2=1.85
cc_606 N_SN_c_655_n N_A_217_617#_c_1196_n 5.85585e-19 $X=1.71 $Y=2.37 $X2=4.49
+ $Y2=1.85
cc_607 N_SN_M1015_g N_A_217_617#_c_1197_n 5.70836e-19 $X=1.925 $Y=1.075
+ $X2=1.855 $Y2=1.85
cc_608 N_SN_c_650_n N_A_217_617#_c_1197_n 9.78592e-19 $X=1.752 $Y=2.205
+ $X2=1.855 $Y2=1.85
cc_609 N_SN_c_651_n N_A_217_617#_c_1197_n 4.80352e-19 $X=1.89 $Y=1.925 $X2=1.855
+ $Y2=1.85
cc_610 N_SN_c_655_n N_A_217_617#_c_1197_n 0.00329414f $X=1.71 $Y=2.37 $X2=1.855
+ $Y2=1.85
cc_611 N_SN_c_657_n N_A_704_89#_M1031_g 0.0108138f $X=7.79 $Y=2.96 $X2=4.195
+ $Y2=4.585
cc_612 N_SN_c_657_n N_A_704_89#_M1025_g 0.00578896f $X=7.79 $Y=2.96 $X2=5.345
+ $Y2=4.585
cc_613 N_SN_c_654_n N_A_704_89#_c_1364_n 0.00228032f $X=7.935 $Y=2.96 $X2=7.22
+ $Y2=3.1
cc_614 N_SN_c_657_n N_A_704_89#_c_1364_n 0.0163748f $X=7.79 $Y=2.96 $X2=7.22
+ $Y2=3.1
cc_615 SN N_A_704_89#_c_1364_n 0.00108239f $X=7.935 $Y=2.96 $X2=7.22 $Y2=3.1
cc_616 N_SN_c_657_n N_A_704_89#_c_1366_n 0.00232295f $X=7.79 $Y=2.96 $X2=7.22
+ $Y2=2.19
cc_617 N_SN_c_657_n N_A_704_89#_c_1377_n 0.0135346f $X=7.79 $Y=2.96 $X2=7.22
+ $Y2=3.185
cc_618 N_SN_c_657_n N_A_1246_89#_M1009_g 0.0105543f $X=7.79 $Y=2.96 $X2=6.305
+ $Y2=4.585
cc_619 N_SN_M1002_g N_A_1246_89#_c_1546_n 0.00967483f $X=8.045 $Y=1.075 $X2=8.26
+ $Y2=0.825
cc_620 N_SN_M1035_g N_A_1246_89#_c_1549_n 3.98669e-19 $X=8.115 $Y=4.585 $X2=8.76
+ $Y2=3.795
cc_621 N_SN_c_652_n N_A_1246_89#_c_1549_n 0.00375577f $X=8.025 $Y=2.255 $X2=8.76
+ $Y2=3.795
cc_622 N_SN_c_654_n N_A_1246_89#_c_1549_n 0.0149392f $X=7.935 $Y=2.96 $X2=8.76
+ $Y2=3.795
cc_623 N_SN_c_656_n N_A_1246_89#_c_1549_n 0.00492795f $X=8.025 $Y=2.255 $X2=8.76
+ $Y2=3.795
cc_624 SN N_A_1246_89#_c_1549_n 0.00496818f $X=7.935 $Y=2.96 $X2=8.76 $Y2=3.795
cc_625 N_SN_M1002_g N_A_1246_89#_c_1550_n 0.00483036f $X=8.045 $Y=1.075
+ $X2=8.845 $Y2=2.19
cc_626 N_SN_c_652_n N_A_1246_89#_c_1550_n 0.0026134f $X=8.025 $Y=2.255 $X2=8.845
+ $Y2=2.19
cc_627 N_SN_c_656_n N_A_1246_89#_c_1550_n 0.00832911f $X=8.025 $Y=2.255
+ $X2=8.845 $Y2=2.19
cc_628 N_SN_c_652_n N_A_1246_89#_c_1552_n 0.00614421f $X=8.025 $Y=2.255
+ $X2=9.235 $Y2=2.19
cc_629 N_SN_c_654_n N_A_1246_89#_c_1552_n 9.11589e-19 $X=7.935 $Y=2.96 $X2=9.235
+ $Y2=2.19
cc_630 N_SN_c_656_n N_A_1246_89#_c_1552_n 0.020493f $X=8.025 $Y=2.255 $X2=9.235
+ $Y2=2.19
cc_631 N_SN_M1002_g N_A_1084_115#_c_1705_n 0.00627778f $X=8.045 $Y=1.075
+ $X2=7.505 $Y2=2.63
cc_632 N_SN_M1035_g N_A_1084_115#_c_1705_n 0.00402616f $X=8.115 $Y=4.585
+ $X2=7.505 $Y2=2.63
cc_633 N_SN_c_652_n N_A_1084_115#_c_1705_n 0.0138276f $X=8.025 $Y=2.255
+ $X2=7.505 $Y2=2.63
cc_634 N_SN_c_654_n N_A_1084_115#_c_1705_n 5.97554e-19 $X=7.935 $Y=2.96
+ $X2=7.505 $Y2=2.63
cc_635 N_SN_c_656_n N_A_1084_115#_c_1705_n 6.33368e-19 $X=8.025 $Y=2.255
+ $X2=7.505 $Y2=2.63
cc_636 N_SN_M1002_g N_A_1084_115#_c_1706_n 0.0853563f $X=8.045 $Y=1.075
+ $X2=7.685 $Y2=1.69
cc_637 N_SN_c_657_n N_A_1084_115#_M1014_g 0.00486063f $X=7.79 $Y=2.96 $X2=7.685
+ $Y2=4.585
cc_638 SN N_A_1084_115#_M1014_g 5.06369e-19 $X=7.935 $Y=2.96 $X2=7.685 $Y2=4.585
cc_639 N_SN_M1035_g N_A_1084_115#_c_1712_n 0.0664f $X=8.115 $Y=4.585 $X2=7.685
+ $Y2=2.765
cc_640 N_SN_c_654_n N_A_1084_115#_c_1712_n 0.00312462f $X=7.935 $Y=2.96
+ $X2=7.685 $Y2=2.765
cc_641 N_SN_c_657_n N_A_1084_115#_c_1712_n 0.00760041f $X=7.79 $Y=2.96 $X2=7.685
+ $Y2=2.765
cc_642 SN N_A_1084_115#_c_1712_n 5.28053e-19 $X=7.935 $Y=2.96 $X2=7.685
+ $Y2=2.765
cc_643 N_SN_c_657_n N_A_1084_115#_c_1713_n 0.0225202f $X=7.79 $Y=2.96 $X2=5.065
+ $Y2=1.85
cc_644 N_SN_c_657_n N_A_1084_115#_c_1757_n 0.0256731f $X=7.79 $Y=2.96 $X2=5.475
+ $Y2=3.185
cc_645 N_SN_M1002_g N_A_1084_115#_c_1717_n 0.00316718f $X=8.045 $Y=1.075
+ $X2=7.595 $Y2=1.85
cc_646 N_SN_c_652_n N_A_1084_115#_c_1717_n 0.00203974f $X=8.025 $Y=2.255
+ $X2=7.595 $Y2=1.85
cc_647 N_SN_c_654_n N_A_1084_115#_c_1717_n 0.0367765f $X=7.935 $Y=2.96 $X2=7.595
+ $Y2=1.85
cc_648 N_SN_c_656_n N_A_1084_115#_c_1717_n 0.0189565f $X=8.025 $Y=2.255
+ $X2=7.595 $Y2=1.85
cc_649 N_SN_c_657_n N_A_1084_115#_c_1717_n 0.0136826f $X=7.79 $Y=2.96 $X2=7.595
+ $Y2=1.85
cc_650 SN N_A_1084_115#_c_1717_n 9.02875e-19 $X=7.935 $Y=2.96 $X2=7.595 $Y2=1.85
cc_651 N_SN_M1002_g N_A_1084_115#_c_1723_n 0.00271237f $X=8.045 $Y=1.075
+ $X2=7.595 $Y2=1.85
cc_652 N_SN_M1000_g N_A_300_617#_c_1949_n 0.0147079f $X=1.855 $Y=4.585 $X2=2.415
+ $Y2=3.63
cc_653 N_SN_c_653_n N_A_300_617#_c_1949_n 8.68455e-19 $X=1.71 $Y=2.96 $X2=2.415
+ $Y2=3.63
cc_654 N_SN_c_657_n N_A_300_617#_c_1949_n 0.0122781f $X=7.79 $Y=2.96 $X2=2.415
+ $Y2=3.63
cc_655 N_SN_c_658_n N_A_300_617#_c_1949_n 0.00326201f $X=1.855 $Y=2.96 $X2=2.415
+ $Y2=3.63
cc_656 N_SN_c_653_n N_A_300_617#_c_1960_n 0.00230057f $X=1.71 $Y=2.96 $X2=1.725
+ $Y2=3.63
cc_657 N_SN_c_658_n N_A_300_617#_c_1960_n 0.00491504f $X=1.855 $Y=2.96 $X2=1.725
+ $Y2=3.63
cc_658 N_SN_M1035_g N_A_1469_617#_c_1973_n 0.0171268f $X=8.115 $Y=4.585
+ $X2=8.245 $Y2=3.63
cc_659 N_SN_c_654_n N_A_1469_617#_c_1973_n 0.0032182f $X=7.935 $Y=2.96 $X2=8.245
+ $Y2=3.63
cc_660 N_SN_c_657_n N_A_1469_617#_c_1973_n 0.0055835f $X=7.79 $Y=2.96 $X2=8.245
+ $Y2=3.63
cc_661 SN N_A_1469_617#_c_1973_n 0.00793147f $X=7.935 $Y=2.96 $X2=8.245 $Y2=3.63
cc_662 N_SN_c_657_n N_A_1469_617#_c_1982_n 0.00594846f $X=7.79 $Y=2.96 $X2=7.555
+ $Y2=3.63
cc_663 N_A_432_520#_c_818_n N_D_M1005_g 0.0123125f $X=3.71 $Y=1.765 $X2=3.235
+ $Y2=1.075
cc_664 N_A_432_520#_c_833_n N_D_M1008_g 0.0167212f $X=3.725 $Y=3.185 $X2=3.235
+ $Y2=4.585
cc_665 N_A_432_520#_c_818_n N_D_c_907_n 0.00207628f $X=3.71 $Y=1.765 $X2=3.295
+ $Y2=2.22
cc_666 N_A_432_520#_c_818_n N_D_c_908_n 0.0086486f $X=3.71 $Y=1.765 $X2=3.295
+ $Y2=2.22
cc_667 N_A_432_520#_c_818_n D 0.00200799f $X=3.71 $Y=1.765 $X2=3.295 $Y2=2.22
cc_668 N_A_432_520#_c_833_n N_CK_M1034_g 0.0150535f $X=3.725 $Y=3.185 $X2=3.595
+ $Y2=4.585
cc_669 N_A_432_520#_c_833_n N_CK_c_943_n 0.00123101f $X=3.725 $Y=3.185 $X2=3.655
+ $Y2=2.765
cc_670 N_A_432_520#_c_818_n N_CK_c_944_n 9.45214e-19 $X=3.71 $Y=1.765 $X2=4.135
+ $Y2=1.85
cc_671 N_A_432_520#_c_844_n N_CK_c_944_n 0.00170561f $X=3.887 $Y=1.415 $X2=4.135
+ $Y2=1.85
cc_672 N_A_432_520#_c_822_n N_CK_c_945_n 0.00464203f $X=3.795 $Y=1.68 $X2=4.135
+ $Y2=1.685
cc_673 N_A_432_520#_c_844_n N_CK_c_945_n 0.00545632f $X=3.887 $Y=1.415 $X2=4.135
+ $Y2=1.685
cc_674 N_A_432_520#_c_818_n N_CK_c_959_n 0.0019742f $X=3.71 $Y=1.765 $X2=4.05
+ $Y2=2.59
cc_675 N_A_432_520#_c_833_n N_CK_c_959_n 0.00786738f $X=3.725 $Y=3.185 $X2=4.05
+ $Y2=2.59
cc_676 N_A_432_520#_c_818_n N_CK_c_960_n 0.012316f $X=3.71 $Y=1.765 $X2=4.135
+ $Y2=1.85
cc_677 N_A_432_520#_c_844_n N_CK_c_960_n 5.28119e-19 $X=3.887 $Y=1.415 $X2=4.135
+ $Y2=1.85
cc_678 N_A_432_520#_c_818_n N_CK_c_965_n 0.00224444f $X=3.71 $Y=1.765 $X2=3.655
+ $Y2=2.59
cc_679 N_A_432_520#_c_833_n N_CK_c_965_n 0.0085861f $X=3.725 $Y=3.185 $X2=3.655
+ $Y2=2.59
cc_680 N_A_432_520#_M1001_g N_A_217_617#_c_1188_n 4.92509e-19 $X=2.285 $Y=1.075
+ $X2=1.625 $Y2=2.02
cc_681 N_A_432_520#_c_817_n N_A_217_617#_c_1188_n 0.00578504f $X=2.295 $Y=2.765
+ $X2=1.625 $Y2=2.02
cc_682 N_A_432_520#_M1001_g N_A_217_617#_c_1190_n 3.35752e-19 $X=2.285 $Y=1.075
+ $X2=1.71 $Y2=0.825
cc_683 N_A_432_520#_c_817_n N_A_217_617#_c_1190_n 0.00179268f $X=2.295 $Y=2.765
+ $X2=1.71 $Y2=0.825
cc_684 N_A_432_520#_c_821_n N_A_217_617#_c_1190_n 0.00488587f $X=2.38 $Y=1.765
+ $X2=1.71 $Y2=0.825
cc_685 N_A_432_520#_M1001_g N_A_217_617#_c_1196_n 8.50336e-19 $X=2.285 $Y=1.075
+ $X2=4.49 $Y2=1.85
cc_686 N_A_432_520#_c_817_n N_A_217_617#_c_1196_n 0.0151086f $X=2.295 $Y=2.765
+ $X2=4.49 $Y2=1.85
cc_687 N_A_432_520#_c_818_n N_A_217_617#_c_1196_n 0.0578899f $X=3.71 $Y=1.765
+ $X2=4.49 $Y2=1.85
cc_688 N_A_432_520#_c_821_n N_A_217_617#_c_1196_n 0.00475107f $X=2.38 $Y=1.765
+ $X2=4.49 $Y2=1.85
cc_689 N_A_432_520#_c_844_n N_A_217_617#_c_1196_n 8.61924e-19 $X=3.887 $Y=1.415
+ $X2=4.49 $Y2=1.85
cc_690 N_A_432_520#_c_817_n N_A_217_617#_c_1197_n 6.43558e-19 $X=2.295 $Y=2.765
+ $X2=1.855 $Y2=1.85
cc_691 N_A_432_520#_c_821_n N_A_217_617#_c_1197_n 6.84883e-19 $X=2.38 $Y=1.765
+ $X2=1.855 $Y2=1.85
cc_692 N_A_432_520#_c_818_n N_A_704_89#_c_1338_n 0.0022787f $X=3.71 $Y=1.765
+ $X2=3.595 $Y2=1.685
cc_693 N_A_432_520#_c_844_n N_A_704_89#_c_1338_n 0.0060945f $X=3.887 $Y=1.415
+ $X2=3.595 $Y2=1.685
cc_694 N_A_432_520#_c_818_n N_A_704_89#_c_1341_n 0.00324141f $X=3.71 $Y=1.765
+ $X2=3.715 $Y2=2.225
cc_695 N_A_432_520#_c_818_n N_A_704_89#_c_1349_n 0.00993431f $X=3.71 $Y=1.765
+ $X2=3.715 $Y2=1.76
cc_696 N_A_432_520#_c_833_n N_A_300_617#_M1003_d 0.00690809f $X=3.725 $Y=3.185
+ $X2=2.36 $Y2=3.085
cc_697 N_A_432_520#_M1003_g N_A_300_617#_c_1949_n 0.0144978f $X=2.285 $Y=4.585
+ $X2=2.415 $Y2=3.63
cc_698 N_A_432_520#_c_833_n N_A_300_617#_c_1949_n 0.00856071f $X=3.725 $Y=3.185
+ $X2=2.415 $Y2=3.63
cc_699 N_A_432_520#_c_863_n N_A_300_617#_c_1949_n 0.0070523f $X=2.38 $Y=3.185
+ $X2=2.415 $Y2=3.63
cc_700 N_A_432_520#_c_833_n A_662_617# 0.00481059f $X=3.725 $Y=3.185 $X2=3.31
+ $Y2=3.085
cc_701 N_D_M1008_g N_CK_c_943_n 0.216757f $X=3.235 $Y=4.585 $X2=3.655 $Y2=2.765
cc_702 N_D_c_907_n N_CK_c_960_n 2.89615e-19 $X=3.295 $Y=2.22 $X2=4.135 $Y2=1.85
cc_703 N_D_c_908_n N_CK_c_960_n 0.00478177f $X=3.295 $Y=2.22 $X2=4.135 $Y2=1.85
cc_704 D N_CK_c_960_n 0.00551577f $X=3.295 $Y=2.22 $X2=4.135 $Y2=1.85
cc_705 N_D_M1008_g N_CK_c_965_n 0.00512934f $X=3.235 $Y=4.585 $X2=3.655 $Y2=2.59
cc_706 N_D_M1008_g N_CK_c_968_n 0.00515433f $X=3.235 $Y=4.585 $X2=3.8 $Y2=2.59
cc_707 D N_CK_c_968_n 0.00375733f $X=3.295 $Y=2.22 $X2=3.8 $Y2=2.59
cc_708 N_D_M1005_g N_A_217_617#_c_1196_n 0.00303372f $X=3.235 $Y=1.075 $X2=4.49
+ $Y2=1.85
cc_709 N_D_c_907_n N_A_217_617#_c_1196_n 7.9412e-19 $X=3.295 $Y=2.22 $X2=4.49
+ $Y2=1.85
cc_710 N_D_c_908_n N_A_217_617#_c_1196_n 0.00111625f $X=3.295 $Y=2.22 $X2=4.49
+ $Y2=1.85
cc_711 D N_A_217_617#_c_1196_n 0.0353362f $X=3.295 $Y=2.22 $X2=4.49 $Y2=1.85
cc_712 N_D_M1005_g N_A_704_89#_c_1338_n 0.0846533f $X=3.235 $Y=1.075 $X2=3.595
+ $Y2=1.685
cc_713 N_D_M1005_g N_A_704_89#_c_1341_n 0.00932846f $X=3.235 $Y=1.075 $X2=3.715
+ $Y2=2.225
cc_714 N_D_c_907_n N_A_704_89#_c_1341_n 0.0210215f $X=3.295 $Y=2.22 $X2=3.715
+ $Y2=2.225
cc_715 N_D_c_908_n N_A_704_89#_c_1341_n 0.00164409f $X=3.295 $Y=2.22 $X2=3.715
+ $Y2=2.225
cc_716 D N_A_704_89#_c_1341_n 0.00342011f $X=3.295 $Y=2.22 $X2=3.715 $Y2=2.225
cc_717 D N_A_704_89#_c_1343_n 4.62757e-19 $X=3.295 $Y=2.22 $X2=3.79 $Y2=2.3
cc_718 N_CK_c_945_n N_A_217_617#_M1021_g 0.0483944f $X=4.135 $Y=1.685 $X2=4.555
+ $Y2=1.075
cc_719 N_CK_c_960_n N_A_217_617#_M1021_g 0.00109079f $X=4.135 $Y=1.85 $X2=4.555
+ $Y2=1.075
cc_720 N_CK_c_948_n N_A_217_617#_c_1178_n 0.0473482f $X=5.405 $Y=1.85 $X2=4.91
+ $Y2=1.85
cc_721 N_CK_c_944_n N_A_217_617#_c_1180_n 0.0483944f $X=4.135 $Y=1.85 $X2=4.63
+ $Y2=1.85
cc_722 N_CK_c_967_n N_A_217_617#_c_1181_n 0.00203319f $X=5.74 $Y=2.59 $X2=4.91
+ $Y2=2.765
cc_723 N_CK_c_967_n N_A_217_617#_c_1182_n 0.00203351f $X=5.74 $Y=2.59 $X2=4.63
+ $Y2=2.765
cc_724 N_CK_c_949_n N_A_217_617#_M1026_g 0.0473482f $X=5.405 $Y=1.685 $X2=4.985
+ $Y2=1.075
cc_725 N_CK_c_961_n N_A_217_617#_M1026_g 3.67139e-19 $X=5.405 $Y=1.85 $X2=4.985
+ $Y2=1.075
cc_726 N_CK_c_944_n N_A_217_617#_c_1193_n 7.30049e-19 $X=4.135 $Y=1.85 $X2=4.725
+ $Y2=2.765
cc_727 N_CK_c_959_n N_A_217_617#_c_1193_n 0.00401809f $X=4.05 $Y=2.59 $X2=4.725
+ $Y2=2.765
cc_728 N_CK_c_960_n N_A_217_617#_c_1193_n 0.0203851f $X=4.135 $Y=1.85 $X2=4.725
+ $Y2=2.765
cc_729 N_CK_c_967_n N_A_217_617#_c_1193_n 0.0154699f $X=5.74 $Y=2.59 $X2=4.725
+ $Y2=2.765
cc_730 N_CK_c_944_n N_A_217_617#_c_1194_n 7.18106e-19 $X=4.135 $Y=1.85 $X2=4.725
+ $Y2=1.85
cc_731 N_CK_c_960_n N_A_217_617#_c_1194_n 0.00742068f $X=4.135 $Y=1.85 $X2=4.725
+ $Y2=1.85
cc_732 N_CK_c_967_n N_A_217_617#_c_1194_n 0.00102309f $X=5.74 $Y=2.59 $X2=4.725
+ $Y2=1.85
cc_733 N_CK_c_944_n N_A_217_617#_c_1196_n 0.00383172f $X=4.135 $Y=1.85 $X2=4.49
+ $Y2=1.85
cc_734 N_CK_c_959_n N_A_217_617#_c_1196_n 0.00443421f $X=4.05 $Y=2.59 $X2=4.49
+ $Y2=1.85
cc_735 N_CK_c_960_n N_A_217_617#_c_1196_n 0.0149977f $X=4.135 $Y=1.85 $X2=4.49
+ $Y2=1.85
cc_736 N_CK_c_965_n N_A_217_617#_c_1196_n 7.12046e-19 $X=3.655 $Y=2.59 $X2=4.49
+ $Y2=1.85
cc_737 N_CK_c_968_n N_A_217_617#_c_1196_n 0.0126164f $X=3.8 $Y=2.59 $X2=4.49
+ $Y2=1.85
cc_738 N_CK_c_944_n N_A_217_617#_c_1247_n 3.3031e-19 $X=4.135 $Y=1.85 $X2=4.635
+ $Y2=1.85
cc_739 N_CK_c_960_n N_A_217_617#_c_1247_n 0.00143592f $X=4.135 $Y=1.85 $X2=4.635
+ $Y2=1.85
cc_740 N_CK_c_967_n N_A_217_617#_c_1247_n 0.0129652f $X=5.74 $Y=2.59 $X2=4.635
+ $Y2=1.85
cc_741 N_CK_c_945_n N_A_704_89#_c_1338_n 0.0252931f $X=4.135 $Y=1.685 $X2=3.595
+ $Y2=1.685
cc_742 N_CK_c_960_n N_A_704_89#_c_1341_n 0.00613747f $X=4.135 $Y=1.85 $X2=3.715
+ $Y2=2.225
cc_743 N_CK_c_944_n N_A_704_89#_c_1342_n 0.0183603f $X=4.135 $Y=1.85 $X2=4.12
+ $Y2=2.3
cc_744 N_CK_c_960_n N_A_704_89#_c_1342_n 0.00630484f $X=4.135 $Y=1.85 $X2=4.12
+ $Y2=2.3
cc_745 N_CK_c_967_n N_A_704_89#_c_1342_n 0.00613485f $X=5.74 $Y=2.59 $X2=4.12
+ $Y2=2.3
cc_746 N_CK_c_943_n N_A_704_89#_c_1343_n 0.00904036f $X=3.655 $Y=2.765 $X2=3.79
+ $Y2=2.3
cc_747 N_CK_c_959_n N_A_704_89#_c_1343_n 0.00878348f $X=4.05 $Y=2.59 $X2=3.79
+ $Y2=2.3
cc_748 N_CK_c_965_n N_A_704_89#_c_1343_n 0.00109468f $X=3.655 $Y=2.59 $X2=3.79
+ $Y2=2.3
cc_749 N_CK_c_968_n N_A_704_89#_c_1343_n 0.00137501f $X=3.8 $Y=2.59 $X2=3.79
+ $Y2=2.3
cc_750 N_CK_M1034_g N_A_704_89#_M1031_g 0.060745f $X=3.595 $Y=4.585 $X2=4.195
+ $Y2=4.585
cc_751 N_CK_c_943_n N_A_704_89#_M1031_g 0.0129692f $X=3.655 $Y=2.765 $X2=4.195
+ $Y2=4.585
cc_752 N_CK_c_959_n N_A_704_89#_M1031_g 0.0081071f $X=4.05 $Y=2.59 $X2=4.195
+ $Y2=4.585
cc_753 N_CK_c_960_n N_A_704_89#_M1031_g 0.00478024f $X=4.135 $Y=1.85 $X2=4.195
+ $Y2=4.585
cc_754 N_CK_c_965_n N_A_704_89#_M1031_g 0.00197555f $X=3.655 $Y=2.59 $X2=4.195
+ $Y2=4.585
cc_755 N_CK_c_967_n N_A_704_89#_M1031_g 0.00462358f $X=5.74 $Y=2.59 $X2=4.195
+ $Y2=4.585
cc_756 N_CK_c_968_n N_A_704_89#_M1031_g 4.2e-19 $X=3.8 $Y=2.59 $X2=4.195
+ $Y2=4.585
cc_757 N_CK_c_967_n N_A_704_89#_c_1345_n 0.00607908f $X=5.74 $Y=2.59 $X2=5.27
+ $Y2=2.3
cc_758 N_CK_M1020_g N_A_704_89#_M1025_g 0.0607514f $X=5.945 $Y=4.585 $X2=5.345
+ $Y2=4.585
cc_759 N_CK_c_952_n N_A_704_89#_M1025_g 0.0122143f $X=5.885 $Y=2.765 $X2=5.345
+ $Y2=4.585
cc_760 N_CK_c_961_n N_A_704_89#_M1025_g 0.00399495f $X=5.405 $Y=1.85 $X2=5.345
+ $Y2=4.585
cc_761 N_CK_c_963_n N_A_704_89#_M1025_g 0.00654233f $X=5.49 $Y=2.59 $X2=5.345
+ $Y2=4.585
cc_762 N_CK_c_966_n N_A_704_89#_M1025_g 0.00130061f $X=5.885 $Y=2.59 $X2=5.345
+ $Y2=4.585
cc_763 N_CK_c_967_n N_A_704_89#_M1025_g 0.00422185f $X=5.74 $Y=2.59 $X2=5.345
+ $Y2=4.585
cc_764 N_CK_c_970_n N_A_704_89#_M1025_g 4.2e-19 $X=6.03 $Y=2.59 $X2=5.345
+ $Y2=4.585
cc_765 N_CK_c_952_n N_A_704_89#_c_1347_n 0.00904036f $X=5.885 $Y=2.765 $X2=5.75
+ $Y2=2.3
cc_766 N_CK_c_961_n N_A_704_89#_c_1347_n 0.00909647f $X=5.405 $Y=1.85 $X2=5.75
+ $Y2=2.3
cc_767 N_CK_c_962_n N_A_704_89#_c_1347_n 0.00924811f $X=5.8 $Y=2.59 $X2=5.75
+ $Y2=2.3
cc_768 N_CK_c_966_n N_A_704_89#_c_1347_n 0.00102633f $X=5.885 $Y=2.59 $X2=5.75
+ $Y2=2.3
cc_769 N_CK_c_967_n N_A_704_89#_c_1347_n 0.00613485f $X=5.74 $Y=2.59 $X2=5.75
+ $Y2=2.3
cc_770 N_CK_c_970_n N_A_704_89#_c_1347_n 0.00137501f $X=6.03 $Y=2.59 $X2=5.75
+ $Y2=2.3
cc_771 N_CK_c_961_n N_A_704_89#_c_1348_n 0.00649764f $X=5.405 $Y=1.85 $X2=5.825
+ $Y2=2.225
cc_772 N_CK_c_944_n N_A_704_89#_c_1349_n 0.0216263f $X=4.135 $Y=1.85 $X2=3.715
+ $Y2=1.76
cc_773 N_CK_c_965_n N_A_704_89#_c_1349_n 2.45465e-19 $X=3.655 $Y=2.59 $X2=3.715
+ $Y2=1.76
cc_774 N_CK_c_960_n N_A_704_89#_c_1350_n 0.00568091f $X=4.135 $Y=1.85 $X2=4.195
+ $Y2=2.3
cc_775 N_CK_c_948_n N_A_704_89#_c_1351_n 0.0183603f $X=5.405 $Y=1.85 $X2=5.345
+ $Y2=2.3
cc_776 N_CK_c_961_n N_A_704_89#_c_1351_n 0.00436024f $X=5.405 $Y=1.85 $X2=5.345
+ $Y2=2.3
cc_777 N_CK_c_948_n N_A_704_89#_c_1352_n 0.0220721f $X=5.405 $Y=1.85 $X2=5.885
+ $Y2=1.85
cc_778 N_CK_c_952_n N_A_704_89#_c_1352_n 0.00227671f $X=5.885 $Y=2.765 $X2=5.885
+ $Y2=1.85
cc_779 N_CK_c_961_n N_A_704_89#_c_1352_n 0.00131283f $X=5.405 $Y=1.85 $X2=5.885
+ $Y2=1.85
cc_780 N_CK_c_966_n N_A_704_89#_c_1352_n 5.27321e-19 $X=5.885 $Y=2.59 $X2=5.885
+ $Y2=1.85
cc_781 N_CK_c_970_n N_A_704_89#_c_1352_n 8.78837e-19 $X=6.03 $Y=2.59 $X2=5.885
+ $Y2=1.85
cc_782 N_CK_c_949_n N_A_704_89#_c_1353_n 0.0268981f $X=5.405 $Y=1.685 $X2=5.885
+ $Y2=1.685
cc_783 N_CK_c_942_n N_A_704_89#_c_1356_n 0.00592387f $X=6.79 $Y=2.6 $X2=6.865
+ $Y2=1.85
cc_784 N_CK_c_948_n N_A_704_89#_c_1356_n 8.05876e-19 $X=5.405 $Y=1.85 $X2=6.865
+ $Y2=1.85
cc_785 N_CK_c_952_n N_A_704_89#_c_1356_n 5.56676e-19 $X=5.885 $Y=2.765 $X2=6.865
+ $Y2=1.85
cc_786 N_CK_c_958_n N_A_704_89#_c_1356_n 0.00762848f $X=6.762 $Y=1.835 $X2=6.865
+ $Y2=1.85
cc_787 N_CK_c_961_n N_A_704_89#_c_1356_n 0.00853323f $X=5.405 $Y=1.85 $X2=6.865
+ $Y2=1.85
cc_788 N_CK_c_962_n N_A_704_89#_c_1356_n 0.00132011f $X=5.8 $Y=2.59 $X2=6.865
+ $Y2=1.85
cc_789 N_CK_c_964_n N_A_704_89#_c_1356_n 8.24249e-19 $X=6.88 $Y=2.59 $X2=6.865
+ $Y2=1.85
cc_790 N_CK_c_966_n N_A_704_89#_c_1356_n 0.00261697f $X=5.885 $Y=2.59 $X2=6.865
+ $Y2=1.85
cc_791 N_CK_c_967_n N_A_704_89#_c_1356_n 3.12599e-19 $X=5.74 $Y=2.59 $X2=6.865
+ $Y2=1.85
cc_792 N_CK_c_969_n N_A_704_89#_c_1356_n 0.00341454f $X=6.735 $Y=2.59 $X2=6.865
+ $Y2=1.85
cc_793 N_CK_c_970_n N_A_704_89#_c_1356_n 0.00221563f $X=6.03 $Y=2.59 $X2=6.865
+ $Y2=1.85
cc_794 N_CK_c_953_n N_A_704_89#_c_1358_n 0.0102351f $X=6.762 $Y=1.685 $X2=6.95
+ $Y2=0.825
cc_795 N_CK_c_958_n N_A_704_89#_c_1358_n 0.00243671f $X=6.762 $Y=1.835 $X2=6.95
+ $Y2=0.825
cc_796 N_CK_c_942_n N_A_704_89#_c_1363_n 0.00495963f $X=6.79 $Y=2.6 $X2=6.95
+ $Y2=2.105
cc_797 N_CK_c_941_n N_A_704_89#_c_1364_n 0.00262756f $X=6.735 $Y=2.93 $X2=7.22
+ $Y2=3.1
cc_798 N_CK_M1012_g N_A_704_89#_c_1364_n 0.00395773f $X=6.735 $Y=4.585 $X2=7.22
+ $Y2=3.1
cc_799 N_CK_c_942_n N_A_704_89#_c_1364_n 0.0049943f $X=6.79 $Y=2.6 $X2=7.22
+ $Y2=3.1
cc_800 N_CK_c_964_n N_A_704_89#_c_1364_n 0.0285927f $X=6.88 $Y=2.59 $X2=7.22
+ $Y2=3.1
cc_801 CK N_A_704_89#_c_1364_n 0.00851352f $X=6.88 $Y=2.59 $X2=7.22 $Y2=3.1
cc_802 N_CK_c_942_n N_A_704_89#_c_1365_n 0.00126782f $X=6.79 $Y=2.6 $X2=6.95
+ $Y2=1.85
cc_803 N_CK_c_958_n N_A_704_89#_c_1365_n 8.92648e-19 $X=6.762 $Y=1.835 $X2=6.95
+ $Y2=1.85
cc_804 N_CK_c_941_n N_A_704_89#_c_1366_n 0.001573f $X=6.735 $Y=2.93 $X2=7.22
+ $Y2=2.19
cc_805 N_CK_c_942_n N_A_704_89#_c_1366_n 0.00236123f $X=6.79 $Y=2.6 $X2=7.22
+ $Y2=2.19
cc_806 N_CK_c_964_n N_A_704_89#_c_1366_n 0.00528683f $X=6.88 $Y=2.59 $X2=7.22
+ $Y2=2.19
cc_807 CK N_A_704_89#_c_1366_n 8.7939e-19 $X=6.88 $Y=2.59 $X2=7.22 $Y2=2.19
cc_808 N_CK_c_941_n N_A_704_89#_c_1377_n 0.00233394f $X=6.735 $Y=2.93 $X2=7.22
+ $Y2=3.185
cc_809 N_CK_c_964_n N_A_704_89#_c_1377_n 0.00601935f $X=6.88 $Y=2.59 $X2=7.22
+ $Y2=3.185
cc_810 N_CK_c_942_n N_A_1246_89#_M1006_g 0.00697006f $X=6.79 $Y=2.6 $X2=6.305
+ $Y2=1.075
cc_811 N_CK_c_953_n N_A_1246_89#_M1006_g 0.0287519f $X=6.762 $Y=1.685 $X2=6.305
+ $Y2=1.075
cc_812 N_CK_c_941_n N_A_1246_89#_M1009_g 0.02899f $X=6.735 $Y=2.93 $X2=6.305
+ $Y2=4.585
cc_813 N_CK_c_942_n N_A_1246_89#_M1009_g 0.0175925f $X=6.79 $Y=2.6 $X2=6.305
+ $Y2=4.585
cc_814 N_CK_c_952_n N_A_1246_89#_M1009_g 0.215582f $X=5.885 $Y=2.765 $X2=6.305
+ $Y2=4.585
cc_815 N_CK_c_964_n N_A_1246_89#_M1009_g 0.00276527f $X=6.88 $Y=2.59 $X2=6.305
+ $Y2=4.585
cc_816 N_CK_c_966_n N_A_1246_89#_M1009_g 0.00472186f $X=5.885 $Y=2.59 $X2=6.305
+ $Y2=4.585
cc_817 N_CK_c_969_n N_A_1246_89#_M1009_g 0.00672311f $X=6.735 $Y=2.59 $X2=6.305
+ $Y2=4.585
cc_818 N_CK_c_970_n N_A_1246_89#_M1009_g 0.00113587f $X=6.03 $Y=2.59 $X2=6.305
+ $Y2=4.585
cc_819 CK N_A_1246_89#_M1009_g 3.05655e-19 $X=6.88 $Y=2.59 $X2=6.305 $Y2=4.585
cc_820 N_CK_c_942_n N_A_1246_89#_c_1539_n 0.0213817f $X=6.79 $Y=2.6 $X2=6.365
+ $Y2=2.19
cc_821 N_CK_c_969_n N_A_1246_89#_c_1539_n 0.00185875f $X=6.735 $Y=2.59 $X2=6.365
+ $Y2=2.19
cc_822 N_CK_c_942_n N_A_1246_89#_c_1545_n 8.95026e-19 $X=6.79 $Y=2.6 $X2=6.365
+ $Y2=2.19
cc_823 N_CK_c_969_n N_A_1246_89#_c_1545_n 0.00488871f $X=6.735 $Y=2.59 $X2=6.365
+ $Y2=2.19
cc_824 N_CK_c_941_n N_A_1246_89#_c_1552_n 2.34467e-19 $X=6.735 $Y=2.93 $X2=9.235
+ $Y2=2.19
cc_825 N_CK_c_942_n N_A_1246_89#_c_1552_n 0.0033485f $X=6.79 $Y=2.6 $X2=9.235
+ $Y2=2.19
cc_826 N_CK_c_964_n N_A_1246_89#_c_1552_n 8.38639e-19 $X=6.88 $Y=2.59 $X2=9.235
+ $Y2=2.19
cc_827 N_CK_c_969_n N_A_1246_89#_c_1552_n 0.0179446f $X=6.735 $Y=2.59 $X2=9.235
+ $Y2=2.19
cc_828 CK N_A_1246_89#_c_1552_n 0.0248956f $X=6.88 $Y=2.59 $X2=9.235 $Y2=2.19
cc_829 N_CK_c_942_n N_A_1246_89#_c_1553_n 8.66236e-19 $X=6.79 $Y=2.6 $X2=6.51
+ $Y2=2.19
cc_830 N_CK_c_969_n N_A_1246_89#_c_1553_n 0.0247156f $X=6.735 $Y=2.59 $X2=6.51
+ $Y2=2.19
cc_831 N_CK_c_941_n N_A_1084_115#_c_1705_n 0.00744372f $X=6.735 $Y=2.93
+ $X2=7.505 $Y2=2.63
cc_832 N_CK_c_942_n N_A_1084_115#_c_1705_n 0.00688829f $X=6.79 $Y=2.6 $X2=7.505
+ $Y2=2.63
cc_833 N_CK_c_941_n N_A_1084_115#_M1014_g 5.00344e-19 $X=6.735 $Y=2.93 $X2=7.685
+ $Y2=4.585
cc_834 N_CK_c_958_n N_A_1084_115#_c_1710_n 0.00688829f $X=6.762 $Y=1.835
+ $X2=7.685 $Y2=1.77
cc_835 N_CK_c_949_n N_A_1084_115#_c_1713_n 0.00554221f $X=5.405 $Y=1.685
+ $X2=5.065 $Y2=1.85
cc_836 N_CK_c_961_n N_A_1084_115#_c_1713_n 0.057541f $X=5.405 $Y=1.85 $X2=5.065
+ $Y2=1.85
cc_837 N_CK_c_963_n N_A_1084_115#_c_1713_n 0.0116326f $X=5.49 $Y=2.59 $X2=5.065
+ $Y2=1.85
cc_838 N_CK_c_966_n N_A_1084_115#_c_1713_n 0.00539276f $X=5.885 $Y=2.59
+ $X2=5.065 $Y2=1.85
cc_839 N_CK_c_967_n N_A_1084_115#_c_1713_n 0.0139004f $X=5.74 $Y=2.59 $X2=5.065
+ $Y2=1.85
cc_840 N_CK_c_970_n N_A_1084_115#_c_1713_n 6.61118e-19 $X=6.03 $Y=2.59 $X2=5.065
+ $Y2=1.85
cc_841 N_CK_c_948_n N_A_1084_115#_c_1738_n 0.00227744f $X=5.405 $Y=1.85
+ $X2=5.475 $Y2=1.43
cc_842 N_CK_c_949_n N_A_1084_115#_c_1738_n 0.0149609f $X=5.405 $Y=1.685
+ $X2=5.475 $Y2=1.43
cc_843 N_CK_c_961_n N_A_1084_115#_c_1738_n 0.0103267f $X=5.405 $Y=1.85 $X2=5.475
+ $Y2=1.43
cc_844 N_CK_c_952_n N_A_1084_115#_c_1757_n 0.00123101f $X=5.885 $Y=2.765
+ $X2=5.475 $Y2=3.185
cc_845 N_CK_c_962_n N_A_1084_115#_c_1757_n 0.00729874f $X=5.8 $Y=2.59 $X2=5.475
+ $Y2=3.185
cc_846 N_CK_c_963_n N_A_1084_115#_c_1757_n 0.00292714f $X=5.49 $Y=2.59 $X2=5.475
+ $Y2=3.185
cc_847 N_CK_c_966_n N_A_1084_115#_c_1757_n 8.86954e-19 $X=5.885 $Y=2.59
+ $X2=5.475 $Y2=3.185
cc_848 N_CK_c_942_n N_A_1084_115#_c_1717_n 2.89967e-19 $X=6.79 $Y=2.6 $X2=7.595
+ $Y2=1.85
cc_849 N_CK_c_958_n N_A_1084_115#_c_1717_n 2.26851e-19 $X=6.762 $Y=1.835
+ $X2=7.595 $Y2=1.85
cc_850 N_CK_c_942_n N_A_1084_115#_c_1719_n 0.00128484f $X=6.79 $Y=2.6 $X2=7.45
+ $Y2=1.85
cc_851 N_CK_c_948_n N_A_1084_115#_c_1719_n 0.00362401f $X=5.405 $Y=1.85 $X2=7.45
+ $Y2=1.85
cc_852 N_CK_c_958_n N_A_1084_115#_c_1719_n 0.00179204f $X=6.762 $Y=1.835
+ $X2=7.45 $Y2=1.85
cc_853 N_CK_c_961_n N_A_1084_115#_c_1719_n 0.0127028f $X=5.405 $Y=1.85 $X2=7.45
+ $Y2=1.85
cc_854 N_CK_c_962_n N_A_1084_115#_c_1719_n 0.00451177f $X=5.8 $Y=2.59 $X2=7.45
+ $Y2=1.85
cc_855 N_CK_c_966_n N_A_1084_115#_c_1719_n 6.39375e-19 $X=5.885 $Y=2.59 $X2=7.45
+ $Y2=1.85
cc_856 N_CK_c_970_n N_A_1084_115#_c_1719_n 0.0144351f $X=6.03 $Y=2.59 $X2=7.45
+ $Y2=1.85
cc_857 N_CK_c_948_n N_A_1084_115#_c_1722_n 9.79344e-19 $X=5.405 $Y=1.85 $X2=5.21
+ $Y2=1.85
cc_858 N_CK_c_961_n N_A_1084_115#_c_1722_n 0.00180575f $X=5.405 $Y=1.85 $X2=5.21
+ $Y2=1.85
cc_859 N_CK_c_967_n N_A_1084_115#_c_1722_n 0.0128239f $X=5.74 $Y=2.59 $X2=5.21
+ $Y2=1.85
cc_860 N_A_217_617#_c_1196_n N_A_704_89#_c_1341_n 0.00253253f $X=4.49 $Y=1.85
+ $X2=3.715 $Y2=2.225
cc_861 N_A_217_617#_c_1196_n N_A_704_89#_c_1342_n 0.00296105f $X=4.49 $Y=1.85
+ $X2=4.12 $Y2=2.3
cc_862 N_A_217_617#_c_1182_n N_A_704_89#_M1031_g 0.215934f $X=4.63 $Y=2.765
+ $X2=4.195 $Y2=4.585
cc_863 N_A_217_617#_c_1193_n N_A_704_89#_M1031_g 0.00493295f $X=4.725 $Y=2.765
+ $X2=4.195 $Y2=4.585
cc_864 N_A_217_617#_c_1180_n N_A_704_89#_c_1345_n 0.0342351f $X=4.63 $Y=1.85
+ $X2=5.27 $Y2=2.3
cc_865 N_A_217_617#_c_1182_n N_A_704_89#_c_1345_n 0.0307748f $X=4.63 $Y=2.765
+ $X2=5.27 $Y2=2.3
cc_866 N_A_217_617#_c_1193_n N_A_704_89#_c_1345_n 0.0113171f $X=4.725 $Y=2.765
+ $X2=5.27 $Y2=2.3
cc_867 N_A_217_617#_c_1194_n N_A_704_89#_c_1345_n 8.69982e-19 $X=4.725 $Y=1.85
+ $X2=5.27 $Y2=2.3
cc_868 N_A_217_617#_c_1196_n N_A_704_89#_c_1345_n 0.00486036f $X=4.49 $Y=1.85
+ $X2=5.27 $Y2=2.3
cc_869 N_A_217_617#_c_1247_n N_A_704_89#_c_1345_n 4.12801e-19 $X=4.635 $Y=1.85
+ $X2=5.27 $Y2=2.3
cc_870 N_A_217_617#_c_1181_n N_A_704_89#_M1025_g 0.21333f $X=4.91 $Y=2.765
+ $X2=5.345 $Y2=4.585
cc_871 N_A_217_617#_M1021_g N_A_1084_115#_c_1713_n 0.001069f $X=4.555 $Y=1.075
+ $X2=5.065 $Y2=1.85
cc_872 N_A_217_617#_M1024_g N_A_1084_115#_c_1713_n 0.0012608f $X=4.555 $Y=4.585
+ $X2=5.065 $Y2=1.85
cc_873 N_A_217_617#_c_1178_n N_A_1084_115#_c_1713_n 0.0061959f $X=4.91 $Y=1.85
+ $X2=5.065 $Y2=1.85
cc_874 N_A_217_617#_c_1181_n N_A_1084_115#_c_1713_n 0.00723389f $X=4.91 $Y=2.765
+ $X2=5.065 $Y2=1.85
cc_875 N_A_217_617#_M1026_g N_A_1084_115#_c_1713_n 0.00502021f $X=4.985 $Y=1.075
+ $X2=5.065 $Y2=1.85
cc_876 N_A_217_617#_M1027_g N_A_1084_115#_c_1713_n 0.0051844f $X=4.985 $Y=4.585
+ $X2=5.065 $Y2=1.85
cc_877 N_A_217_617#_c_1193_n N_A_1084_115#_c_1713_n 0.0700853f $X=4.725 $Y=2.765
+ $X2=5.065 $Y2=1.85
cc_878 N_A_217_617#_c_1194_n N_A_1084_115#_c_1713_n 0.0157315f $X=4.725 $Y=1.85
+ $X2=5.065 $Y2=1.85
cc_879 N_A_217_617#_c_1247_n N_A_1084_115#_c_1713_n 4.18442e-19 $X=4.635 $Y=1.85
+ $X2=5.065 $Y2=1.85
cc_880 N_A_217_617#_M1021_g N_A_1084_115#_c_1739_n 0.00136315f $X=4.555 $Y=1.075
+ $X2=5.15 $Y2=1.43
cc_881 N_A_217_617#_M1026_g N_A_1084_115#_c_1739_n 0.0099627f $X=4.985 $Y=1.075
+ $X2=5.15 $Y2=1.43
cc_882 N_A_217_617#_M1024_g N_A_1084_115#_c_1805_n 9.13132e-19 $X=4.555 $Y=4.585
+ $X2=5.15 $Y2=3.185
cc_883 N_A_217_617#_M1027_g N_A_1084_115#_c_1805_n 0.0096885f $X=4.985 $Y=4.585
+ $X2=5.15 $Y2=3.185
cc_884 N_A_217_617#_c_1178_n N_A_1084_115#_c_1722_n 0.00229064f $X=4.91 $Y=1.85
+ $X2=5.21 $Y2=1.85
cc_885 N_A_217_617#_c_1194_n N_A_1084_115#_c_1722_n 0.0012094f $X=4.725 $Y=1.85
+ $X2=5.21 $Y2=1.85
cc_886 N_A_217_617#_c_1247_n N_A_1084_115#_c_1722_n 0.0241863f $X=4.635 $Y=1.85
+ $X2=5.21 $Y2=1.85
cc_887 N_A_704_89#_c_1348_n N_A_1246_89#_M1006_g 0.0073696f $X=5.825 $Y=2.225
+ $X2=6.305 $Y2=1.075
cc_888 N_A_704_89#_c_1353_n N_A_1246_89#_M1006_g 0.0974852f $X=5.885 $Y=1.685
+ $X2=6.305 $Y2=1.075
cc_889 N_A_704_89#_c_1356_n N_A_1246_89#_M1006_g 0.0107575f $X=6.865 $Y=1.85
+ $X2=6.305 $Y2=1.075
cc_890 N_A_704_89#_c_1347_n N_A_1246_89#_c_1539_n 0.0073696f $X=5.75 $Y=2.3
+ $X2=6.365 $Y2=2.19
cc_891 N_A_704_89#_c_1356_n N_A_1246_89#_c_1539_n 0.00290516f $X=6.865 $Y=1.85
+ $X2=6.365 $Y2=2.19
cc_892 N_A_704_89#_c_1366_n N_A_1246_89#_c_1539_n 2.96928e-19 $X=7.22 $Y=2.19
+ $X2=6.365 $Y2=2.19
cc_893 N_A_704_89#_c_1348_n N_A_1246_89#_c_1545_n 0.0035305f $X=5.825 $Y=2.225
+ $X2=6.365 $Y2=2.19
cc_894 N_A_704_89#_c_1356_n N_A_1246_89#_c_1545_n 0.0219931f $X=6.865 $Y=1.85
+ $X2=6.365 $Y2=2.19
cc_895 N_A_704_89#_c_1366_n N_A_1246_89#_c_1545_n 0.00559532f $X=7.22 $Y=2.19
+ $X2=6.365 $Y2=2.19
cc_896 N_A_704_89#_c_1356_n N_A_1246_89#_c_1552_n 0.00314603f $X=6.865 $Y=1.85
+ $X2=9.235 $Y2=2.19
cc_897 N_A_704_89#_c_1363_n N_A_1246_89#_c_1552_n 6.94255e-19 $X=6.95 $Y=2.105
+ $X2=9.235 $Y2=2.19
cc_898 N_A_704_89#_c_1364_n N_A_1246_89#_c_1552_n 0.00464833f $X=7.22 $Y=3.1
+ $X2=9.235 $Y2=2.19
cc_899 N_A_704_89#_c_1366_n N_A_1246_89#_c_1552_n 0.0207528f $X=7.22 $Y=2.19
+ $X2=9.235 $Y2=2.19
cc_900 N_A_704_89#_c_1348_n N_A_1246_89#_c_1553_n 9.14174e-19 $X=5.825 $Y=2.225
+ $X2=6.51 $Y2=2.19
cc_901 N_A_704_89#_c_1356_n N_A_1246_89#_c_1553_n 0.0010261f $X=6.865 $Y=1.85
+ $X2=6.51 $Y2=2.19
cc_902 N_A_704_89#_c_1363_n N_A_1246_89#_c_1553_n 0.00122156f $X=6.95 $Y=2.105
+ $X2=6.51 $Y2=2.19
cc_903 N_A_704_89#_c_1363_n N_A_1084_115#_c_1705_n 0.00130229f $X=6.95 $Y=2.105
+ $X2=7.505 $Y2=2.63
cc_904 N_A_704_89#_c_1364_n N_A_1084_115#_c_1705_n 0.00568165f $X=7.22 $Y=3.1
+ $X2=7.505 $Y2=2.63
cc_905 N_A_704_89#_c_1366_n N_A_1084_115#_c_1705_n 0.00134862f $X=7.22 $Y=2.19
+ $X2=7.505 $Y2=2.63
cc_906 N_A_704_89#_c_1358_n N_A_1084_115#_c_1706_n 0.00649036f $X=6.95 $Y=0.825
+ $X2=7.685 $Y2=1.69
cc_907 N_A_704_89#_c_1373_n N_A_1084_115#_M1014_g 0.00664364f $X=6.95 $Y=3.455
+ $X2=7.685 $Y2=4.585
cc_908 N_A_704_89#_c_1364_n N_A_1084_115#_M1014_g 0.00331798f $X=7.22 $Y=3.1
+ $X2=7.685 $Y2=4.585
cc_909 N_A_704_89#_c_1377_n N_A_1084_115#_M1014_g 0.00560488f $X=7.22 $Y=3.185
+ $X2=7.685 $Y2=4.585
cc_910 N_A_704_89#_c_1358_n N_A_1084_115#_c_1710_n 0.00137598f $X=6.95 $Y=0.825
+ $X2=7.685 $Y2=1.77
cc_911 N_A_704_89#_c_1365_n N_A_1084_115#_c_1710_n 9.86466e-19 $X=6.95 $Y=1.85
+ $X2=7.685 $Y2=1.77
cc_912 N_A_704_89#_c_1345_n N_A_1084_115#_c_1713_n 0.0124213f $X=5.27 $Y=2.3
+ $X2=5.065 $Y2=1.85
cc_913 N_A_704_89#_M1025_g N_A_1084_115#_c_1713_n 0.0105859f $X=5.345 $Y=4.585
+ $X2=5.065 $Y2=1.85
cc_914 N_A_704_89#_c_1352_n N_A_1084_115#_c_1738_n 0.00174784f $X=5.885 $Y=1.85
+ $X2=5.475 $Y2=1.43
cc_915 N_A_704_89#_c_1353_n N_A_1084_115#_c_1738_n 0.00205316f $X=5.885 $Y=1.685
+ $X2=5.475 $Y2=1.43
cc_916 N_A_704_89#_c_1356_n N_A_1084_115#_c_1738_n 0.00436807f $X=6.865 $Y=1.85
+ $X2=5.475 $Y2=1.43
cc_917 N_A_704_89#_M1025_g N_A_1084_115#_c_1757_n 0.0157833f $X=5.345 $Y=4.585
+ $X2=5.475 $Y2=3.185
cc_918 N_A_704_89#_c_1363_n N_A_1084_115#_c_1717_n 0.00520507f $X=6.95 $Y=2.105
+ $X2=7.595 $Y2=1.85
cc_919 N_A_704_89#_c_1364_n N_A_1084_115#_c_1717_n 0.039533f $X=7.22 $Y=3.1
+ $X2=7.595 $Y2=1.85
cc_920 N_A_704_89#_c_1365_n N_A_1084_115#_c_1717_n 0.00358095f $X=6.95 $Y=1.85
+ $X2=7.595 $Y2=1.85
cc_921 N_A_704_89#_c_1366_n N_A_1084_115#_c_1717_n 0.00955403f $X=7.22 $Y=2.19
+ $X2=7.595 $Y2=1.85
cc_922 N_A_704_89#_c_1345_n N_A_1084_115#_c_1719_n 0.00156696f $X=5.27 $Y=2.3
+ $X2=7.45 $Y2=1.85
cc_923 N_A_704_89#_c_1347_n N_A_1084_115#_c_1719_n 0.00244106f $X=5.75 $Y=2.3
+ $X2=7.45 $Y2=1.85
cc_924 N_A_704_89#_c_1351_n N_A_1084_115#_c_1719_n 5.19983e-19 $X=5.345 $Y=2.3
+ $X2=7.45 $Y2=1.85
cc_925 N_A_704_89#_c_1352_n N_A_1084_115#_c_1719_n 0.00455939f $X=5.885 $Y=1.85
+ $X2=7.45 $Y2=1.85
cc_926 N_A_704_89#_c_1356_n N_A_1084_115#_c_1719_n 0.0492477f $X=6.865 $Y=1.85
+ $X2=7.45 $Y2=1.85
cc_927 N_A_704_89#_c_1365_n N_A_1084_115#_c_1719_n 0.0117855f $X=6.95 $Y=1.85
+ $X2=7.45 $Y2=1.85
cc_928 N_A_704_89#_c_1366_n N_A_1084_115#_c_1719_n 0.00219678f $X=7.22 $Y=2.19
+ $X2=7.45 $Y2=1.85
cc_929 N_A_704_89#_c_1345_n N_A_1084_115#_c_1722_n 0.00120486f $X=5.27 $Y=2.3
+ $X2=5.21 $Y2=1.85
cc_930 N_A_704_89#_c_1358_n N_A_1084_115#_c_1723_n 0.0010241f $X=6.95 $Y=0.825
+ $X2=7.595 $Y2=1.85
cc_931 N_A_704_89#_c_1363_n N_A_1084_115#_c_1723_n 6.33705e-19 $X=6.95 $Y=2.105
+ $X2=7.595 $Y2=1.85
cc_932 N_A_704_89#_c_1373_n N_A_1469_617#_c_1970_n 0.101221f $X=6.95 $Y=3.455
+ $X2=7.47 $Y2=3.795
cc_933 N_A_704_89#_c_1373_n N_A_1469_617#_c_1982_n 0.00811594f $X=6.95 $Y=3.455
+ $X2=7.555 $Y2=3.63
cc_934 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1705_n 0.00586968f $X=9.235 $Y=2.19
+ $X2=7.505 $Y2=2.63
cc_935 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1710_n 6.8924e-19 $X=9.235 $Y=2.19
+ $X2=7.685 $Y2=1.77
cc_936 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1712_n 0.00207076f $X=9.235 $Y=2.19
+ $X2=7.685 $Y2=2.765
cc_937 N_A_1246_89#_c_1546_n N_A_1084_115#_c_1717_n 0.0010677f $X=8.26 $Y=0.825
+ $X2=7.595 $Y2=1.85
cc_938 N_A_1246_89#_c_1550_n N_A_1084_115#_c_1717_n 0.00422342f $X=8.845 $Y=2.19
+ $X2=7.595 $Y2=1.85
cc_939 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1717_n 0.0169834f $X=9.235 $Y=2.19
+ $X2=7.595 $Y2=1.85
cc_940 N_A_1246_89#_M1006_g N_A_1084_115#_c_1719_n 0.00231271f $X=6.305 $Y=1.075
+ $X2=7.45 $Y2=1.85
cc_941 N_A_1246_89#_c_1539_n N_A_1084_115#_c_1719_n 0.00187603f $X=6.365 $Y=2.19
+ $X2=7.45 $Y2=1.85
cc_942 N_A_1246_89#_c_1545_n N_A_1084_115#_c_1719_n 0.00166223f $X=6.365 $Y=2.19
+ $X2=7.45 $Y2=1.85
cc_943 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1719_n 0.0841111f $X=9.235 $Y=2.19
+ $X2=7.45 $Y2=1.85
cc_944 N_A_1246_89#_c_1553_n N_A_1084_115#_c_1719_n 0.0289631f $X=6.51 $Y=2.19
+ $X2=7.45 $Y2=1.85
cc_945 N_A_1246_89#_c_1546_n N_A_1084_115#_c_1723_n 0.00247064f $X=8.26 $Y=0.825
+ $X2=7.595 $Y2=1.85
cc_946 N_A_1246_89#_c_1550_n N_A_1084_115#_c_1723_n 0.00385422f $X=8.845 $Y=2.19
+ $X2=7.595 $Y2=1.85
cc_947 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1723_n 0.027605f $X=9.235 $Y=2.19
+ $X2=7.595 $Y2=1.85
cc_948 N_A_1246_89#_M1007_g N_QN_M1010_g 0.0391431f $X=9.495 $Y=0.945 $X2=9.925
+ $Y2=0.945
cc_949 N_A_1246_89#_c_1541_n N_QN_M1010_g 0.0153129f $X=9.382 $Y=2.025 $X2=9.925
+ $Y2=0.945
cc_950 N_A_1246_89#_c_1551_n N_QN_M1010_g 4.79563e-19 $X=9.38 $Y=2.19 $X2=9.925
+ $Y2=0.945
cc_951 N_A_1246_89#_c_1543_n N_QN_M1029_g 0.0102953f $X=9.47 $Y=2.855 $X2=9.925
+ $Y2=5.085
cc_952 N_A_1246_89#_c_1544_n N_QN_M1029_g 0.0662174f $X=9.47 $Y=3.005 $X2=9.925
+ $Y2=5.085
cc_953 N_A_1246_89#_c_1540_n N_QN_c_1866_n 0.021196f $X=9.38 $Y=2.19 $X2=9.865
+ $Y2=2.395
cc_954 N_A_1246_89#_c_1551_n N_QN_c_1866_n 3.0115e-19 $X=9.38 $Y=2.19 $X2=9.865
+ $Y2=2.395
cc_955 N_A_1246_89#_c_1554_n N_QN_c_1866_n 4.60229e-19 $X=9.38 $Y=2.19 $X2=9.865
+ $Y2=2.395
cc_956 N_A_1246_89#_M1007_g N_QN_c_1867_n 0.016723f $X=9.495 $Y=0.945 $X2=9.28
+ $Y2=0.825
cc_957 N_A_1246_89#_c_1542_n N_QN_c_1867_n 0.00312124f $X=9.47 $Y=1.8 $X2=9.28
+ $Y2=0.825
cc_958 N_A_1246_89#_M1028_g N_QN_c_1871_n 0.0462756f $X=9.495 $Y=5.085 $X2=9.28
+ $Y2=2.96
cc_959 N_A_1246_89#_c_1543_n N_QN_c_1871_n 0.00516467f $X=9.47 $Y=2.855 $X2=9.28
+ $Y2=2.96
cc_960 N_A_1246_89#_c_1549_n N_QN_c_1871_n 0.136786f $X=8.76 $Y=3.795 $X2=9.28
+ $Y2=2.96
cc_961 N_A_1246_89#_c_1541_n N_QN_c_1872_n 0.00722072f $X=9.382 $Y=2.025
+ $X2=9.78 $Y2=1.85
cc_962 N_A_1246_89#_c_1542_n N_QN_c_1872_n 0.0108332f $X=9.47 $Y=1.8 $X2=9.78
+ $Y2=1.85
cc_963 N_A_1246_89#_c_1551_n N_QN_c_1872_n 0.0110498f $X=9.38 $Y=2.19 $X2=9.78
+ $Y2=1.85
cc_964 N_A_1246_89#_c_1554_n N_QN_c_1872_n 0.00387586f $X=9.38 $Y=2.19 $X2=9.78
+ $Y2=1.85
cc_965 N_A_1246_89#_c_1540_n N_QN_c_1873_n 0.00308111f $X=9.38 $Y=2.19 $X2=9.365
+ $Y2=1.85
cc_966 N_A_1246_89#_c_1550_n N_QN_c_1873_n 0.00372477f $X=8.845 $Y=2.19
+ $X2=9.365 $Y2=1.85
cc_967 N_A_1246_89#_c_1551_n N_QN_c_1873_n 0.0120703f $X=9.38 $Y=2.19 $X2=9.365
+ $Y2=1.85
cc_968 N_A_1246_89#_c_1552_n N_QN_c_1873_n 0.0010572f $X=9.235 $Y=2.19 $X2=9.365
+ $Y2=1.85
cc_969 N_A_1246_89#_c_1554_n N_QN_c_1873_n 0.00336135f $X=9.38 $Y=2.19 $X2=9.365
+ $Y2=1.85
cc_970 N_A_1246_89#_c_1543_n N_QN_c_1874_n 0.0151488f $X=9.47 $Y=2.855 $X2=9.78
+ $Y2=2.765
cc_971 N_A_1246_89#_c_1544_n N_QN_c_1874_n 0.00248624f $X=9.47 $Y=3.005 $X2=9.78
+ $Y2=2.765
cc_972 N_A_1246_89#_c_1551_n N_QN_c_1874_n 0.00426371f $X=9.38 $Y=2.19 $X2=9.78
+ $Y2=2.765
cc_973 N_A_1246_89#_c_1554_n N_QN_c_1874_n 0.00253233f $X=9.38 $Y=2.19 $X2=9.78
+ $Y2=2.765
cc_974 N_A_1246_89#_c_1540_n N_QN_c_1875_n 0.00265611f $X=9.38 $Y=2.19 $X2=9.365
+ $Y2=2.765
cc_975 N_A_1246_89#_c_1549_n N_QN_c_1875_n 0.00792667f $X=8.76 $Y=3.795
+ $X2=9.365 $Y2=2.765
cc_976 N_A_1246_89#_c_1551_n N_QN_c_1875_n 0.00471962f $X=9.38 $Y=2.19 $X2=9.365
+ $Y2=2.765
cc_977 N_A_1246_89#_c_1552_n N_QN_c_1875_n 9.40773e-19 $X=9.235 $Y=2.19
+ $X2=9.365 $Y2=2.765
cc_978 N_A_1246_89#_c_1554_n N_QN_c_1875_n 0.00140341f $X=9.38 $Y=2.19 $X2=9.365
+ $Y2=2.765
cc_979 N_A_1246_89#_c_1540_n N_QN_c_1876_n 0.00216137f $X=9.38 $Y=2.19 $X2=9.865
+ $Y2=2.395
cc_980 N_A_1246_89#_c_1541_n N_QN_c_1876_n 0.00323473f $X=9.382 $Y=2.025
+ $X2=9.865 $Y2=2.395
cc_981 N_A_1246_89#_c_1543_n N_QN_c_1876_n 0.00226435f $X=9.47 $Y=2.855
+ $X2=9.865 $Y2=2.395
cc_982 N_A_1246_89#_c_1551_n N_QN_c_1876_n 0.00987106f $X=9.38 $Y=2.19 $X2=9.865
+ $Y2=2.395
cc_983 N_A_1246_89#_c_1554_n N_QN_c_1876_n 0.00377439f $X=9.38 $Y=2.19 $X2=9.865
+ $Y2=2.395
cc_984 N_A_1246_89#_M1028_g QN 0.00233857f $X=9.495 $Y=5.085 $X2=9.285 $Y2=2.96
cc_985 N_A_1246_89#_c_1544_n QN 0.00481276f $X=9.47 $Y=3.005 $X2=9.285 $Y2=2.96
cc_986 N_A_1246_89#_c_1549_n QN 0.00717706f $X=8.76 $Y=3.795 $X2=9.285 $Y2=2.96
cc_987 N_A_1246_89#_c_1551_n QN 0.00359685f $X=9.38 $Y=2.19 $X2=9.285 $Y2=2.96
cc_988 N_A_1246_89#_c_1554_n QN 0.00842298f $X=9.38 $Y=2.19 $X2=9.285 $Y2=2.96
cc_989 N_A_1246_89#_M1028_g Q 0.0011399f $X=9.495 $Y=5.085 $X2=10.135 $Y2=3.33
cc_990 N_A_1084_115#_c_1757_n A_1012_617# 0.00310684f $X=5.475 $Y=3.185 $X2=5.06
+ $Y2=3.085
cc_991 N_A_1084_115#_c_1805_n A_1012_617# 0.00144354f $X=5.15 $Y=3.185 $X2=5.06
+ $Y2=3.085
cc_992 N_A_1084_115#_M1014_g N_A_1469_617#_c_1973_n 0.0155681f $X=7.685 $Y=4.585
+ $X2=8.245 $Y2=3.63
cc_993 N_A_1084_115#_c_1717_n N_A_1469_617#_c_1973_n 0.00125278f $X=7.595
+ $Y=1.85 $X2=8.245 $Y2=3.63
cc_994 N_A_1084_115#_c_1712_n N_A_1469_617#_c_1982_n 0.0020255f $X=7.685
+ $Y=2.765 $X2=7.555 $Y2=3.63
cc_995 N_A_1084_115#_c_1717_n N_A_1469_617#_c_1982_n 7.57421e-19 $X=7.595
+ $Y=1.85 $X2=7.555 $Y2=3.63
cc_996 N_A_1084_115#_c_1713_n A_1012_115# 9.4749e-19 $X=5.065 $Y=1.85 $X2=5.06
+ $Y2=0.575
cc_997 N_A_1084_115#_c_1738_n A_1012_115# 0.00337089f $X=5.475 $Y=1.43 $X2=5.06
+ $Y2=0.575
cc_998 N_A_1084_115#_c_1739_n A_1012_115# 0.00148865f $X=5.15 $Y=1.43 $X2=5.06
+ $Y2=0.575
cc_999 N_QN_M1010_g N_Q_c_1989_n 0.011148f $X=9.925 $Y=0.945 $X2=10.14 $Y2=0.825
cc_1000 N_QN_M1029_g N_Q_c_1993_n 0.0305875f $X=9.925 $Y=5.085 $X2=10.14
+ $Y2=4.475
cc_1001 N_QN_M1010_g N_Q_c_1991_n 0.0383548f $X=9.925 $Y=0.945 $X2=10.255
+ $Y2=3.16
cc_1002 N_QN_c_1872_n N_Q_c_1991_n 0.0111776f $X=9.78 $Y=1.85 $X2=10.255
+ $Y2=3.16
cc_1003 N_QN_c_1874_n N_Q_c_1991_n 0.0111776f $X=9.78 $Y=2.765 $X2=10.255
+ $Y2=3.16
cc_1004 N_QN_c_1876_n N_Q_c_1991_n 0.0438362f $X=9.865 $Y=2.395 $X2=10.255
+ $Y2=3.16
cc_1005 N_QN_M1010_g N_Q_c_1992_n 0.00695117f $X=9.925 $Y=0.945 $X2=10.255
+ $Y2=1.515
cc_1006 N_QN_M1029_g N_Q_c_1997_n 0.00911548f $X=9.925 $Y=5.085 $X2=10.14
+ $Y2=3.287
cc_1007 N_QN_M1029_g Q 0.0145232f $X=9.925 $Y=5.085 $X2=10.135 $Y2=3.33
cc_1008 N_QN_c_1871_n Q 0.00553023f $X=9.28 $Y=2.96 $X2=10.135 $Y2=3.33
cc_1009 N_QN_c_1874_n Q 0.00245821f $X=9.78 $Y=2.765 $X2=10.135 $Y2=3.33
