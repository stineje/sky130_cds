magic
tech sky130A
magscale 1 2
timestamp 1604007754
<< checkpaint >>
rect -1269 2461 1439 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1439 -1129
<< nwell >>
rect -9 529 179 1119
<< locali >>
rect 0 1049 176 1110
rect 0 0 176 61
<< metal1 >>
rect 0 1049 176 1110
rect 0 0 176 61
<< labels >>
rlabel metal1 112 28 112 28 1 gnd
rlabel metal1 111 1081 111 1081 1 vdd
<< end >>
