* File: sky130_osu_sc_15T_ls__inv_8.pex.spice
* Created: Fri Nov 12 14:57:56 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__INV_8%GND 1 2 3 4 5 51 55 57 64 66 73 75 82 84
+ 92 104 106
r110 104 106 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.06 $Y2=0.152
r111 90 92 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.865
r112 85 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r113 84 90 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=3.615 $Y=0.152
+ $X2=3.7 $Y2=0.305
r114 80 100 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r115 80 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.865
r116 76 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r117 75 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r118 71 99 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r119 71 73 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.865
r120 67 98 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r121 66 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r122 62 98 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r123 62 64 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.865
r124 57 98 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r125 53 55 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r126 51 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=0.19
+ $X2=3.06 $Y2=0.19
r127 51 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r128 51 53 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r129 51 58 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r130 51 84 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r131 51 85 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r132 51 75 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r133 51 76 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r134 51 66 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r135 51 67 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r136 51 57 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r137 51 58 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r138 5 92 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.865
r139 4 82 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.865
r140 3 73 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.865
r141 2 64 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r142 1 55 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__INV_8%VDD 1 2 3 4 5 41 45 49 55 59 65 69 75 79
+ 86 97 101
r77 97 101 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=3.06 $Y2=5.397
r78 91 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r79 86 89 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.7 $Y=3.205
+ $X2=3.7 $Y2=4.565
r80 84 89 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=5.245 $X2=3.7
+ $Y2=4.565
r81 82 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=5.36
+ $X2=3.06 $Y2=5.36
r82 80 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=2.84 $Y2=5.397
r83 80 82 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=3.06 $Y2=5.397
r84 79 84 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.7 $Y2=5.245
r85 79 82 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.06 $Y2=5.397
r86 75 78 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.205
+ $X2=2.84 $Y2=4.565
r87 73 95 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=5.397
r88 73 78 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.565
r89 70 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r90 70 72 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r91 69 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.397
r92 69 72 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r93 65 68 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.205
+ $X2=1.98 $Y2=4.565
r94 63 94 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r95 63 68 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.565
r96 60 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r97 60 62 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r98 59 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r99 59 62 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r100 55 58 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=3.205
+ $X2=1.12 $Y2=4.565
r101 53 93 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r102 53 58 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r103 50 91 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r104 50 52 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r105 49 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r106 49 52 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r107 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r108 43 91 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r109 43 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r110 41 82 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r111 41 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r112 41 62 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r113 41 52 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r114 41 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r115 5 89 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=4.565
r116 5 86 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=3.205
r117 4 78 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.565
r118 4 75 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.205
r119 3 68 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.565
r120 3 65 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.205
r121 2 58 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r122 2 55 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.205
r123 1 48 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r124 1 45 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__INV_8%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 45 47 49 50 52 53 55 57 59 60 62 63 65 67 69
+ 70 72 73 75 77 79 80 82 83 85 86 88 89 90 91 92 93 94 95 96 97 98 99 100 103
+ 105 107 110
c234 70 0 1.33323e-19 $X=3.055 $Y=2.7
c235 67 0 1.33323e-19 $X=3.055 $Y=1.44
c236 60 0 1.33323e-19 $X=2.625 $Y=2.7
c237 57 0 1.33323e-19 $X=2.625 $Y=1.44
c238 50 0 1.33323e-19 $X=2.195 $Y=2.7
c239 45 0 1.33323e-19 $X=2.195 $Y=1.44
c240 38 0 1.33323e-19 $X=1.765 $Y=2.7
c241 35 0 1.33323e-19 $X=1.765 $Y=1.44
c242 28 0 1.33323e-19 $X=1.335 $Y=2.7
c243 25 0 1.33323e-19 $X=1.335 $Y=1.44
c244 18 0 1.33323e-19 $X=0.905 $Y=2.7
c245 15 0 1.33323e-19 $X=0.905 $Y=1.44
r246 110 113 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=3.065
+ $X2=0.405 $Y2=3.07
r247 105 107 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.045
+ $X2=0.535 $Y2=2.045
r248 103 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r249 101 105 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.405 $Y2=2.045
r250 101 103 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.32 $Y2=3.07
r251 85 107 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.045 $X2=0.535 $Y2=2.045
r252 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=2.21
r253 85 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=1.88
r254 80 82 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=3.825
r255 77 79 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.485 $Y2=0.945
r256 76 100 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.625
+ $X2=3.055 $Y2=2.625
r257 75 80 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.485 $Y2=2.7
r258 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.13 $Y2=2.625
r259 74 99 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.055 $Y2=1.515
r260 73 77 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.515
+ $X2=3.485 $Y2=1.44
r261 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.515
+ $X2=3.13 $Y2=1.515
r262 70 100 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=2.625
r263 70 72 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=3.825
r264 67 99 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=1.515
r265 67 69 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=0.945
r266 66 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.625
+ $X2=2.625 $Y2=2.625
r267 65 100 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=3.055 $Y2=2.625
r268 65 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=2.7 $Y2=2.625
r269 64 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.625 $Y2=1.515
r270 63 99 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=3.055 $Y2=1.515
r271 63 64 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=2.7 $Y2=1.515
r272 60 98 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=2.625
r273 60 62 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r274 57 97 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=1.515
r275 57 59 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=0.945
r276 56 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r277 55 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.625
r278 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r279 54 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.515
+ $X2=2.195 $Y2=1.515
r280 53 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.625 $Y2=1.515
r281 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.27 $Y2=1.515
r282 50 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7 $X2=2.195
+ $Y2=2.625
r283 50 52 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r284 49 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.55
+ $X2=2.195 $Y2=2.625
r285 48 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.59
+ $X2=2.195 $Y2=1.515
r286 48 49 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.59
+ $X2=2.195 $Y2=2.55
r287 45 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.44
+ $X2=2.195 $Y2=1.515
r288 45 47 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.195 $Y=1.44
+ $X2=2.195 $Y2=0.945
r289 44 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r290 43 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r291 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r292 42 93 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.515
+ $X2=1.765 $Y2=1.515
r293 41 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.515
+ $X2=2.195 $Y2=1.515
r294 41 42 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.515
+ $X2=1.84 $Y2=1.515
r295 38 94 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r296 38 40 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r297 35 93 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.44
+ $X2=1.765 $Y2=1.515
r298 35 37 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.765 $Y=1.44
+ $X2=1.765 $Y2=0.945
r299 34 92 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.625
+ $X2=1.335 $Y2=2.625
r300 33 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r301 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.41 $Y2=2.625
r302 32 91 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.335 $Y2=1.515
r303 31 93 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.765 $Y2=1.515
r304 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.41 $Y2=1.515
r305 28 92 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=2.625
r306 28 30 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r307 25 91 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.44
+ $X2=1.335 $Y2=1.515
r308 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.335 $Y=1.44
+ $X2=1.335 $Y2=0.945
r309 24 90 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.625
+ $X2=0.905 $Y2=2.625
r310 23 92 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.625
+ $X2=1.335 $Y2=2.625
r311 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.625
+ $X2=0.98 $Y2=2.625
r312 22 89 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.515
+ $X2=0.905 $Y2=1.515
r313 21 91 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=1.335 $Y2=1.515
r314 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=0.98 $Y2=1.515
r315 18 90 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.7
+ $X2=0.905 $Y2=2.625
r316 18 20 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=2.7
+ $X2=0.905 $Y2=3.825
r317 15 89 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.44
+ $X2=0.905 $Y2=1.515
r318 15 17 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.905 $Y=1.44
+ $X2=0.905 $Y2=0.945
r319 14 88 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.625
+ $X2=0.475 $Y2=2.625
r320 13 90 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.625
+ $X2=0.905 $Y2=2.625
r321 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.625
+ $X2=0.55 $Y2=2.625
r322 12 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.515
+ $X2=0.475 $Y2=1.515
r323 11 89 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.515
+ $X2=0.905 $Y2=1.515
r324 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.515
+ $X2=0.55 $Y2=1.515
r325 8 88 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.7
+ $X2=0.475 $Y2=2.625
r326 8 10 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.475 $Y=2.7
+ $X2=0.475 $Y2=3.825
r327 7 88 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.55
+ $X2=0.475 $Y2=2.625
r328 7 87 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.55
+ $X2=0.475 $Y2=2.21
r329 4 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.59
+ $X2=0.475 $Y2=1.515
r330 4 86 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.59
+ $X2=0.475 $Y2=1.88
r331 1 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=1.515
r332 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__INV_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68 76
+ 82 89 90 92 94 96 99 100 101 102 103 105 106 107 108 109 110 111
c171 111 0 1.33323e-19 $X=3.27 $Y=2.585
c172 110 0 1.33323e-19 $X=3.27 $Y=1.335
c173 109 0 2.66647e-19 $X=2.555 $Y=2.7
c174 107 0 2.66647e-19 $X=2.555 $Y=1.22
c175 103 0 2.66647e-19 $X=1.695 $Y=2.7
c176 101 0 2.66647e-19 $X=1.695 $Y=1.22
c177 90 0 1.33323e-19 $X=0.69 $Y=2.585
c178 89 0 1.33323e-19 $X=0.69 $Y=1.335
r179 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.585
+ $X2=3.27 $Y2=2.7
r180 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=1.22
r181 110 111 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=2.585
r182 109 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.7
+ $X2=2.41 $Y2=2.7
r183 108 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.7
+ $X2=3.27 $Y2=2.7
r184 108 109 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.7
+ $X2=2.555 $Y2=2.7
r185 107 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.22
+ $X2=2.41 $Y2=1.22
r186 106 125 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=3.27 $Y2=1.22
r187 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=2.555 $Y2=1.22
r188 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.585
+ $X2=2.41 $Y2=2.7
r189 104 121 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r190 104 105 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.585
r191 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.7
+ $X2=1.55 $Y2=2.7
r192 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.7
+ $X2=2.41 $Y2=2.7
r193 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.7
+ $X2=1.695 $Y2=2.7
r194 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r195 100 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r196 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r197 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.585
+ $X2=1.55 $Y2=2.7
r198 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r199 98 99 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=2.585
r200 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.7
+ $X2=0.69 $Y2=2.7
r201 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.7
+ $X2=1.55 $Y2=2.7
r202 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.7
+ $X2=0.835 $Y2=2.7
r203 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.22
+ $X2=0.69 $Y2=1.22
r204 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.22
+ $X2=1.55 $Y2=1.22
r205 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.22
+ $X2=0.835 $Y2=1.22
r206 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=2.7
r207 90 92 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=1.94
r208 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.22
r209 89 92 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.94
r210 85 87 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.27 $Y=3.205
+ $X2=3.27 $Y2=4.565
r211 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.7
+ $X2=3.27 $Y2=2.7
r212 82 85 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.27 $Y=2.7
+ $X2=3.27 $Y2=3.205
r213 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.22
+ $X2=3.27 $Y2=1.22
r214 76 79 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.27 $Y=0.865
+ $X2=3.27 $Y2=1.22
r215 71 73 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.205
+ $X2=2.41 $Y2=4.565
r216 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.7
+ $X2=2.41 $Y2=2.7
r217 68 71 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.41 $Y=2.7
+ $X2=2.41 $Y2=3.205
r218 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r219 62 65 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.41 $Y=0.865
+ $X2=2.41 $Y2=1.22
r220 57 59 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.205
+ $X2=1.55 $Y2=4.565
r221 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.7
+ $X2=1.55 $Y2=2.7
r222 54 57 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.55 $Y=2.7
+ $X2=1.55 $Y2=3.205
r223 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r224 48 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.55 $Y=0.865
+ $X2=1.55 $Y2=1.22
r225 43 45 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r226 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=2.7
r227 40 43 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=3.205
r228 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.22
+ $X2=0.69 $Y2=1.22
r229 34 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.69 $Y=0.865
+ $X2=0.69 $Y2=1.22
r230 12 87 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=4.565
r231 12 85 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=3.205
r232 11 73 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.565
r233 11 71 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.205
r234 10 59 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.565
r235 10 57 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.205
r236 9 45 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r237 9 43 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r238 4 76 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.865
r239 3 62 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.865
r240 2 48 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.865
r241 1 34 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

