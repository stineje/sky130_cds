* File: sky130_osu_sc_12T_ls__inv_4.pex.spice
* Created: Fri Nov 12 15:37:56 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__INV_4%GND 1 2 3 31 35 37 44 46 54 64 66
r57 64 66 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r58 52 54 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r59 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r60 46 52 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.305
r61 42 60 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r62 42 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r63 37 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r64 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r65 31 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r66 31 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r67 31 33 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r68 31 38 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r69 31 46 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r70 31 47 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r71 31 37 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r72 31 38 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r73 3 54 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84 $Y=0.575
+ $X2=1.98 $Y2=0.755
r74 2 44 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
r75 1 35 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_4%VDD 1 2 3 25 29 31 37 41 48 57 61
r39 57 61 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.7 $Y2=4.287
r40 53 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r41 48 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r42 46 51 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135 $X2=1.98
+ $Y2=3.635
r43 44 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=4.25 $X2=1.7
+ $Y2=4.25
r44 42 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r45 42 44 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r46 41 46 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.135
r47 41 44 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r48 37 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r49 35 55 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r50 35 40 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135 $X2=1.12
+ $Y2=3.635
r51 32 53 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r52 32 34 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r53 31 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r54 31 34 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r55 27 53 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r56 27 29 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135 $X2=0.26
+ $Y2=3.635
r57 25 44 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r58 25 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r59 25 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r60 3 51 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r61 3 48 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r62 2 40 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r63 2 37 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r64 1 29 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_4%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 44 46 47 48 49 50 53 55 57 60
c120 43 0 1.50926e-19 $X=0.535 $Y=1.825
c121 28 0 1.33323e-19 $X=1.335 $Y=2.48
c122 25 0 1.33323e-19 $X=1.335 $Y=1.22
c123 18 0 1.33323e-19 $X=0.905 $Y=2.48
c124 15 0 1.33323e-19 $X=0.905 $Y=1.22
r125 60 63 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=2.845
+ $X2=0.405 $Y2=2.85
r126 55 57 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=1.825
+ $X2=0.535 $Y2=1.825
r127 53 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r128 51 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.405 $Y2=1.825
r129 51 53 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.32 $Y2=2.85
r130 43 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.825 $X2=0.535 $Y2=1.825
r131 43 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.99
r132 43 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.66
r133 38 40 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r134 35 37 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.765 $Y=1.22
+ $X2=1.765 $Y2=0.835
r135 34 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.405
+ $X2=1.335 $Y2=2.405
r136 33 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.48
r137 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.41 $Y2=2.405
r138 32 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.335 $Y2=1.295
r139 31 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=1.295
+ $X2=1.765 $Y2=1.22
r140 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.295
+ $X2=1.41 $Y2=1.295
r141 28 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=2.405
r142 28 30 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r143 25 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=1.295
r144 25 27 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=0.835
r145 24 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.405
+ $X2=0.905 $Y2=2.405
r146 23 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=1.335 $Y2=2.405
r147 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=0.98 $Y2=2.405
r148 22 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.295
+ $X2=0.905 $Y2=1.295
r149 21 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=1.335 $Y2=1.295
r150 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=0.98 $Y2=1.295
r151 18 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=2.405
r152 18 20 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=3.235
r153 15 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=1.295
r154 15 17 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=0.835
r155 14 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.405
+ $X2=0.475 $Y2=2.405
r156 13 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.905 $Y2=2.405
r157 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.55 $Y2=2.405
r158 12 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.475 $Y2=1.295
r159 11 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.905 $Y2=1.295
r160 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.55 $Y2=1.295
r161 8 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=2.405
r162 8 10 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=3.235
r163 7 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=2.405
r164 7 45 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=1.99
r165 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.295
r166 4 44 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.66
r167 1 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=1.295
r168 1 3 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_4%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c88 55 0 1.33323e-19 $X=1.55 $Y=2.365
c89 54 0 1.33323e-19 $X=1.55 $Y=1.115
c90 46 0 1.33323e-19 $X=0.69 $Y=2.365
c91 45 0 1.33323e-19 $X=0.69 $Y=1.115
c92 18 0 1.50926e-19 $X=0.69 $Y=0.755
r93 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.48
r94 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r95 54 55 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=2.365
r96 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.48
+ $X2=0.69 $Y2=2.48
r97 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=1.55 $Y2=2.48
r98 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=0.835 $Y2=2.48
r99 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1
+ $X2=0.69 $Y2=1
r100 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=1.55 $Y2=1
r101 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=0.835 $Y2=1
r102 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.48
r103 46 48 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=1.72
r104 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1
r105 45 48 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1.72
r106 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r107 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.48
r108 38 41 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.955
r109 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r110 32 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r111 27 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r112 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r113 24 27 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.955
r114 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1 $X2=0.69
+ $Y2=1
r115 18 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0.755
+ $X2=0.69 $Y2=1
r116 6 43 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r117 6 41 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r118 5 29 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r119 5 27 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r120 2 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
r121 1 18 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

