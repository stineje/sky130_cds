* File: sky130_osu_sc_12T_ms__or2_1.pex.spice
* Created: Fri Nov 12 15:26:02 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__OR2_1%GND 1 2 21 25 27 35 42 44 47
r38 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r39 33 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r40 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r41 27 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r42 23 25 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r43 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r44 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r45 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r46 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r47 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r48 2 35 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
r49 1 25 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_1%VDD 1 13 15 24 28 30 33
r23 30 33 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r24 22 28 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r25 22 24 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135 $X2=1.12
+ $Y2=3.635
r26 20 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r27 17 20 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r28 15 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r29 15 20 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r30 13 20 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r31 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r32 1 24 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_1%B 3 7 12 15 21
r28 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.48
r29 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.195
+ $X2=0.27 $Y2=2.48
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.195 $X2=0.27 $Y2=2.195
r31 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.195
+ $X2=0.475 $Y2=2.195
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=2.195
r33 5 7 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=3.235
r34 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.03
+ $X2=0.475 $Y2=2.195
r35 1 3 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.475 $Y=2.03
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_1%A 3 7 10 14 20
r44 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.85
+ $X2=0.95 $Y2=2.85
r45 14 17 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=2.85
r46 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.905 $X2=0.95 $Y2=1.905
r47 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=2.07
r48 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=1.74
r49 7 12 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.07
r50 3 11 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=0.905 $Y=0.835
+ $X2=0.905 $Y2=1.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_1%A_27_521# 1 3 11 15 16 18 19 24 26 27 29
+ 32 36 38
r70 34 38 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.455
+ $X2=0.65 $Y2=1.455
r71 34 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.455
+ $X2=1.43 $Y2=1.455
r72 30 38 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.65 $Y2=1.455
r73 30 32 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.69 $Y2=0.755
r74 28 38 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.65 $Y2=1.455
r75 28 29 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=3.065
r76 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.15
+ $X2=0.61 $Y2=3.065
r77 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.15
+ $X2=0.345 $Y2=3.15
r78 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.235
+ $X2=0.345 $Y2=3.15
r79 22 24 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.26 $Y=3.235 $X2=0.26
+ $Y2=3.295
r80 21 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.455 $X2=1.43 $Y2=1.455
r81 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.33
+ $X2=1.352 $Y2=2.48
r82 16 21 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.412 $Y2=1.455
r83 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=2.33
r84 15 19 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=3.235
+ $X2=1.335 $Y2=2.48
r85 9 21 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.412 $Y2=1.455
r86 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.835
r87 3 24 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.295
r88 1 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_1%Y 1 3 10 16 26 29 32
r36 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=2.11
r37 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=1.74
r38 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r39 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.74
r40 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r41 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.11
r42 16 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.955
r43 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r44 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r45 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r46 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r47 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41 $Y=0.575
+ $X2=1.55 $Y2=0.755
.ends

