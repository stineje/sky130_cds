* File: sky130_osu_sc_18T_ls__oai21_l.spice
* Created: Fri Nov 12 14:18:52 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_ls__oai21_l.pex.spice"
.subckt sky130_osu_sc_18T_ls__oai21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1005 N_GND_M1005_d N_A0_M1005_g N_A_27_115#_M1005_s N_GND_M1005_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1001 N_A_27_115#_M1001_d N_A1_M1001_g N_GND_M1005_d N_GND_M1005_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_115#_M1001_d N_GND_M1005_b NSHORT L=0.15
+ W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 A_110_617# N_A0_M1004_g N_Y_M1004_s N_VDD_M1004_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.9 A=0.45 P=6.3 MULT=1
MM1003 N_VDD_M1003_d N_A1_M1003_g A_110_617# N_VDD_M1004_b PHIGHVT L=0.15 W=3
+ AD=0.567 AS=0.315 PD=4.008 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75000.5
+ SB=75000.5 A=0.45 P=6.3 MULT=1
MM1000 N_Y_M1000_d N_B0_M1000_g N_VDD_M1003_d N_VDD_M1004_b PHIGHVT L=0.15 W=2
+ AD=0.53 AS=0.378 PD=4.53 PS=2.672 NRD=0 NRS=5.8903 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1005_b N_VDD_M1004_b NWDIODE A=7.277 P=11.43
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__oai21_l.pxi.spice"
*
.ends
*
*
