* File: sky130_osu_sc_18T_hs__addh_l.spice
* Created: Thu Oct 29 17:05:39 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_hs__addh_l.pex.spice"
.subckt sky130_osu_sc_18T_hs__addh_l  GND VDD CON B A S CO
* 
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1005 N_GND_M1005_d N_CON_M1005_g N_S_M1005_s N_GND_M1005_b NLOWVT L=0.15
+ W=0.64 AD=0.122146 AS=0.1696 PD=1.04585 PS=1.81 NRD=11.712 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1008 A_208_115# N_B_M1008_g N_GND_M1005_d N_GND_M1005_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.190854 PD=1.21 PS=1.63415 NRD=5.988 NRS=0 M=1 R=6.66667
+ SA=75000.5 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1009 N_A_208_617#_M1009_d N_A_M1009_g A_208_115# N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_GND_M1002_d N_A_208_617#_M1002_g N_CO_M1002_s N_GND_M1005_b NLOWVT
+ L=0.15 W=0.64 AD=0.122146 AS=0.1696 PD=1.04585 PS=1.81 NRD=11.712 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1010 N_A_570_115#_M1010_d N_A_208_617#_M1010_g N_GND_M1002_d N_GND_M1005_b
+ NLOWVT L=0.15 W=1 AD=0.14 AS=0.190854 PD=1.28 PS=1.63415 NRD=0 NRS=0 M=1
+ R=6.66667 SA=75000.5 SB=75001 A=0.15 P=2.3 MULT=1
MM1003 N_CON_M1003_d N_B_M1003_g N_A_570_115#_M1010_d N_GND_M1005_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.9 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1004 N_A_570_115#_M1004_d N_A_M1004_g N_CON_M1003_d N_GND_M1005_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_VDD_M1001_d N_CON_M1001_g N_S_M1001_s N_VDD_M1001_b PSHORT L=0.15
+ W=1.65 AD=0.326008 AS=0.43725 PD=2.37032 PS=3.83 NRD=7.2693 NRS=0 M=1 R=11
+ SA=75000.2 SB=75001.6 A=0.2475 P=3.6 MULT=1
MM1006 N_A_208_617#_M1006_d N_B_M1006_g N_VDD_M1001_d N_VDD_M1001_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.592742 PD=3.28 PS=4.30968 NRD=0 NRS=0 M=1 R=20
+ SA=75000.5 SB=75000.9 A=0.45 P=6.3 MULT=1
MM1007 N_VDD_M1007_d N_A_M1007_g N_A_208_617#_M1006_d N_VDD_M1001_b PSHORT
+ L=0.15 W=3 AD=0.592742 AS=0.42 PD=4.30968 PS=3.28 NRD=0 NRS=0 M=1 R=20
+ SA=75000.9 SB=75000.5 A=0.45 P=6.3 MULT=1
MM1011 N_CO_M1011_d N_A_208_617#_M1011_g N_VDD_M1007_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.65 AD=0.43725 AS=0.326008 PD=3.83 PS=2.37032 NRD=0 NRS=7.2693 M=1
+ R=11 SA=75001.6 SB=75000.2 A=0.2475 P=3.6 MULT=1
MM1000 N_VDD_M1000_d N_A_208_617#_M1000_g N_CON_M1000_s N_VDD_M1001_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1012 A_668_617# N_B_M1012_g N_VDD_M1000_d N_VDD_M1001_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1013 N_CON_M1013_d N_A_M1013_g A_668_617# N_VDD_M1001_b PSHORT L=0.15 W=3
+ AD=0.84 AS=0.315 PD=6.56 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX14_noxref N_GND_M1005_b N_VDD_M1001_b NWDIODE A=16.074 P=16.06
pX15_noxref noxref_12 S S PROBETYPE=1
pX16_noxref noxref_13 CO CO PROBETYPE=1
pX17_noxref noxref_14 B B PROBETYPE=1
pX18_noxref noxref_15 CON CON PROBETYPE=1
pX19_noxref noxref_16 A A PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__addh_l.pxi.spice"
*
.ends
*
*
