* File: sky130_osu_sc_15T_hs__buf_2.spice
* Created: Fri Nov 12 14:28:09 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__buf_2.pex.spice"
.subckt sky130_osu_sc_15T_hs__buf_2  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1004_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_Y_M1000_d N_A_27_115#_M1001_g N_GND_M1001_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VDD_M1005_d N_A_M1005_g N_A_27_115#_M1005_s N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1002 N_Y_M1002_d N_A_27_115#_M1002_g N_VDD_M1005_d N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1003 N_Y_M1002_d N_A_27_115#_M1003_g N_VDD_M1003_s N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1005_b NWDIODE A=5.67875 P=9.75
pX7_noxref noxref_6 A A PROBETYPE=1
pX8_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__buf_2.pxi.spice"
*
.ends
*
*
