* File: sky130_osu_sc_18T_ls__and2_2.spice
* Created: Thu Oct 29 17:33:42 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ls__and2_2.pex.spice"
.subckt sky130_osu_sc_18T_ls__and2_2  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 A_110_115# N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1004_b NSHORT L=0.15 W=1
+ AD=0.175 AS=0.105 PD=1.35 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75000.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1001_d N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.175 PD=1.28 PS=1.35 NRD=0 NRS=8.388 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1000_d N_A_27_115#_M1006_g N_GND_M1006_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_27_115#_M1003_d N_A_M1003_g N_VDD_M1003_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001.5 A=0.45 P=6.3 MULT=1
MM1007 N_VDD_M1007_d N_B_M1007_g N_A_27_115#_M1003_d N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1002 N_VDD_M1007_d N_A_27_115#_M1002_g N_Y_M1002_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1005 N_VDD_M1005_d N_A_27_115#_M1005_g N_Y_M1002_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.5
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX8_noxref N_GND_M1004_b N_VDD_M1003_b NWDIODE A=8.949 P=12.31
pX9_noxref noxref_8 A A PROBETYPE=1
pX10_noxref noxref_9 B B PROBETYPE=1
pX11_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__and2_2.pxi.spice"
*
.ends
*
*
