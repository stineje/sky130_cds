* File: sky130_osu_sc_12T_hs__dffsr_1.spice
* Created: Fri Nov 12 15:09:47 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__dffsr_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffsr_1  GND VDD RN SN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* RN	RN
* VDD	VDD
* GND	GND
MM1016 N_A_110_115#_M1016_d N_RN_M1016_g N_GND_M1016_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1034 N_A_217_521#_M1034_d N_A_110_115#_M1034_g N_GND_M1034_s N_GND_M1016_b
+ NLOWVT L=0.15 W=0.42 AD=0.0767474 AS=0.1113 PD=0.770722 PS=1.37 NRD=17.136
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1015 A_400_115# N_SN_M1015_g N_A_217_521#_M1034_d N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.100503 PD=0.76 PS=1.00928 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1003 N_GND_M1003_d N_A_432_424#_M1003_g A_400_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.9 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 A_662_115# N_D_M1005_g N_GND_M1005_s N_GND_M1016_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1035 N_A_432_424#_M1035_d N_A_704_89#_M1035_g A_662_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1026 A_854_115# N_CK_M1026_g N_A_432_424#_M1035_d N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1020 N_GND_M1020_d N_A_217_521#_M1020_g A_854_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1023 A_1012_115# N_A_217_521#_M1023_g N_GND_M1020_d N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1021 N_A_1084_115#_M1021_d N_CK_M1021_g A_1012_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1017 A_1204_115# N_A_704_89#_M1017_g N_A_1084_115#_M1021_d N_GND_M1016_b
+ NLOWVT L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54
+ M=1 R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1006 N_GND_M1006_d N_A_1246_89#_M1006_g A_1204_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_A_704_89#_M1011_d N_CK_M1011_g N_GND_M1006_d N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1013 A_1552_115# N_A_1084_115#_M1013_g N_GND_M1013_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1004 N_A_1246_89#_M1004_d N_SN_M1004_g A_1552_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.100503 AS=0.05775 PD=1.00928 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1022 N_GND_M1022_d N_A_110_115#_M1022_g N_A_1246_89#_M1004_d N_GND_M1016_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0767474 PD=1.37 PS=0.770722 NRD=0
+ NRS=17.136 M=1 R=2.8 SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_GND_M1007_d N_A_1246_89#_M1007_g N_QN_M1007_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1008 N_Q_M1008_d N_QN_M1008_g N_GND_M1007_d N_GND_M1016_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1001 N_A_110_115#_M1001_d N_RN_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_300_521#_M1000_d N_A_110_115#_M1000_g N_A_217_521#_M1000_s
+ N_VDD_M1001_b PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0
+ NRS=0 M=1 R=8.4 SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1024 N_VDD_M1024_d N_SN_M1024_g N_A_300_521#_M1000_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_A_300_521#_M1027_d N_A_432_424#_M1027_g N_VDD_M1024_d N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1028 A_662_521# N_D_M1028_g N_VDD_M1028_s N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1018 N_A_432_424#_M1018_d N_CK_M1018_g A_662_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1014 A_854_521# N_A_704_89#_M1014_g N_A_432_424#_M1018_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1009 N_VDD_M1009_d N_A_217_521#_M1009_g A_854_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1012 A_1012_521# N_A_217_521#_M1012_g N_VDD_M1009_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1010 N_A_1084_115#_M1010_d N_A_704_89#_M1010_g A_1012_521# N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778
+ NRS=7.8012 M=1 R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 A_1204_521# N_CK_M1002_g N_A_1084_115#_M1010_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1029 N_VDD_M1029_d N_A_1246_89#_M1029_g A_1204_521# N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1031 N_A_704_89#_M1031_d N_CK_M1031_g N_VDD_M1029_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1033 N_VDD_M1033_d N_A_1084_115#_M1033_g N_A_1469_521#_M1033_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1019 N_A_1469_521#_M1019_d N_SN_M1019_g N_VDD_M1033_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_A_1246_89#_M1025_d N_A_110_115#_M1025_g N_A_1469_521#_M1019_d
+ N_VDD_M1001_b PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0
+ NRS=0 M=1 R=8.4 SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1030 N_VDD_M1030_d N_A_1246_89#_M1030_g N_QN_M1030_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1032 N_Q_M1032_d N_QN_M1032_g N_VDD_M1030_d N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref N_GND_M1016_b N_VDD_M1001_b NWDIODE A=21.63 P=25.12
pX37_noxref noxref_27 RN RN PROBETYPE=1
pX38_noxref noxref_28 D D PROBETYPE=1
pX39_noxref noxref_29 CK CK PROBETYPE=1
pX40_noxref noxref_30 SN SN PROBETYPE=1
pX41_noxref noxref_31 QN QN PROBETYPE=1
pX42_noxref noxref_32 Q Q PROBETYPE=1
c_2169 A_1012_521# 0 1.57671e-19 $X=5.06 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffsr_1.pxi.spice"
*
.ends
*
*
