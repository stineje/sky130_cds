* File: sky130_osu_sc_18T_ms__nand2_l.pex.spice
* Created: Thu Oct 29 17:30:36 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_L%GND 1 12 14 21 24 27
r24 24 27 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r25 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r26 12 19 4.26217 $w=1.7e-07 $l=2.14243e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=1.05 $Y2=0.305
r27 12 14 3.29607 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=0.965 $Y2=0.152
r28 12 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r29 12 14 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r30 1 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_L%VDD 1 2 13 17 23 30 32 35
r15 35 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r16 32 35 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r17 30 39 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r18 27 39 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r19 27 29 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r20 23 26 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=4.815
+ $X2=1.12 $Y2=5.835
r21 21 30 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.035 $Y2=6.507
r22 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r23 17 20 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=4.815
+ $X2=0.26 $Y2=5.835
r24 15 29 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r25 15 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r26 13 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r27 13 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r28 2 26 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=5.835
r29 2 23 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=4.815
r30 1 20 300 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=5.835
r31 1 17 300 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=4.815
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_L%A 3 7 10 15 16
r27 16 18 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.685
+ $X2=0.367 $Y2=2.85
r28 16 17 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.685
+ $X2=0.367 $Y2=2.52
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.685 $X2=0.32 $Y2=2.685
r30 12 15 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=2.685
r31 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r32 7 18 1146.03 $w=1.5e-07 $l=2.235e-06 $layer=POLY_cond $X=0.475 $Y=5.085
+ $X2=0.475 $Y2=2.85
r33 3 17 807.606 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=2.52
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_L%B 3 7 11 13 17 19
c35 11 0 1.91696e-19 $X=0.915 $Y=1.935
c36 3 0 1.57512e-19 $X=0.835 $Y=0.945
r37 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.06 $Y=2.96
+ $X2=1.06 $Y2=2.96
r38 14 19 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.06 $Y=2.02
+ $X2=1.06 $Y2=2.96
r39 13 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.935
+ $X2=1.06 $Y2=2.02
r40 11 22 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.935
+ $X2=0.905 $Y2=1.77
r41 10 13 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.915 $Y=1.935
+ $X2=1.06 $Y2=1.935
r42 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=1.935 $X2=0.915 $Y2=1.935
r43 5 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.1
+ $X2=0.905 $Y2=1.935
r44 5 7 1530.61 $w=1.5e-07 $l=2.985e-06 $layer=POLY_cond $X=0.905 $Y=2.1
+ $X2=0.905 $Y2=5.085
r45 3 22 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=1.77
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_L%Y 1 2 7 8 12 19 20 23
c37 20 0 1.91696e-19 $X=0.69 $Y=2.59
c38 8 0 1.57512e-19 $X=0.405 $Y=1.48
r39 30 32 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=4.815
+ $X2=0.69 $Y2=5.835
r40 20 30 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=0.69 $Y=2.59
+ $X2=0.69 $Y2=4.815
r41 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.59
+ $X2=0.69 $Y2=2.59
r42 16 23 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.26 $Y=1.48
+ $X2=0.26 $Y2=0.825
r43 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.48
+ $X2=0.26 $Y2=1.48
r44 10 19 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.475
+ $X2=0.69 $Y2=2.59
r45 10 12 0.12036 $w=1.7e-07 $l=1.25e-07 $layer=MET1_cond $X=0.69 $Y=2.475
+ $X2=0.69 $Y2=2.35
r46 9 12 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=0.69 $Y=1.565
+ $X2=0.69 $Y2=2.35
r47 8 15 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=1.48
+ $X2=0.26 $Y2=1.48
r48 7 9 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=1.48
+ $X2=0.69 $Y2=1.565
r49 7 8 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=1.48 $X2=0.405
+ $Y2=1.48
r50 2 32 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=5.835
r51 2 30 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=4.815
r52 1 23 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

