* File: sky130_osu_sc_15T_hs__aoi21_l.spice
* Created: Fri Nov 12 14:27:44 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__aoi21_l.pex.spice"
.subckt sky130_osu_sc_15T_hs__aoi21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A0_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_110_115# N_GND_M1003_b NLOWVT L=0.15 W=0.64
+ AD=0.113398 AS=0.0672 PD=1.05412 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1004 N_GND_M1004_d N_B0_M1004_g N_Y_M1000_d N_GND_M1003_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.0974517 PD=1.63 PS=0.905882 NRD=0 NRS=13.08 M=1 R=3.66667
+ SA=75001 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 N_VDD_M1005_d N_A0_M1005_g N_A_27_565#_M1005_s N_VDD_M1005_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1001 N_A_27_565#_M1001_d N_A1_M1001_g N_VDD_M1005_d N_VDD_M1005_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_565#_M1001_d N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1005_b NWDIODE A=5.64925 P=9.73
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__aoi21_l.pxi.spice"
*
.ends
*
*
