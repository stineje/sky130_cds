* File: sky130_osu_sc_15T_ms__nor2_l.spice
* Created: Fri Nov 12 14:45:27 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__nor2_l.pex.spice"
.subckt sky130_osu_sc_15T_ms__nor2_l  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_Y_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NSHORT L=0.15 W=0.52
+ AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1003_d N_GND_M1003_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1002 A_110_713# N_B_M1002_g N_Y_M1002_s N_VDD_M1002_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g A_110_713# N_VDD_M1002_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=4.35125 P=8.85
pX5_noxref noxref_7 B B PROBETYPE=1
pX6_noxref noxref_8 Y Y PROBETYPE=1
pX7_noxref noxref_9 A A PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__nor2_l.pxi.spice"
*
.ends
*
*
