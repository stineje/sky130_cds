* File: sky130_osu_sc_12T_hs__inv_8.spice
* Created: Fri Nov 12 15:11:19 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__inv_8.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_8  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1006 N_GND_M1002_d N_A_M1006_g N_Y_M1006_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1011 N_GND_M1011_d N_A_M1011_g N_Y_M1006_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1012 N_GND_M1011_d N_A_M1012_g N_Y_M1012_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1013 N_GND_M1013_d N_A_M1013_g N_Y_M1012_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1014 N_GND_M1013_d N_A_M1014_g N_Y_M1014_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1015 N_GND_M1015_d N_A_M1015_g N_Y_M1014_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_VDD_M1008_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VDD_M1008_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1009_d N_A_M1010_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=8.4769 P=12.35
pX17_noxref noxref_5 A A PROBETYPE=1
pX18_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_8.pxi.spice"
*
.ends
*
*
