* File: sky130_osu_sc_12T_hs__xnor2_l.pex.spice
* Created: Fri Nov 12 15:14:07 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%GND 1 2 33 35 43 45 55 67 69
r74 67 69 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r75 53 55 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.74
r76 46 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r77 41 59 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r78 41 43 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r79 35 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r80 33 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r81 33 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r82 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r83 33 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r84 33 45 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r85 33 46 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r86 33 35 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r87 2 55 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.575 $X2=2.44 $Y2=0.74
r88 1 43 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%VDD 1 2 25 27 34 38 46 54 57 61
c40 34 0 1.59951e-19 $X=0.69 $Y=2.955
r41 57 61 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=2.38 $Y2=4.287
r42 54 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=4.25
+ $X2=2.38 $Y2=4.25
r43 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.44 $Y=2.955
+ $X2=2.44 $Y2=3.635
r44 44 54 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=4.135
+ $X2=2.44 $Y2=4.287
r45 44 49 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.44 $Y=4.135 $X2=2.44
+ $Y2=3.635
r46 41 43 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r47 39 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r48 39 41 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r49 38 54 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=4.287
+ $X2=2.44 $Y2=4.287
r50 38 43 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=4.287
+ $X2=1.7 $Y2=4.287
r51 34 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r52 32 52 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r53 32 37 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135 $X2=0.69
+ $Y2=3.635
r54 29 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r55 27 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r56 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r57 25 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r58 25 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r59 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r60 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r61 2 49 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.605 $X2=2.44 $Y2=3.635
r62 2 46 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.605 $X2=2.44 $Y2=2.955
r63 1 37 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r64 1 34 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A 3 5 8 9 13 16 18 19 20 21 22 26 30 36
+ 40 41 42 46 51 52
c121 36 0 1.96463e-19 $X=2.105 $Y=1.74
r122 51 52 0.0806629 $w=2.95e-07 $l=1.15e-07 $layer=MET1_cond $X=2.107 $Y=1.74
+ $X2=2.107 $Y2=1.625
r123 43 52 0.519956 $w=1.7e-07 $l=5.4e-07 $layer=MET1_cond $X=2.105 $Y=1.085
+ $X2=2.105 $Y2=1.625
r124 41 43 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=2.02 $Y=1
+ $X2=2.105 $Y2=1.085
r125 41 42 1.04954 $w=1.7e-07 $l=1.09e-06 $layer=MET1_cond $X=2.02 $Y=1 $X2=0.93
+ $Y2=1
r126 40 46 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.845 $Y=1.255
+ $X2=0.845 $Y2=1.37
r127 39 42 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.845
+ $Y=1.085 $X2=0.93 $Y2=1
r128 39 40 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=0.845 $Y=1.085
+ $X2=0.845 $Y2=1.255
r129 36 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.105 $Y=1.74
+ $X2=2.105 $Y2=1.74
r130 36 38 9.34866 $w=2.61e-07 $l=2e-07 $layer=LI1_cond $X=2.19 $Y=1.74 $X2=2.19
+ $Y2=1.94
r131 30 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.845 $Y=1.37
+ $X2=0.845 $Y2=1.37
r132 30 33 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.845 $Y=1.37
+ $X2=0.845 $Y2=1.4
r133 28 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=1.94 $X2=2.225 $Y2=1.94
r134 26 28 73.8383 $w=2.35e-07 $l=3.6e-07 $layer=POLY_cond $X=1.865 $Y=1.955
+ $X2=2.225 $Y2=1.955
r135 24 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.4 $X2=0.845 $Y2=1.4
r136 21 24 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=0.845 $Y=1.275
+ $X2=0.845 $Y2=1.4
r137 21 22 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.275
+ $X2=0.845 $Y2=1.2
r138 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.45 $Y=2.38 $X2=0.45
+ $Y2=2.53
r139 14 26 13.2911 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.865 $Y=2.105
+ $X2=1.865 $Y2=1.955
r140 14 16 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=1.865 $Y=2.105
+ $X2=1.865 $Y2=3.235
r141 13 22 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.905 $Y=0.85
+ $X2=0.905 $Y2=1.2
r142 10 18 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=1.275
+ $X2=0.45 $Y2=1.275
r143 9 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=1.275
+ $X2=0.845 $Y2=1.275
r144 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=1.275
+ $X2=0.55 $Y2=1.275
r145 8 20 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=2.53
r146 3 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=1.2
+ $X2=0.45 $Y2=1.275
r147 3 5 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.475 $Y=1.2
+ $X2=0.475 $Y2=0.85
r148 1 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=1.35
+ $X2=0.45 $Y2=1.275
r149 1 19 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=0.425 $Y=1.35
+ $X2=0.425 $Y2=2.38
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A_27_115# 1 3 11 13 15 17 21 25 29 33
+ 39 41
r84 37 39 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.765 $Y=1.855
+ $X2=1.765 $Y2=1.4
r85 34 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.94
+ $X2=0.26 $Y2=1.94
r86 34 36 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=1.94
+ $X2=0.845 $Y2=1.94
r87 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=1.94
+ $X2=1.765 $Y2=1.855
r88 33 36 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.68 $Y=1.94
+ $X2=0.845 $Y2=1.94
r89 29 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r90 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.025
+ $X2=0.26 $Y2=1.94
r91 27 29 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.26 $Y=2.025
+ $X2=0.26 $Y2=2.955
r92 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.855
+ $X2=0.26 $Y2=1.94
r93 23 25 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=0.26 $Y=1.855
+ $X2=0.26 $Y2=0.755
r94 21 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.4 $X2=1.765 $Y2=1.4
r95 21 22 15.9603 $w=3.02e-07 $l=1e-07 $layer=POLY_cond $X=1.765 $Y=1.4
+ $X2=1.865 $Y2=1.4
r96 17 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.94 $X2=0.845 $Y2=1.94
r97 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=1.94
+ $X2=0.845 $Y2=2.105
r98 13 22 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.235
+ $X2=1.865 $Y2=1.4
r99 13 15 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.865 $Y=1.235
+ $X2=1.865 $Y2=0.85
r100 11 19 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.105
r101 3 31 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r102 3 29 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r103 1 25 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A_238_89# 1 3 11 15 18 21 27 31 35
r64 31 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.87 $Y=2.955
+ $X2=2.87 $Y2=3.635
r65 29 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.37 $X2=2.87
+ $Y2=2.285
r66 29 31 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.87 $Y=2.37
+ $X2=2.87 $Y2=2.955
r67 25 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.2 $X2=2.87
+ $Y2=2.285
r68 25 27 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=2.87 $Y=2.2
+ $X2=2.87 $Y2=0.755
r69 21 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=2.285
+ $X2=2.87 $Y2=2.285
r70 21 23 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=2.285
+ $X2=1.325 $Y2=2.285
r71 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.285 $X2=1.325 $Y2=2.285
r72 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.285
+ $X2=1.325 $Y2=2.45
r73 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.285
+ $X2=1.325 $Y2=2.12
r74 15 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.265 $Y=3.235
+ $X2=1.265 $Y2=2.45
r75 11 19 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.265 $Y=0.85
+ $X2=1.265 $Y2=2.12
r76 3 33 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.605 $X2=2.87 $Y2=3.635
r77 3 31 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.605 $X2=2.87 $Y2=2.955
r78 1 27 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.73 $Y=0.575
+ $X2=2.87 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 20 21 23 31
c57 31 0 1.96463e-19 $X=2.53 $Y=1.4
r58 29 31 0.0101078 $w=3.71e-07 $l=3e-08 $layer=MET1_cond $X=2.585 $Y=1.37
+ $X2=2.585 $Y2=1.4
r59 23 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.37
+ $X2=2.53 $Y2=1.37
r60 23 26 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.53 $Y=1.37 $X2=2.53
+ $Y2=1.4
r61 19 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.4 $X2=2.53 $Y2=1.4
r62 19 20 21.9891 $w=2.74e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=1.382
+ $X2=2.655 $Y2=1.382
r63 14 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=2.53
+ $X2=2.655 $Y2=2.455
r64 14 16 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.655 $Y=2.53
+ $X2=2.655 $Y2=3.235
r65 13 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=2.38
+ $X2=2.655 $Y2=2.455
r66 12 20 16.847 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=2.655 $Y=1.565
+ $X2=2.655 $Y2=1.382
r67 12 13 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.655 $Y=1.565
+ $X2=2.655 $Y2=2.38
r68 9 20 16.847 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.655 $Y=1.2
+ $X2=2.655 $Y2=1.382
r69 9 11 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.655 $Y=1.2
+ $X2=2.655 $Y2=0.85
r70 7 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=2.455
+ $X2=2.655 $Y2=2.455
r71 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=2.455 $X2=2.3
+ $Y2=2.455
r72 4 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=2.53
+ $X2=2.3 $Y2=2.455
r73 4 6 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.225 $Y=2.53
+ $X2=2.225 $Y2=3.235
r74 1 19 53.6533 $w=2.74e-07 $l=3.85402e-07 $layer=POLY_cond $X=2.225 $Y=1.2
+ $X2=2.53 $Y2=1.382
r75 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.225 $Y=1.2 $X2=2.225
+ $Y2=0.85
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XNOR2_L%Y 1 3 11 13 15 17 27 30 33
c59 27 0 1.59951e-19 $X=1.42 $Y=1.655
r60 25 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=2.735
+ $X2=1.425 $Y2=2.85
r61 25 27 1.03991 $w=1.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.425 $Y=2.735
+ $X2=1.425 $Y2=1.655
r62 24 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.485
+ $X2=1.425 $Y2=1.37
r63 24 27 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.425 $Y=1.485
+ $X2=1.425 $Y2=1.655
r64 21 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=2.85
+ $X2=1.425 $Y2=2.85
r65 21 23 3.32727 $w=3.85e-07 $l=1.05e-07 $layer=LI1_cond $X=1.537 $Y=2.85
+ $X2=1.537 $Y2=2.955
r66 17 19 5.12913 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.425 $Y=0.755
+ $X2=1.565 $Y2=0.755
r67 13 23 0.513842 $w=3.85e-07 $l=3.2619e-08 $layer=LI1_cond $X=1.565 $Y=2.965
+ $X2=1.537 $Y2=2.955
r68 13 15 22.7099 $w=3.38e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=2.965
+ $X2=1.565 $Y2=3.635
r69 11 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=1.37
+ $X2=1.425 $Y2=1.37
r70 9 17 4.67747 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.425 $Y=0.935
+ $X2=1.425 $Y2=0.755
r71 9 11 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.425 $Y=0.935
+ $X2=1.425 $Y2=1.37
r72 3 15 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.565 $Y2=3.635
r73 3 23 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.565 $Y2=2.955
r74 1 19 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.755
.ends

