* File: sky130_osu_sc_15T_ls__dff_l.pex.spice
* Created: Fri Nov 12 14:55:42 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%GND 1 2 3 4 5 81 83 91 93 103 105 115 117
+ 124 126 133 152 154
c172 81 0 1.27355e-19 $X=-0.045 $Y=0
r173 152 154 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r174 131 133 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.545 $Y=0.305
+ $X2=6.545 $Y2=0.74
r175 122 124 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.165 $Y=0.305
+ $X2=5.165 $Y2=0.865
r176 118 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.152
+ $X2=4.215 $Y2=0.152
r177 113 141 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.152
r178 113 115 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.865
r179 105 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.152
+ $X2=4.215 $Y2=0.152
r180 101 103 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.465 $Y=0.305
+ $X2=2.465 $Y2=0.74
r181 94 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.152
+ $X2=0.715 $Y2=0.152
r182 89 137 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.152
r183 89 91 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.865
r184 83 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.152
+ $X2=0.715 $Y2=0.152
r185 81 154 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r186 81 152 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r187 81 131 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.545 $Y2=0.305
r188 81 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.46 $Y2=0.152
r189 81 122 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.165 $Y2=0.305
r190 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.08 $Y2=0.152
r191 81 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.25 $Y2=0.152
r192 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.465 $Y2=0.305
r193 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.38 $Y2=0.152
r194 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.55 $Y2=0.152
r195 81 126 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.46 $Y2=0.152
r196 81 127 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.25 $Y2=0.152
r197 81 117 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=5.08 $Y2=0.152
r198 81 118 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.3 $Y2=0.152
r199 81 105 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.13 $Y2=0.152
r200 81 106 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.55 $Y2=0.152
r201 81 93 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.38 $Y2=0.152
r202 81 94 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.8 $Y2=0.152
r203 81 83 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.63 $Y2=0.152
r204 5 133 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.405
+ $Y=0.575 $X2=6.545 $Y2=0.74
r205 4 124 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.575 $X2=5.165 $Y2=0.865
r206 3 115 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.575 $X2=4.215 $Y2=0.865
r207 2 103 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.74
r208 1 91 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.575 $X2=0.715 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%VDD 1 2 3 4 5 61 63 70 74 82 86 94 98 104
+ 108 114 125 128 132
c98 70 0 5.41559e-20 $X=0.715 $Y=3.545
c99 1 0 1.59851e-19 $X=0.575 $Y=2.825
r100 128 132 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=6.46 $Y2=5.397
r101 125 132 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=5.36
+ $X2=6.46 $Y2=5.36
r102 112 125 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=5.245
+ $X2=6.545 $Y2=5.397
r103 112 114 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.545 $Y=5.245
+ $X2=6.545 $Y2=4.565
r104 109 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.25 $Y=5.397
+ $X2=5.165 $Y2=5.397
r105 109 111 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.25 $Y=5.397
+ $X2=5.78 $Y2=5.397
r106 108 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=5.397
+ $X2=6.545 $Y2=5.397
r107 108 111 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.46 $Y=5.397
+ $X2=5.78 $Y2=5.397
r108 104 107 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=5.165 $Y=3.545
+ $X2=5.165 $Y2=4.565
r109 102 123 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.165 $Y=5.245
+ $X2=5.165 $Y2=5.397
r110 102 107 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.165 $Y=5.245
+ $X2=5.165 $Y2=4.565
r111 99 121 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=5.397
+ $X2=4.215 $Y2=5.397
r112 99 101 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.3 $Y=5.397
+ $X2=4.42 $Y2=5.397
r113 98 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=5.397
+ $X2=5.165 $Y2=5.397
r114 98 101 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.08 $Y=5.397
+ $X2=4.42 $Y2=5.397
r115 94 97 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.215 $Y=3.205
+ $X2=4.215 $Y2=4.565
r116 92 121 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.215 $Y=5.245
+ $X2=4.215 $Y2=5.397
r117 92 97 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.215 $Y=5.245
+ $X2=4.215 $Y2=4.565
r118 89 91 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=5.397
+ $X2=3.74 $Y2=5.397
r119 87 120 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=5.397
+ $X2=2.465 $Y2=5.397
r120 87 89 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=2.55 $Y=5.397
+ $X2=3.06 $Y2=5.397
r121 86 121 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=5.397
+ $X2=4.215 $Y2=5.397
r122 86 91 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=4.13 $Y=5.397
+ $X2=3.74 $Y2=5.397
r123 82 85 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.465 $Y=3.545
+ $X2=2.465 $Y2=4.565
r124 80 120 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.465 $Y=5.245
+ $X2=2.465 $Y2=5.397
r125 80 85 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.465 $Y=5.245
+ $X2=2.465 $Y2=4.565
r126 77 79 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=5.397
+ $X2=1.7 $Y2=5.397
r127 75 118 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=5.397
+ $X2=0.715 $Y2=5.397
r128 75 77 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=0.8 $Y=5.397
+ $X2=1.02 $Y2=5.397
r129 74 120 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=5.397
+ $X2=2.465 $Y2=5.397
r130 74 79 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=5.397
+ $X2=1.7 $Y2=5.397
r131 70 73 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.715 $Y=3.545
+ $X2=0.715 $Y2=4.565
r132 68 118 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.715 $Y=5.245
+ $X2=0.715 $Y2=5.397
r133 68 73 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.715 $Y=5.245
+ $X2=0.715 $Y2=4.565
r134 65 128 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r135 63 118 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=5.397
+ $X2=0.715 $Y2=5.397
r136 63 65 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.63 $Y=5.397
+ $X2=0.34 $Y2=5.397
r137 61 125 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=5.245 $X2=6.46 $Y2=5.33
r138 61 111 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=5.245 $X2=5.78 $Y2=5.33
r139 61 123 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=5.245 $X2=5.1 $Y2=5.33
r140 61 101 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=5.245 $X2=4.42 $Y2=5.33
r141 61 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r142 61 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r143 61 120 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r144 61 79 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r145 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r146 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r147 5 114 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=3.565 $X2=6.545 $Y2=4.565
r148 4 107 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=2.825 $X2=5.165 $Y2=4.565
r149 4 104 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=2.825 $X2=5.165 $Y2=3.545
r150 3 97 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.075
+ $Y=2.825 $X2=4.215 $Y2=4.565
r151 3 94 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=4.075
+ $Y=2.825 $X2=4.215 $Y2=3.205
r152 2 85 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=2.825 $X2=2.465 $Y2=4.565
r153 2 82 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=2.825 $X2=2.465 $Y2=3.545
r154 1 73 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.825 $X2=0.715 $Y2=4.565
r155 1 70 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.825 $X2=0.715 $Y2=3.545
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%A_75_292# 1 3 13 17 20 22 23 28 29 30 31
+ 32 34 37 41 46 47 50
c86 29 0 1.29912e-19 $X=1.405 $Y=1.505
c87 28 0 1.59851e-19 $X=0.625 $Y=2.84
c88 22 0 5.41559e-20 $X=0.51 $Y=2.505
r89 49 50 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.582 $Y=0.985
+ $X2=1.582 $Y2=1.155
r90 46 48 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.505
+ $X2=0.567 $Y2=2.67
r91 46 47 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.505
+ $X2=0.567 $Y2=2.34
r92 41 43 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=1.59 $Y=3.205
+ $X2=1.59 $Y2=4.565
r93 39 41 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=3.115 $X2=1.59
+ $Y2=3.205
r94 37 49 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.59 $Y=0.865
+ $X2=1.59 $Y2=0.985
r95 34 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.49 $Y=1.42
+ $X2=1.49 $Y2=1.155
r96 31 39 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=1.42 $Y=2.925
+ $X2=1.59 $Y2=3.115
r97 31 32 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.42 $Y=2.925
+ $X2=0.71 $Y2=2.925
r98 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.505
+ $X2=1.49 $Y2=1.42
r99 29 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.405 $Y=1.505
+ $X2=0.71 $Y2=1.505
r100 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=2.84
+ $X2=0.71 $Y2=2.925
r101 28 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.625 $Y=2.84
+ $X2=0.625 $Y2=2.67
r102 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.59
+ $X2=0.71 $Y2=1.505
r103 25 47 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.625 $Y=1.59
+ $X2=0.625 $Y2=2.34
r104 22 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=2.505 $X2=0.51 $Y2=2.505
r105 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.505
+ $X2=0.51 $Y2=2.67
r106 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.505
+ $X2=0.51 $Y2=2.34
r107 20 23 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.45 $Y=1.61
+ $X2=0.45 $Y2=2.34
r108 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.475 $Y=1.46
+ $X2=0.475 $Y2=1.61
r109 17 24 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=0.5 $Y=3.825
+ $X2=0.5 $Y2=2.67
r110 13 19 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.5 $Y=0.945
+ $X2=0.5 $Y2=1.46
r111 3 43 240 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=1.365
+ $Y=2.825 $X2=1.59 $Y2=4.565
r112 3 41 240 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=2 $X=1.365
+ $Y=2.825 $X2=1.59 $Y2=3.205
r113 1 37 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.575 $X2=1.59 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%D 3 7 10 14 19
c43 19 0 1.41836e-19 $X=0.99 $Y=1.96
c44 10 0 1.12321e-19 $X=0.99 $Y=1.96
r45 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=1.96
+ $X2=0.99 $Y2=1.96
r46 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.96 $X2=0.99 $Y2=1.96
r47 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.96
+ $X2=0.99 $Y2=2.125
r48 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.96
+ $X2=0.99 $Y2=1.795
r49 7 12 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=0.93 $Y=3.825
+ $X2=0.93 $Y2=2.125
r50 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.93 $Y=0.945
+ $X2=0.93 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c213 55 0 6.79641e-20 $X=3.185 $Y=2.33
c214 48 0 1.98654e-19 $X=1.83 $Y=1.59
c215 44 0 1.86602e-19 $X=1.745 $Y=2.33
c216 30 0 1.29912e-19 $X=1.83 $Y=1.425
c217 25 0 1.41836e-19 $X=1.35 $Y=2.505
r218 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.725 $Y=2.33
+ $X2=3.58 $Y2=2.33
r219 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.43 $Y=2.33
+ $X2=4.575 $Y2=2.33
r220 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=4.43 $Y=2.33
+ $X2=3.725 $Y2=2.33
r221 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.495 $Y=2.33
+ $X2=1.35 $Y2=2.33
r222 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.435 $Y=2.33
+ $X2=3.58 $Y2=2.33
r223 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=3.435 $Y=2.33
+ $X2=1.495 $Y2=2.33
r224 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.33
+ $X2=3.58 $Y2=2.33
r225 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.58 $Y=2.33
+ $X2=3.58 $Y2=2.505
r226 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.35 $Y=2.33
+ $X2=1.35 $Y2=2.33
r227 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.35 $Y=2.33
+ $X2=1.35 $Y2=2.505
r228 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.575 $Y=2.33
+ $X2=4.575 $Y2=2.33
r229 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.33
+ $X2=4.575 $Y2=2.505
r230 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.33
+ $X2=3.58 $Y2=2.33
r231 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.495 $Y=2.33
+ $X2=3.185 $Y2=2.33
r232 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.245
+ $X2=3.185 $Y2=2.33
r233 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.1 $Y=2.245
+ $X2=3.1 $Y2=1.59
r234 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.83 $Y=2.245
+ $X2=1.83 $Y2=1.59
r235 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.33
+ $X2=1.35 $Y2=2.33
r236 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=2.33
+ $X2=1.83 $Y2=2.245
r237 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.745 $Y=2.33
+ $X2=1.435 $Y2=2.33
r238 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=2.505 $X2=4.575 $Y2=2.505
r239 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=4.457 $Y=1.425
+ $X2=4.457 $Y2=1.575
r240 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=2.505 $X2=3.58 $Y2=2.505
r241 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=2.505
+ $X2=3.58 $Y2=2.67
r242 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.59 $X2=3.1 $Y2=1.59
r243 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.59
+ $X2=3.1 $Y2=1.425
r244 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.59 $X2=1.83 $Y2=1.59
r245 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.59
+ $X2=1.83 $Y2=1.425
r246 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=2.505 $X2=1.35 $Y2=2.505
r247 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=2.505
+ $X2=1.35 $Y2=2.67
r248 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=4.485 $Y=2.34
+ $X2=4.532 $Y2=2.505
r249 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.485 $Y=2.34
+ $X2=4.485 $Y2=1.575
r250 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=4.43 $Y=2.67
+ $X2=4.532 $Y2=2.505
r251 18 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=4.43 $Y=2.67
+ $X2=4.43 $Y2=3.825
r252 17 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.43 $Y=0.945
+ $X2=4.43 $Y2=1.425
r253 13 39 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=3.64 $Y=3.825
+ $X2=3.64 $Y2=2.67
r254 10 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.04 $Y=0.945
+ $X2=3.04 $Y2=1.425
r255 7 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.89 $Y=0.945
+ $X2=1.89 $Y2=1.425
r256 3 27 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=1.29 $Y=3.825
+ $X2=1.29 $Y2=2.67
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%A_32_115# 1 3 11 15 17 18 21 22 27 31 34
+ 37 41 47 52 56 61 62 63 68
c116 47 0 1.5821e-19 $X=2.42 $Y=2.505
c117 31 0 6.36774e-20 $X=2.68 $Y=3.825
c118 22 0 1.86602e-19 $X=2.325 $Y=2.505
c119 21 0 6.79641e-20 $X=2.605 $Y=2.505
c120 15 0 6.36774e-20 $X=2.25 $Y=3.825
r121 63 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.43 $Y=1.59
+ $X2=0.285 $Y2=1.59
r122 62 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.185 $Y=1.59
+ $X2=2.33 $Y2=1.59
r123 62 63 1.68986 $w=1.7e-07 $l=1.755e-06 $layer=MET1_cond $X=2.185 $Y=1.59
+ $X2=0.43 $Y2=1.59
r124 59 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.33 $Y=1.59
+ $X2=2.33 $Y2=1.59
r125 59 61 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=2.33 $Y=1.55 $X2=2.42
+ $Y2=1.55
r126 54 56 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=3
+ $X2=0.285 $Y2=3
r127 52 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.285 $Y=1.59
+ $X2=0.285 $Y2=1.59
r128 49 52 4.81931 $w=2.73e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=1.537
+ $X2=0.285 $Y2=1.537
r129 45 61 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.42 $Y=1.675
+ $X2=2.42 $Y2=1.55
r130 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.42 $Y=1.675
+ $X2=2.42 $Y2=2.505
r131 41 43 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.285 $Y=3.205
+ $X2=0.285 $Y2=4.565
r132 39 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=3.085
+ $X2=0.285 $Y2=3
r133 39 41 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.285 $Y=3.085
+ $X2=0.285 $Y2=3.205
r134 35 52 3.55113 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.285 $Y=1.4
+ $X2=0.285 $Y2=1.537
r135 35 37 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.285 $Y=1.4
+ $X2=0.285 $Y2=0.865
r136 34 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=2.915
+ $X2=0.17 $Y2=3
r137 33 49 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.17 $Y=1.675
+ $X2=0.17 $Y2=1.537
r138 33 34 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=0.17 $Y=1.675
+ $X2=0.17 $Y2=2.915
r139 29 31 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=2.68 $Y=2.64
+ $X2=2.68 $Y2=3.825
r140 25 27 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.68 $Y=1.455
+ $X2=2.68 $Y2=0.945
r141 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=2.505 $X2=2.42 $Y2=2.505
r142 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=2.505
+ $X2=2.42 $Y2=2.505
r143 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=2.505
+ $X2=2.68 $Y2=2.64
r144 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=2.505
+ $X2=2.42 $Y2=2.505
r145 20 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.59 $X2=2.42 $Y2=1.59
r146 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=1.59
+ $X2=2.42 $Y2=1.59
r147 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=1.59
+ $X2=2.68 $Y2=1.455
r148 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=1.59
+ $X2=2.42 $Y2=1.59
r149 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=2.64
+ $X2=2.325 $Y2=2.505
r150 13 15 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=2.25 $Y=2.64
+ $X2=2.25 $Y2=3.825
r151 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=1.455
+ $X2=2.325 $Y2=1.59
r152 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.25 $Y=1.455
+ $X2=2.25 $Y2=0.945
r153 3 43 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.825 $X2=0.285 $Y2=4.565
r154 3 41 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.825 $X2=0.285 $Y2=3.205
r155 1 37 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%A_243_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c174 35 0 1.98654e-19 $X=1.41 $Y=1.5
c175 18 0 1.12321e-19 $X=1.89 $Y=3.825
r176 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=2.925
+ $X2=4.915 $Y2=2.925
r177 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=1.93
+ $X2=4.915 $Y2=1.93
r178 60 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.84
+ $X2=4.915 $Y2=2.925
r179 59 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.015
+ $X2=4.915 $Y2=1.93
r180 59 60 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.915 $Y=2.015
+ $X2=4.915 $Y2=2.84
r181 55 57 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.645 $Y=3.205
+ $X2=4.645 $Y2=4.565
r182 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=3.01
+ $X2=4.645 $Y2=2.925
r183 53 55 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.645 $Y=3.01
+ $X2=4.645 $Y2=3.205
r184 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.845
+ $X2=4.645 $Y2=1.93
r185 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.675
+ $X2=4.645 $Y2=1.59
r186 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.645 $Y=1.675
+ $X2=4.645 $Y2=1.845
r187 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.505
+ $X2=4.645 $Y2=1.59
r188 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.645 $Y=1.505
+ $X2=4.645 $Y2=0.865
r189 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=1.59
+ $X2=4.645 $Y2=1.59
r190 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.56 $Y=1.59
+ $X2=3.58 $Y2=1.59
r191 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.59 $X2=3.58 $Y2=1.59
r192 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.59
+ $X2=3.58 $Y2=1.755
r193 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.59
+ $X2=3.58 $Y2=1.425
r194 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.29 $Y=1.5
+ $X2=1.41 $Y2=1.5
r195 32 41 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.64 $Y=0.945
+ $X2=3.64 $Y2=1.425
r196 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.52 $Y=1.965
+ $X2=3.52 $Y2=1.755
r197 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.115 $Y=2.04
+ $X2=3.04 $Y2=2.04
r198 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.445 $Y=2.04
+ $X2=3.52 $Y2=1.965
r199 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.445 $Y=2.04
+ $X2=3.115 $Y2=2.04
r200 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.04 $Y=2.115
+ $X2=3.04 $Y2=2.04
r201 22 24 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=3.04 $Y=2.115
+ $X2=3.04 $Y2=3.825
r202 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=2.04
+ $X2=1.89 $Y2=2.04
r203 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.965 $Y=2.04
+ $X2=3.04 $Y2=2.04
r204 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.965 $Y=2.04
+ $X2=1.965 $Y2=2.04
r205 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=2.115
+ $X2=1.89 $Y2=2.04
r206 16 18 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=1.89 $Y=2.115
+ $X2=1.89 $Y2=3.825
r207 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=2.04
+ $X2=1.89 $Y2=2.04
r208 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.815 $Y=2.04
+ $X2=1.485 $Y2=2.04
r209 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.965
+ $X2=1.485 $Y2=2.04
r210 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.575
+ $X2=1.41 $Y2=1.5
r211 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.41 $Y=1.575
+ $X2=1.41 $Y2=1.965
r212 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.425
+ $X2=1.29 $Y2=1.5
r213 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.29 $Y=1.425
+ $X2=1.29 $Y2=0.945
r214 3 57 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=2.825 $X2=4.645 $Y2=4.565
r215 3 55 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=2.825 $X2=4.645 $Y2=3.205
r216 1 49 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.575 $X2=4.645 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%A_785_89# 1 3 11 15 23 27 30 34 35 38 39
+ 40 42 48 52 58 61 62 63 68
c134 39 0 8.77106e-20 $X=6.305 $Y=2.595
c135 34 0 2.20654e-19 $X=6.215 $Y=1.93
r136 63 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.205 $Y=1.93
+ $X2=4.06 $Y2=1.93
r137 62 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.07 $Y=1.93
+ $X2=6.215 $Y2=1.93
r138 62 63 1.79578 $w=1.7e-07 $l=1.865e-06 $layer=MET1_cond $X=6.07 $Y=1.93
+ $X2=4.205 $Y2=1.93
r139 58 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=1.93
+ $X2=6.215 $Y2=1.93
r140 56 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=1.93
+ $X2=5.595 $Y2=1.93
r141 56 58 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.68 $Y=1.93
+ $X2=6.215 $Y2=1.93
r142 52 54 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=5.595 $Y=3.205
+ $X2=5.595 $Y2=4.565
r143 50 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=2.015
+ $X2=5.595 $Y2=1.93
r144 50 52 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.595 $Y=2.015
+ $X2=5.595 $Y2=3.205
r145 46 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.845
+ $X2=5.595 $Y2=1.93
r146 46 48 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.595 $Y=1.845
+ $X2=5.595 $Y2=0.865
r147 42 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.06 $Y=1.93
+ $X2=4.06 $Y2=1.93
r148 39 40 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=2.595
+ $X2=6.305 $Y2=2.745
r149 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=1.39
+ $X2=6.305 $Y2=1.54
r150 36 39 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.28 $Y=2.095
+ $X2=6.28 $Y2=2.595
r151 35 38 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.28 $Y=1.765
+ $X2=6.28 $Y2=1.54
r152 34 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.93 $X2=6.215 $Y2=1.93
r153 34 36 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.217 $Y=1.93
+ $X2=6.217 $Y2=2.095
r154 34 35 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.217 $Y=1.93
+ $X2=6.217 $Y2=1.765
r155 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.93 $X2=4.06 $Y2=1.93
r156 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.93
+ $X2=4.06 $Y2=2.095
r157 30 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.93
+ $X2=4.06 $Y2=1.765
r158 27 40 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=6.33 $Y=4.195
+ $X2=6.33 $Y2=2.745
r159 23 37 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.33 $Y=0.835
+ $X2=6.33 $Y2=1.39
r160 15 32 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=4 $Y=3.825 $X2=4
+ $Y2=2.095
r161 11 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4 $Y=0.945 $X2=4
+ $Y2=1.765
r162 3 54 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=5.455
+ $Y=2.825 $X2=5.595 $Y2=4.565
r163 3 52 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=5.455
+ $Y=2.825 $X2=5.595 $Y2=3.205
r164 1 48 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.575 $X2=5.595 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%A_623_115# 1 3 9 11 14 19 24 25 26 27 28
+ 31 35 40 44 45 50
c115 45 0 1.5821e-19 $X=2.905 $Y=1.59
c116 24 0 1.57671e-19 $X=2.76 $Y=1.59
r117 45 47 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.905 $Y=1.59
+ $X2=2.76 $Y2=1.59
r118 44 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.59
+ $X2=5.175 $Y2=1.59
r119 44 45 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=5.03 $Y=1.59
+ $X2=2.905 $Y2=1.59
r120 40 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.59
+ $X2=5.175 $Y2=1.59
r121 35 37 34.5733 $w=3.38e-07 $l=1.02e-06 $layer=LI1_cond $X=3.34 $Y=3.545
+ $X2=3.34 $Y2=4.565
r122 33 35 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=3.34 $Y=3.01
+ $X2=3.34 $Y2=3.545
r123 29 31 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=3.34 $Y=1.085
+ $X2=3.34 $Y2=0.865
r124 27 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=2.925
+ $X2=3.34 $Y2=3.01
r125 27 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=2.925
+ $X2=2.845 $Y2=2.925
r126 25 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=1.17
+ $X2=3.34 $Y2=1.085
r127 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=1.17
+ $X2=2.845 $Y2=1.17
r128 24 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.76 $Y=1.59
+ $X2=2.76 $Y2=1.59
r129 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=2.84
+ $X2=2.845 $Y2=2.925
r130 22 24 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.76 $Y=2.84
+ $X2=2.76 $Y2=1.59
r131 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=1.255
+ $X2=2.845 $Y2=1.17
r132 21 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.76 $Y=1.255
+ $X2=2.76 $Y2=1.59
r133 17 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.59 $X2=5.175 $Y2=1.59
r134 17 19 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.175 $Y=1.59
+ $X2=5.38 $Y2=1.59
r135 12 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.755
+ $X2=5.38 $Y2=1.59
r136 12 14 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=5.38 $Y=1.755
+ $X2=5.38 $Y2=3.825
r137 9 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.425
+ $X2=5.38 $Y2=1.59
r138 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.38 $Y=1.425
+ $X2=5.38 $Y2=0.945
r139 3 37 300 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=3.115
+ $Y=2.825 $X2=3.34 $Y2=4.565
r140 3 35 300 $w=1.7e-07 $l=8.24864e-07 $layer=licon1_PDIFF $count=2 $X=3.115
+ $Y=2.825 $X2=3.34 $Y2=3.545
r141 1 31 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.575 $X2=3.34 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c77 42 0 8.77106e-20 $X=6.12 $Y=2.7
c78 33 0 9.99996e-20 $X=6.615 $Y=2.505
c79 31 0 1.20654e-19 $X=6.615 $Y=1.59
r80 40 42 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=6.115 $Y=2.7
+ $X2=6.12 $Y2=2.7
r81 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.7 $Y=2.42 $X2=6.7
+ $Y2=2.135
r82 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.7 $Y=1.675 $X2=6.7
+ $Y2=2.135
r83 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=2.505
+ $X2=6.7 $Y2=2.42
r84 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=2.505
+ $X2=6.2 $Y2=2.505
r85 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=1.59
+ $X2=6.7 $Y2=1.675
r86 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=1.59
+ $X2=6.2 $Y2=1.59
r87 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.115 $Y=2.7
+ $X2=6.115 $Y2=2.7
r88 27 29 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=6.115 $Y=2.7
+ $X2=6.115 $Y2=4.565
r89 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=2.59
+ $X2=6.2 $Y2=2.505
r90 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.115 $Y=2.59
+ $X2=6.115 $Y2=2.7
r91 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=1.505
+ $X2=6.2 $Y2=1.59
r92 21 23 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.115 $Y=1.505
+ $X2=6.115 $Y2=0.74
r93 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=2.135 $X2=6.7 $Y2=2.135
r94 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.135
+ $X2=6.7 $Y2=2.3
r95 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.135
+ $X2=6.7 $Y2=1.97
r96 15 20 971.691 $w=1.5e-07 $l=1.895e-06 $layer=POLY_cond $X=6.76 $Y=4.195
+ $X2=6.76 $Y2=2.3
r97 11 19 581.989 $w=1.5e-07 $l=1.135e-06 $layer=POLY_cond $X=6.76 $Y=0.835
+ $X2=6.76 $Y2=1.97
r98 3 29 600 $w=1.7e-07 $l=1.06066e-06 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=3.565 $X2=6.115 $Y2=4.565
r99 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.575 $X2=6.115 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__DFF_L%Q 1 3 11 15 18 21 25 28
r22 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=3.027
+ $X2=7.09 $Y2=3.027
r23 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.97 $Y=3.07
+ $X2=6.97 $Y2=3.07
r24 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=6.97 $Y=3.027
+ $X2=6.975 $Y2=3.027
r25 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=1.255
+ $X2=7.09 $Y2=1.255
r26 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.09 $Y=2.9 $X2=7.09
+ $Y2=3.027
r27 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.34
+ $X2=7.09 $Y2=1.255
r28 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=7.09 $Y=1.34
+ $X2=7.09 $Y2=2.9
r29 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=6.975 $Y=3.155
+ $X2=6.975 $Y2=3.027
r30 13 15 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=6.975 $Y=3.155
+ $X2=6.975 $Y2=4.565
r31 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=1.17
+ $X2=6.975 $Y2=1.255
r32 9 11 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.975 $Y=1.17
+ $X2=6.975 $Y2=0.74
r33 3 15 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=6.835
+ $Y=3.565 $X2=6.975 $Y2=4.565
r34 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.575 $X2=6.975 $Y2=0.74
.ends

