* File: sky130_osu_sc_15T_hs__tnbufi_1.spice
* Created: Fri Nov 12 14:33:47 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__tnbufi_1.pex.spice"
.subckt sky130_osu_sc_15T_hs__tnbufi_1  GND VDD OE A Y
* 
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_OE_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1001 A_196_115# N_A_27_115#_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.64 AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g A_196_115# N_GND_M1003_b NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75001
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VDD_M1004_d N_OE_M1004_g N_A_27_115#_M1004_s N_VDD_M1004_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1002 A_196_565# N_OE_M1002_g N_VDD_M1004_d N_VDD_M1004_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.5 A=0.3 P=4.3 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g A_196_565# N_VDD_M1004_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.21 PD=4.53 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1004_b NWDIODE A=5.664 P=9.74
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__tnbufi_1.pxi.spice"
*
.ends
*
*
