* File: sky130_osu_sc_18T_ls__oai21_l.pex.spice
* Created: Fri Nov 12 14:18:52 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%GND 1 17 19 26 35 38
r37 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r38 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r39 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r40 24 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r41 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r42 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r43 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r44 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r45 1 26 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%VDD 1 13 15 21 28 31 34
r26 31 34 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r27 28 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r28 21 24 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.05 $Y=4.475
+ $X2=1.05 $Y2=5.835
r29 19 28 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.05 $Y=6.355
+ $X2=1.05 $Y2=6.507
r30 19 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=6.355
+ $X2=1.05 $Y2=5.835
r31 15 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=6.507
+ $X2=1.05 $Y2=6.507
r32 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=6.507
+ $X2=0.34 $Y2=6.507
r33 13 28 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r34 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r35 1 24 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=3.085 $X2=1.05 $Y2=5.835
r36 1 21 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=3.085 $X2=1.05 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%A0 3 5 8 12 15 16 19 25
r37 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.415 $Y=3.33
+ $X2=0.415 $Y2=3.33
r38 19 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.415 $Y=2.76
+ $X2=0.415 $Y2=3.33
r39 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=2.76 $X2=0.415 $Y2=2.76
r40 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.76
+ $X2=0.415 $Y2=2.925
r41 15 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.76
+ $X2=0.415 $Y2=2.595
r42 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=0.355 $Y=1.775
+ $X2=0.475 $Y2=1.775
r43 8 17 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.925
r44 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.775
r45 3 5 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.075
r46 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.355 $Y=1.85
+ $X2=0.355 $Y2=1.775
r47 1 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.355 $Y=1.85
+ $X2=0.355 $Y2=2.595
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%A1 3 7 10 15 18 22
r55 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.895 $Y=2.96
+ $X2=0.895 $Y2=2.96
r56 18 19 5.0779 $w=2.18e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.96 $X2=0.87
+ $Y2=2.875
r57 15 19 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.845 $Y=2.22
+ $X2=0.845 $Y2=2.875
r58 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.22 $X2=0.845 $Y2=2.22
r59 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.845 $Y=2.22
+ $X2=0.845 $Y2=2.355
r60 10 11 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.845 $Y=2.22
+ $X2=0.845 $Y2=2.085
r61 7 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.085
r62 3 12 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=0.835 $Y=4.585
+ $X2=0.835 $Y2=2.355
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%B0 1 3 7 13 15 17 20
r52 15 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.285 $Y=1.88
+ $X2=1.395 $Y2=1.88
r53 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.59 $X2=1.2
+ $Y2=2.59
r54 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=1.965
+ $X2=1.285 $Y2=1.88
r55 11 13 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.2 $Y=1.965
+ $X2=1.2 $Y2=2.59
r56 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.88 $X2=1.395 $Y2=1.88
r57 5 10 38.8629 $w=2.72e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.335 $Y=1.715
+ $X2=1.39 $Y2=1.88
r58 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.335 $Y=1.715
+ $X2=1.335 $Y2=1.075
r59 1 10 38.8629 $w=2.72e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.325 $Y=2.045
+ $X2=1.39 $Y2=1.88
r60 1 3 1558.81 $w=1.5e-07 $l=3.04e-06 $layer=POLY_cond $X=1.325 $Y=2.045
+ $X2=1.325 $Y2=5.085
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%Y 1 3 4 15 19 20 23 27 32 37 41 42 47
r57 41 42 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.54 $Y=2.22
+ $X2=1.54 $Y2=2.105
r58 38 47 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r59 38 42 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.105
r60 35 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r61 32 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.55 $Y=0.82
+ $X2=1.55 $Y2=1.48
r62 27 29 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.54 $Y=4.475
+ $X2=1.54 $Y2=5.835
r63 25 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.755
+ $X2=1.54 $Y2=3.67
r64 25 27 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.54 $Y=3.755
+ $X2=1.54 $Y2=4.475
r65 23 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.54 $Y=2.22
+ $X2=1.54 $Y2=2.22
r66 21 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.585
+ $X2=1.54 $Y2=3.67
r67 21 23 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.54 $Y=3.585
+ $X2=1.54 $Y2=2.22
r68 19 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=3.67
+ $X2=1.54 $Y2=3.67
r69 19 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.455 $Y=3.67
+ $X2=0.345 $Y2=3.67
r70 15 17 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r71 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.755
+ $X2=0.345 $Y2=3.67
r72 13 15 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.26 $Y=3.755
+ $X2=0.26 $Y2=4.135
r73 4 29 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=4.085 $X2=1.54 $Y2=5.835
r74 4 27 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=4.085 $X2=1.54 $Y2=4.475
r75 3 17 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r76 3 15 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
r77 1 32 91 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.82
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__OAI21_L%A_27_115# 1 2 11 13 14 17
r14 15 17 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=0.825
r15 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.42
+ $X2=1.12 $Y2=1.335
r16 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.42
+ $X2=0.345 $Y2=1.42
r17 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.335
+ $X2=0.345 $Y2=1.42
r18 9 11 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.26 $Y=1.335
+ $X2=0.26 $Y2=0.825
r19 2 17 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r20 1 11 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

