* File: sky130_osu_sc_18T_hs__buf_8.pxi.spice
* Created: Fri Nov 12 13:48:22 2021
* 
x_PM_SKY130_OSU_SC_18T_HS__BUF_8%GND N_GND_M1006_d N_GND_M1003_s N_GND_M1010_s
+ N_GND_M1014_s N_GND_M1017_s N_GND_M1006_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p
+ N_GND_c_15_p N_GND_c_24_p N_GND_c_30_p N_GND_c_37_p N_GND_c_44_p N_GND_c_51_p
+ N_GND_c_57_p GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_HS__BUF_8%GND
x_PM_SKY130_OSU_SC_18T_HS__BUF_8%VDD N_VDD_M1004_d N_VDD_M1002_s N_VDD_M1008_s
+ N_VDD_M1012_s N_VDD_M1016_s N_VDD_M1004_b N_VDD_c_121_p N_VDD_c_122_p
+ N_VDD_c_131_p N_VDD_c_136_p N_VDD_c_143_p N_VDD_c_148_p N_VDD_c_154_p
+ N_VDD_c_159_p N_VDD_c_165_p N_VDD_c_170_p VDD N_VDD_c_123_p
+ PM_SKY130_OSU_SC_18T_HS__BUF_8%VDD
x_PM_SKY130_OSU_SC_18T_HS__BUF_8%A N_A_M1006_g N_A_M1004_g N_A_c_207_n
+ N_A_c_208_n A PM_SKY130_OSU_SC_18T_HS__BUF_8%A
x_PM_SKY130_OSU_SC_18T_HS__BUF_8%A_27_115# N_A_27_115#_M1006_s
+ N_A_27_115#_M1004_s N_A_27_115#_M1001_g N_A_27_115#_c_311_n
+ N_A_27_115#_M1000_g N_A_27_115#_c_246_n N_A_27_115#_M1003_g
+ N_A_27_115#_c_315_n N_A_27_115#_M1002_g N_A_27_115#_c_251_n
+ N_A_27_115#_c_253_n N_A_27_115#_c_254_n N_A_27_115#_c_255_n
+ N_A_27_115#_M1007_g N_A_27_115#_c_323_n N_A_27_115#_M1005_g
+ N_A_27_115#_c_260_n N_A_27_115#_c_261_n N_A_27_115#_M1010_g
+ N_A_27_115#_c_328_n N_A_27_115#_M1008_g N_A_27_115#_c_266_n
+ N_A_27_115#_c_268_n N_A_27_115#_M1011_g N_A_27_115#_c_273_n
+ N_A_27_115#_c_334_n N_A_27_115#_M1009_g N_A_27_115#_c_274_n
+ N_A_27_115#_c_275_n N_A_27_115#_M1014_g N_A_27_115#_c_339_n
+ N_A_27_115#_M1012_g N_A_27_115#_c_280_n N_A_27_115#_c_282_n
+ N_A_27_115#_M1015_g N_A_27_115#_c_345_n N_A_27_115#_M1013_g
+ N_A_27_115#_c_287_n N_A_27_115#_c_288_n N_A_27_115#_M1017_g
+ N_A_27_115#_c_350_n N_A_27_115#_M1016_g N_A_27_115#_c_293_n
+ N_A_27_115#_c_294_n N_A_27_115#_c_295_n N_A_27_115#_c_296_n
+ N_A_27_115#_c_297_n N_A_27_115#_c_298_n N_A_27_115#_c_299_n
+ N_A_27_115#_c_300_n N_A_27_115#_c_301_n N_A_27_115#_c_302_n
+ N_A_27_115#_c_303_n N_A_27_115#_c_306_n N_A_27_115#_c_307_n
+ N_A_27_115#_c_309_n N_A_27_115#_c_310_n
+ PM_SKY130_OSU_SC_18T_HS__BUF_8%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__BUF_8%Y N_Y_M1001_d N_Y_M1007_d N_Y_M1011_d
+ N_Y_M1015_d N_Y_M1000_d N_Y_M1005_d N_Y_M1009_d N_Y_M1013_d N_Y_c_474_n
+ N_Y_c_517_n N_Y_c_478_n N_Y_c_520_n N_Y_c_483_n N_Y_c_523_n N_Y_c_488_n
+ N_Y_c_526_n N_Y_c_492_n N_Y_c_495_n Y N_Y_c_497_n N_Y_c_530_n N_Y_c_499_n
+ N_Y_c_500_n N_Y_c_502_n N_Y_c_532_n N_Y_c_505_n N_Y_c_506_n N_Y_c_507_n
+ N_Y_c_509_n N_Y_c_535_n N_Y_c_512_n N_Y_c_513_n N_Y_c_516_n
+ PM_SKY130_OSU_SC_18T_HS__BUF_8%Y
cc_1 N_GND_M1006_b N_A_M1006_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1006_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1006_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_A_M1006_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.475 $Y2=1.075
cc_5 N_GND_M1006_b N_A_M1004_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_6 N_GND_M1006_b N_A_c_207_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_7 N_GND_M1006_b N_A_c_208_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_8 N_GND_M1006_b N_A_27_115#_M1001_g 0.0207501f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=1.075
cc_9 N_GND_c_3_p N_A_27_115#_M1001_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=1.075
cc_10 N_GND_c_10_p N_A_27_115#_M1001_g 0.00606474f $X=1.465 $Y=0.152 $X2=0.905
+ $Y2=1.075
cc_11 N_GND_c_4_p N_A_27_115#_M1001_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.905
+ $Y2=1.075
cc_12 N_GND_M1006_b N_A_27_115#_c_246_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.86
cc_13 N_GND_M1006_b N_A_27_115#_M1003_g 0.020212f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_14 N_GND_c_10_p N_A_27_115#_M1003_g 0.00606474f $X=1.465 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_15 N_GND_c_15_p N_A_27_115#_M1003_g 0.00356864f $X=1.55 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_16 N_GND_c_4_p N_A_27_115#_M1003_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_M1006_b N_A_27_115#_c_251_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.845
cc_18 N_GND_c_15_p N_A_27_115#_c_251_n 0.00256938f $X=1.55 $Y=0.825 $X2=1.69
+ $Y2=1.845
cc_19 N_GND_M1006_b N_A_27_115#_c_253_n 0.0429274f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.845
cc_20 N_GND_M1006_b N_A_27_115#_c_254_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.935
cc_21 N_GND_M1006_b N_A_27_115#_c_255_n 0.0196789f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.935
cc_22 N_GND_M1006_b N_A_27_115#_M1007_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_23 N_GND_c_15_p N_A_27_115#_M1007_g 0.00356864f $X=1.55 $Y=0.825 $X2=1.765
+ $Y2=1.075
cc_24 N_GND_c_24_p N_A_27_115#_M1007_g 0.00606474f $X=2.325 $Y=0.152 $X2=1.765
+ $Y2=1.075
cc_25 N_GND_c_4_p N_A_27_115#_M1007_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.765
+ $Y2=1.075
cc_26 N_GND_M1006_b N_A_27_115#_c_260_n 0.0195339f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.845
cc_27 N_GND_M1006_b N_A_27_115#_c_261_n 0.0107618f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.935
cc_28 N_GND_M1006_b N_A_27_115#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.075
cc_29 N_GND_c_24_p N_A_27_115#_M1010_g 0.00606474f $X=2.325 $Y=0.152 $X2=2.195
+ $Y2=1.075
cc_30 N_GND_c_30_p N_A_27_115#_M1010_g 0.00356864f $X=2.41 $Y=0.825 $X2=2.195
+ $Y2=1.075
cc_31 N_GND_c_4_p N_A_27_115#_M1010_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.195
+ $Y2=1.075
cc_32 N_GND_M1006_b N_A_27_115#_c_266_n 0.0165886f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.845
cc_33 N_GND_c_30_p N_A_27_115#_c_266_n 0.00256938f $X=2.41 $Y=0.825 $X2=2.55
+ $Y2=1.845
cc_34 N_GND_M1006_b N_A_27_115#_c_268_n 0.0109555f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.935
cc_35 N_GND_M1006_b N_A_27_115#_M1011_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.075
cc_36 N_GND_c_30_p N_A_27_115#_M1011_g 0.00356864f $X=2.41 $Y=0.825 $X2=2.625
+ $Y2=1.075
cc_37 N_GND_c_37_p N_A_27_115#_M1011_g 0.00606474f $X=3.185 $Y=0.152 $X2=2.625
+ $Y2=1.075
cc_38 N_GND_c_4_p N_A_27_115#_M1011_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.625
+ $Y2=1.075
cc_39 N_GND_M1006_b N_A_27_115#_c_273_n 0.0668243f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.86
cc_40 N_GND_M1006_b N_A_27_115#_c_274_n 0.0195339f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.845
cc_41 N_GND_M1006_b N_A_27_115#_c_275_n 0.0107618f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.935
cc_42 N_GND_M1006_b N_A_27_115#_M1014_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.075
cc_43 N_GND_c_37_p N_A_27_115#_M1014_g 0.00606474f $X=3.185 $Y=0.152 $X2=3.055
+ $Y2=1.075
cc_44 N_GND_c_44_p N_A_27_115#_M1014_g 0.00356864f $X=3.27 $Y=0.825 $X2=3.055
+ $Y2=1.075
cc_45 N_GND_c_4_p N_A_27_115#_M1014_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.055
+ $Y2=1.075
cc_46 N_GND_M1006_b N_A_27_115#_c_280_n 0.0215078f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.845
cc_47 N_GND_c_44_p N_A_27_115#_c_280_n 0.00256938f $X=3.27 $Y=0.825 $X2=3.41
+ $Y2=1.845
cc_48 N_GND_M1006_b N_A_27_115#_c_282_n 0.0158747f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.935
cc_49 N_GND_M1006_b N_A_27_115#_M1015_g 0.020212f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.075
cc_50 N_GND_c_44_p N_A_27_115#_M1015_g 0.00356864f $X=3.27 $Y=0.825 $X2=3.485
+ $Y2=1.075
cc_51 N_GND_c_51_p N_A_27_115#_M1015_g 0.00606474f $X=4.045 $Y=0.152 $X2=3.485
+ $Y2=1.075
cc_52 N_GND_c_4_p N_A_27_115#_M1015_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.485
+ $Y2=1.075
cc_53 N_GND_M1006_b N_A_27_115#_c_287_n 0.0385034f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.845
cc_54 N_GND_M1006_b N_A_27_115#_c_288_n 0.0221499f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.935
cc_55 N_GND_M1006_b N_A_27_115#_M1017_g 0.0264941f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=1.075
cc_56 N_GND_c_51_p N_A_27_115#_M1017_g 0.00606474f $X=4.045 $Y=0.152 $X2=3.915
+ $Y2=1.075
cc_57 N_GND_c_57_p N_A_27_115#_M1017_g 0.00713292f $X=4.13 $Y=0.825 $X2=3.915
+ $Y2=1.075
cc_58 N_GND_c_4_p N_A_27_115#_M1017_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.915
+ $Y2=1.075
cc_59 N_GND_M1006_b N_A_27_115#_c_293_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.845
cc_60 N_GND_M1006_b N_A_27_115#_c_294_n 0.00890086f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.935
cc_61 N_GND_M1006_b N_A_27_115#_c_295_n 0.0106787f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.845
cc_62 N_GND_M1006_b N_A_27_115#_c_296_n 0.00890086f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.935
cc_63 N_GND_M1006_b N_A_27_115#_c_297_n 0.0023879f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.845
cc_64 N_GND_M1006_b N_A_27_115#_c_298_n 7.16371e-19 $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.935
cc_65 N_GND_M1006_b N_A_27_115#_c_299_n 0.0106787f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.845
cc_66 N_GND_M1006_b N_A_27_115#_c_300_n 0.00890086f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.935
cc_67 N_GND_M1006_b N_A_27_115#_c_301_n 0.0106787f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.845
cc_68 N_GND_M1006_b N_A_27_115#_c_302_n 0.00890086f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.935
cc_69 N_GND_M1006_b N_A_27_115#_c_303_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_70 N_GND_c_2_p N_A_27_115#_c_303_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_71 N_GND_c_4_p N_A_27_115#_c_303_n 0.00476261f $X=3.74 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_72 N_GND_M1006_b N_A_27_115#_c_306_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.455
cc_73 N_GND_M1006_b N_A_27_115#_c_307_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.935
cc_74 N_GND_c_3_p N_A_27_115#_c_307_n 0.00702738f $X=0.69 $Y=0.825 $X2=0.88
+ $Y2=1.935
cc_75 N_GND_M1006_b N_A_27_115#_c_309_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.935
cc_76 N_GND_M1006_b N_A_27_115#_c_310_n 0.00592383f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.935
cc_77 N_GND_M1006_b N_Y_c_474_n 0.00155118f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.825
cc_78 N_GND_c_10_p N_Y_c_474_n 0.00734006f $X=1.465 $Y=0.152 $X2=1.12 $Y2=0.825
cc_79 N_GND_c_15_p N_Y_c_474_n 8.14297e-19 $X=1.55 $Y=0.825 $X2=1.12 $Y2=0.825
cc_80 N_GND_c_4_p N_Y_c_474_n 0.00475776f $X=3.74 $Y=0.19 $X2=1.12 $Y2=0.825
cc_81 N_GND_M1006_b N_Y_c_478_n 0.00155118f $X=-0.045 $Y=0 $X2=1.98 $Y2=0.825
cc_82 N_GND_c_15_p N_Y_c_478_n 8.14297e-19 $X=1.55 $Y=0.825 $X2=1.98 $Y2=0.825
cc_83 N_GND_c_24_p N_Y_c_478_n 0.00754406f $X=2.325 $Y=0.152 $X2=1.98 $Y2=0.825
cc_84 N_GND_c_30_p N_Y_c_478_n 8.14297e-19 $X=2.41 $Y=0.825 $X2=1.98 $Y2=0.825
cc_85 N_GND_c_4_p N_Y_c_478_n 0.00475776f $X=3.74 $Y=0.19 $X2=1.98 $Y2=0.825
cc_86 N_GND_M1006_b N_Y_c_483_n 0.00155118f $X=-0.045 $Y=0 $X2=2.84 $Y2=0.825
cc_87 N_GND_c_30_p N_Y_c_483_n 8.14297e-19 $X=2.41 $Y=0.825 $X2=2.84 $Y2=0.825
cc_88 N_GND_c_37_p N_Y_c_483_n 0.00746708f $X=3.185 $Y=0.152 $X2=2.84 $Y2=0.825
cc_89 N_GND_c_44_p N_Y_c_483_n 8.14297e-19 $X=3.27 $Y=0.825 $X2=2.84 $Y2=0.825
cc_90 N_GND_c_4_p N_Y_c_483_n 0.00475776f $X=3.74 $Y=0.19 $X2=2.84 $Y2=0.825
cc_91 N_GND_M1006_b N_Y_c_488_n 0.00155118f $X=-0.045 $Y=0 $X2=3.7 $Y2=0.825
cc_92 N_GND_c_44_p N_Y_c_488_n 8.14297e-19 $X=3.27 $Y=0.825 $X2=3.7 $Y2=0.825
cc_93 N_GND_c_51_p N_Y_c_488_n 0.00734006f $X=4.045 $Y=0.152 $X2=3.7 $Y2=0.825
cc_94 N_GND_c_4_p N_Y_c_488_n 0.00475776f $X=3.74 $Y=0.19 $X2=3.7 $Y2=0.825
cc_95 N_GND_M1006_b N_Y_c_492_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.595
cc_96 N_GND_c_3_p N_Y_c_492_n 0.00134236f $X=0.69 $Y=0.825 $X2=1.12 $Y2=1.595
cc_97 N_GND_c_15_p N_Y_c_492_n 7.53951e-19 $X=1.55 $Y=0.825 $X2=1.12 $Y2=1.595
cc_98 N_GND_M1006_b N_Y_c_495_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.845
cc_99 N_GND_M1006_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=2.27
cc_100 N_GND_M1003_s N_Y_c_497_n 0.0127884f $X=1.41 $Y=0.575 $X2=1.835 $Y2=1.48
cc_101 N_GND_c_15_p N_Y_c_497_n 0.0142303f $X=1.55 $Y=0.825 $X2=1.835 $Y2=1.48
cc_102 N_GND_M1006_b N_Y_c_499_n 0.0437239f $X=-0.045 $Y=0 $X2=1.98 $Y2=2.845
cc_103 N_GND_M1010_s N_Y_c_500_n 0.0127884f $X=2.27 $Y=0.575 $X2=2.695 $Y2=1.48
cc_104 N_GND_c_30_p N_Y_c_500_n 0.0142303f $X=2.41 $Y=0.825 $X2=2.695 $Y2=1.48
cc_105 N_GND_M1006_b N_Y_c_502_n 0.00409378f $X=-0.045 $Y=0 $X2=2.125 $Y2=1.48
cc_106 N_GND_c_15_p N_Y_c_502_n 7.53951e-19 $X=1.55 $Y=0.825 $X2=2.125 $Y2=1.48
cc_107 N_GND_c_30_p N_Y_c_502_n 7.53951e-19 $X=2.41 $Y=0.825 $X2=2.125 $Y2=1.48
cc_108 N_GND_M1006_b N_Y_c_505_n 0.00560779f $X=-0.045 $Y=0 $X2=2.125 $Y2=2.96
cc_109 N_GND_M1006_b N_Y_c_506_n 0.0575129f $X=-0.045 $Y=0 $X2=2.84 $Y2=2.845
cc_110 N_GND_M1014_s N_Y_c_507_n 0.0127884f $X=3.13 $Y=0.575 $X2=3.555 $Y2=1.48
cc_111 N_GND_c_44_p N_Y_c_507_n 0.0142303f $X=3.27 $Y=0.825 $X2=3.555 $Y2=1.48
cc_112 N_GND_M1006_b N_Y_c_509_n 0.00409378f $X=-0.045 $Y=0 $X2=2.985 $Y2=1.48
cc_113 N_GND_c_30_p N_Y_c_509_n 7.53951e-19 $X=2.41 $Y=0.825 $X2=2.985 $Y2=1.48
cc_114 N_GND_c_44_p N_Y_c_509_n 7.53951e-19 $X=3.27 $Y=0.825 $X2=2.985 $Y2=1.48
cc_115 N_GND_M1006_b N_Y_c_512_n 0.00485078f $X=-0.045 $Y=0 $X2=2.985 $Y2=2.96
cc_116 N_GND_M1006_b N_Y_c_513_n 0.00409378f $X=-0.045 $Y=0 $X2=3.7 $Y2=1.595
cc_117 N_GND_c_44_p N_Y_c_513_n 7.53951e-19 $X=3.27 $Y=0.825 $X2=3.7 $Y2=1.595
cc_118 N_GND_c_57_p N_Y_c_513_n 0.00134236f $X=4.13 $Y=0.825 $X2=3.7 $Y2=1.595
cc_119 N_GND_M1006_b N_Y_c_516_n 0.0800785f $X=-0.045 $Y=0 $X2=3.7 $Y2=2.845
cc_120 N_VDD_M1004_b N_A_M1004_g 0.0245629f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_121 N_VDD_c_121_p N_A_M1004_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_122 N_VDD_c_122_p N_A_M1004_g 0.00354579f $X=0.69 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_123 N_VDD_c_123_p N_A_M1004_g 0.00468827f $X=3.74 $Y=6.47 $X2=0.475 $Y2=4.585
cc_124 N_VDD_M1004_d N_A_c_208_n 0.00628533f $X=0.55 $Y=3.085 $X2=0.635 $Y2=2.48
cc_125 N_VDD_M1004_b N_A_c_208_n 0.00328912f $X=-0.045 $Y=2.905 $X2=0.635
+ $Y2=2.48
cc_126 N_VDD_c_122_p N_A_c_208_n 0.00264661f $X=0.69 $Y=4.135 $X2=0.635 $Y2=2.48
cc_127 N_VDD_M1004_d A 0.00797576f $X=0.55 $Y=3.085 $X2=0.635 $Y2=3.33
cc_128 N_VDD_c_122_p A 0.00510982f $X=0.69 $Y=4.135 $X2=0.635 $Y2=3.33
cc_129 N_VDD_M1004_b N_A_27_115#_c_311_n 0.014249f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=3.01
cc_130 N_VDD_c_122_p N_A_27_115#_c_311_n 0.00354579f $X=0.69 $Y=4.135 $X2=0.905
+ $Y2=3.01
cc_131 N_VDD_c_131_p N_A_27_115#_c_311_n 0.00606474f $X=1.465 $Y=6.507 $X2=0.905
+ $Y2=3.01
cc_132 N_VDD_c_123_p N_A_27_115#_c_311_n 0.00468827f $X=3.74 $Y=6.47 $X2=0.905
+ $Y2=3.01
cc_133 N_VDD_M1004_b N_A_27_115#_c_315_n 0.0141063f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=3.01
cc_134 N_VDD_c_122_p N_A_27_115#_c_315_n 3.67508e-19 $X=0.69 $Y=4.135 $X2=1.335
+ $Y2=3.01
cc_135 N_VDD_c_131_p N_A_27_115#_c_315_n 0.00610567f $X=1.465 $Y=6.507 $X2=1.335
+ $Y2=3.01
cc_136 N_VDD_c_136_p N_A_27_115#_c_315_n 0.00373985f $X=1.55 $Y=3.455 $X2=1.335
+ $Y2=3.01
cc_137 N_VDD_c_123_p N_A_27_115#_c_315_n 0.00470215f $X=3.74 $Y=6.47 $X2=1.335
+ $Y2=3.01
cc_138 N_VDD_M1004_b N_A_27_115#_c_254_n 0.00647677f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.935
cc_139 N_VDD_c_136_p N_A_27_115#_c_254_n 0.00364479f $X=1.55 $Y=3.455 $X2=1.69
+ $Y2=2.935
cc_140 N_VDD_M1004_b N_A_27_115#_c_255_n 0.0113915f $X=-0.045 $Y=2.905 $X2=1.41
+ $Y2=2.935
cc_141 N_VDD_M1004_b N_A_27_115#_c_323_n 0.0137901f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=3.01
cc_142 N_VDD_c_136_p N_A_27_115#_c_323_n 0.00354579f $X=1.55 $Y=3.455 $X2=1.765
+ $Y2=3.01
cc_143 N_VDD_c_143_p N_A_27_115#_c_323_n 0.00606474f $X=2.325 $Y=6.507 $X2=1.765
+ $Y2=3.01
cc_144 N_VDD_c_123_p N_A_27_115#_c_323_n 0.00468827f $X=3.74 $Y=6.47 $X2=1.765
+ $Y2=3.01
cc_145 N_VDD_M1004_b N_A_27_115#_c_261_n 0.00596183f $X=-0.045 $Y=2.905 $X2=2.12
+ $Y2=2.935
cc_146 N_VDD_M1004_b N_A_27_115#_c_328_n 0.0137901f $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=3.01
cc_147 N_VDD_c_143_p N_A_27_115#_c_328_n 0.00606474f $X=2.325 $Y=6.507 $X2=2.195
+ $Y2=3.01
cc_148 N_VDD_c_148_p N_A_27_115#_c_328_n 0.00354579f $X=2.41 $Y=3.455 $X2=2.195
+ $Y2=3.01
cc_149 N_VDD_c_123_p N_A_27_115#_c_328_n 0.00468827f $X=3.74 $Y=6.47 $X2=2.195
+ $Y2=3.01
cc_150 N_VDD_M1004_b N_A_27_115#_c_268_n 0.00647677f $X=-0.045 $Y=2.905 $X2=2.55
+ $Y2=2.935
cc_151 N_VDD_c_148_p N_A_27_115#_c_268_n 0.00364479f $X=2.41 $Y=3.455 $X2=2.55
+ $Y2=2.935
cc_152 N_VDD_M1004_b N_A_27_115#_c_334_n 0.0137901f $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=3.01
cc_153 N_VDD_c_148_p N_A_27_115#_c_334_n 0.00354579f $X=2.41 $Y=3.455 $X2=2.625
+ $Y2=3.01
cc_154 N_VDD_c_154_p N_A_27_115#_c_334_n 0.00606474f $X=3.185 $Y=6.507 $X2=2.625
+ $Y2=3.01
cc_155 N_VDD_c_123_p N_A_27_115#_c_334_n 0.00468827f $X=3.74 $Y=6.47 $X2=2.625
+ $Y2=3.01
cc_156 N_VDD_M1004_b N_A_27_115#_c_275_n 0.00596183f $X=-0.045 $Y=2.905 $X2=2.98
+ $Y2=2.935
cc_157 N_VDD_M1004_b N_A_27_115#_c_339_n 0.0137901f $X=-0.045 $Y=2.905 $X2=3.055
+ $Y2=3.01
cc_158 N_VDD_c_154_p N_A_27_115#_c_339_n 0.00606474f $X=3.185 $Y=6.507 $X2=3.055
+ $Y2=3.01
cc_159 N_VDD_c_159_p N_A_27_115#_c_339_n 0.00354579f $X=3.27 $Y=3.455 $X2=3.055
+ $Y2=3.01
cc_160 N_VDD_c_123_p N_A_27_115#_c_339_n 0.00468827f $X=3.74 $Y=6.47 $X2=3.055
+ $Y2=3.01
cc_161 N_VDD_M1004_b N_A_27_115#_c_282_n 0.00647677f $X=-0.045 $Y=2.905 $X2=3.41
+ $Y2=2.935
cc_162 N_VDD_c_159_p N_A_27_115#_c_282_n 0.00364479f $X=3.27 $Y=3.455 $X2=3.41
+ $Y2=2.935
cc_163 N_VDD_M1004_b N_A_27_115#_c_345_n 0.0137901f $X=-0.045 $Y=2.905 $X2=3.485
+ $Y2=3.01
cc_164 N_VDD_c_159_p N_A_27_115#_c_345_n 0.00354579f $X=3.27 $Y=3.455 $X2=3.485
+ $Y2=3.01
cc_165 N_VDD_c_165_p N_A_27_115#_c_345_n 0.00606474f $X=4.045 $Y=6.507 $X2=3.485
+ $Y2=3.01
cc_166 N_VDD_c_123_p N_A_27_115#_c_345_n 0.00468827f $X=3.74 $Y=6.47 $X2=3.485
+ $Y2=3.01
cc_167 N_VDD_M1004_b N_A_27_115#_c_288_n 0.0134369f $X=-0.045 $Y=2.905 $X2=3.84
+ $Y2=2.935
cc_168 N_VDD_M1004_b N_A_27_115#_c_350_n 0.0166569f $X=-0.045 $Y=2.905 $X2=3.915
+ $Y2=3.01
cc_169 N_VDD_c_165_p N_A_27_115#_c_350_n 0.00606474f $X=4.045 $Y=6.507 $X2=3.915
+ $Y2=3.01
cc_170 N_VDD_c_170_p N_A_27_115#_c_350_n 0.00713292f $X=4.13 $Y=3.455 $X2=3.915
+ $Y2=3.01
cc_171 N_VDD_c_123_p N_A_27_115#_c_350_n 0.00468827f $X=3.74 $Y=6.47 $X2=3.915
+ $Y2=3.01
cc_172 N_VDD_M1004_b N_A_27_115#_c_294_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.935
cc_173 N_VDD_M1004_b N_A_27_115#_c_296_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.935
cc_174 N_VDD_M1004_b N_A_27_115#_c_298_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=2.935
cc_175 N_VDD_M1004_b N_A_27_115#_c_300_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=3.055 $Y2=2.935
cc_176 N_VDD_M1004_b N_A_27_115#_c_302_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=3.485 $Y2=2.935
cc_177 N_VDD_M1004_b N_A_27_115#_c_306_n 0.00996008f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.455
cc_178 N_VDD_c_121_p N_A_27_115#_c_306_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=3.455
cc_179 N_VDD_c_123_p N_A_27_115#_c_306_n 0.00476261f $X=3.74 $Y=6.47 $X2=0.26
+ $Y2=3.455
cc_180 N_VDD_M1004_b N_Y_c_517_n 0.00290209f $X=-0.045 $Y=2.905 $X2=1.12
+ $Y2=2.96
cc_181 N_VDD_c_131_p N_Y_c_517_n 0.00734006f $X=1.465 $Y=6.507 $X2=1.12 $Y2=2.96
cc_182 N_VDD_c_123_p N_Y_c_517_n 0.00475776f $X=3.74 $Y=6.47 $X2=1.12 $Y2=2.96
cc_183 N_VDD_M1004_b N_Y_c_520_n 0.00337919f $X=-0.045 $Y=2.905 $X2=1.98
+ $Y2=2.96
cc_184 N_VDD_c_143_p N_Y_c_520_n 0.00754406f $X=2.325 $Y=6.507 $X2=1.98 $Y2=2.96
cc_185 N_VDD_c_123_p N_Y_c_520_n 0.00475776f $X=3.74 $Y=6.47 $X2=1.98 $Y2=2.96
cc_186 N_VDD_M1004_b N_Y_c_523_n 0.00337919f $X=-0.045 $Y=2.905 $X2=2.84
+ $Y2=2.96
cc_187 N_VDD_c_154_p N_Y_c_523_n 0.00746708f $X=3.185 $Y=6.507 $X2=2.84 $Y2=2.96
cc_188 N_VDD_c_123_p N_Y_c_523_n 0.00475776f $X=3.74 $Y=6.47 $X2=2.84 $Y2=2.96
cc_189 N_VDD_M1004_b N_Y_c_526_n 0.00337919f $X=-0.045 $Y=2.905 $X2=3.7 $Y2=2.96
cc_190 N_VDD_c_165_p N_Y_c_526_n 0.00734006f $X=4.045 $Y=6.507 $X2=3.7 $Y2=2.96
cc_191 N_VDD_c_123_p N_Y_c_526_n 0.00475776f $X=3.74 $Y=6.47 $X2=3.7 $Y2=2.96
cc_192 N_VDD_M1004_b N_Y_c_495_n 0.00409378f $X=-0.045 $Y=2.905 $X2=1.12
+ $Y2=2.845
cc_193 N_VDD_M1004_b N_Y_c_530_n 0.00520877f $X=-0.045 $Y=2.905 $X2=1.835
+ $Y2=2.96
cc_194 N_VDD_c_136_p N_Y_c_530_n 0.0090257f $X=1.55 $Y=3.455 $X2=1.835 $Y2=2.96
cc_195 N_VDD_M1004_b N_Y_c_532_n 0.00520877f $X=-0.045 $Y=2.905 $X2=2.695
+ $Y2=2.96
cc_196 N_VDD_c_148_p N_Y_c_532_n 0.0090257f $X=2.41 $Y=3.455 $X2=2.695 $Y2=2.96
cc_197 N_VDD_M1004_b N_Y_c_505_n 0.00409378f $X=-0.045 $Y=2.905 $X2=2.125
+ $Y2=2.96
cc_198 N_VDD_M1004_b N_Y_c_535_n 0.00520877f $X=-0.045 $Y=2.905 $X2=3.555
+ $Y2=2.96
cc_199 N_VDD_c_159_p N_Y_c_535_n 0.0090257f $X=3.27 $Y=3.455 $X2=3.555 $Y2=2.96
cc_200 N_VDD_M1004_b N_Y_c_512_n 0.00409378f $X=-0.045 $Y=2.905 $X2=2.985
+ $Y2=2.96
cc_201 N_VDD_M1004_b N_Y_c_516_n 0.00409378f $X=-0.045 $Y=2.905 $X2=3.7
+ $Y2=2.845
cc_202 A N_A_27_115#_M1004_s 0.00414531f $X=0.635 $Y=3.33 $X2=0.135 $Y2=3.085
cc_203 N_A_M1006_g N_A_27_115#_M1001_g 0.0387262f $X=0.475 $Y=1.075 $X2=0.905
+ $Y2=1.075
cc_204 A N_A_27_115#_c_311_n 0.00419145f $X=0.635 $Y=3.33 $X2=0.905 $Y2=3.01
cc_205 N_A_M1006_g N_A_27_115#_c_246_n 0.00260138f $X=0.475 $Y=1.075 $X2=1.18
+ $Y2=2.86
cc_206 N_A_M1004_g N_A_27_115#_c_246_n 0.00209773f $X=0.475 $Y=4.585 $X2=1.18
+ $Y2=2.86
cc_207 N_A_c_207_n N_A_27_115#_c_246_n 0.0139096f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_208 N_A_c_208_n N_A_27_115#_c_246_n 0.00361737f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_209 N_A_M1004_g N_A_27_115#_c_255_n 0.0499373f $X=0.475 $Y=4.585 $X2=1.41
+ $Y2=2.935
cc_210 N_A_c_208_n N_A_27_115#_c_255_n 0.00477416f $X=0.635 $Y=2.48 $X2=1.41
+ $Y2=2.935
cc_211 N_A_M1006_g N_A_27_115#_c_303_n 0.0148408f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_212 N_A_M1006_g N_A_27_115#_c_306_n 0.0337582f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=3.455
cc_213 N_A_c_208_n N_A_27_115#_c_306_n 0.0548951f $X=0.635 $Y=2.48 $X2=0.26
+ $Y2=3.455
cc_214 A N_A_27_115#_c_306_n 0.0155137f $X=0.635 $Y=3.33 $X2=0.26 $Y2=3.455
cc_215 N_A_M1006_g N_A_27_115#_c_307_n 0.0207696f $X=0.475 $Y=1.075 $X2=0.88
+ $Y2=1.935
cc_216 N_A_c_207_n N_A_27_115#_c_307_n 0.00273049f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_217 N_A_c_208_n N_A_27_115#_c_307_n 0.00886797f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_218 N_A_M1006_g N_A_27_115#_c_310_n 6.59135e-19 $X=0.475 $Y=1.075 $X2=0.965
+ $Y2=1.935
cc_219 N_A_c_208_n N_Y_c_517_n 0.0135622f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_220 A N_Y_c_517_n 0.00731851f $X=0.635 $Y=3.33 $X2=1.12 $Y2=2.96
cc_221 N_A_M1006_g N_Y_c_492_n 8.23842e-19 $X=0.475 $Y=1.075 $X2=1.12 $Y2=1.595
cc_222 N_A_c_208_n N_Y_c_495_n 0.00677552f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.845
cc_223 N_A_M1006_g Y 0.00310306f $X=0.475 $Y=1.075 $X2=1.055 $Y2=2.27
cc_224 N_A_c_207_n Y 0.00441844f $X=0.635 $Y=2.48 $X2=1.055 $Y2=2.27
cc_225 N_A_c_208_n Y 0.0200396f $X=0.635 $Y=2.48 $X2=1.055 $Y2=2.27
cc_226 N_A_27_115#_M1001_g N_Y_c_474_n 0.00231637f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_227 N_A_27_115#_M1003_g N_Y_c_474_n 0.00231637f $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_228 N_A_27_115#_c_253_n N_Y_c_474_n 0.0030245f $X=1.41 $Y=1.845 $X2=1.12
+ $Y2=0.825
cc_229 N_A_27_115#_c_310_n N_Y_c_474_n 7.32051e-19 $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_230 N_A_27_115#_c_311_n N_Y_c_517_n 0.00155107f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_231 N_A_27_115#_c_315_n N_Y_c_517_n 0.00250481f $X=1.335 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_232 N_A_27_115#_c_255_n N_Y_c_517_n 0.0126676f $X=1.41 $Y=2.935 $X2=1.12
+ $Y2=2.96
cc_233 N_A_27_115#_M1007_g N_Y_c_478_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.98
+ $Y2=0.825
cc_234 N_A_27_115#_c_260_n N_Y_c_478_n 0.00280419f $X=2.12 $Y=1.845 $X2=1.98
+ $Y2=0.825
cc_235 N_A_27_115#_M1010_g N_Y_c_478_n 0.00231637f $X=2.195 $Y=1.075 $X2=1.98
+ $Y2=0.825
cc_236 N_A_27_115#_c_323_n N_Y_c_520_n 0.00250481f $X=1.765 $Y=3.01 $X2=1.98
+ $Y2=2.96
cc_237 N_A_27_115#_c_261_n N_Y_c_520_n 0.0138847f $X=2.12 $Y=2.935 $X2=1.98
+ $Y2=2.96
cc_238 N_A_27_115#_c_328_n N_Y_c_520_n 0.00250481f $X=2.195 $Y=3.01 $X2=1.98
+ $Y2=2.96
cc_239 N_A_27_115#_M1011_g N_Y_c_483_n 0.00231637f $X=2.625 $Y=1.075 $X2=2.84
+ $Y2=0.825
cc_240 N_A_27_115#_c_274_n N_Y_c_483_n 0.00280419f $X=2.98 $Y=1.845 $X2=2.84
+ $Y2=0.825
cc_241 N_A_27_115#_M1014_g N_Y_c_483_n 0.00231637f $X=3.055 $Y=1.075 $X2=2.84
+ $Y2=0.825
cc_242 N_A_27_115#_c_334_n N_Y_c_523_n 0.00250481f $X=2.625 $Y=3.01 $X2=2.84
+ $Y2=2.96
cc_243 N_A_27_115#_c_275_n N_Y_c_523_n 0.0138847f $X=2.98 $Y=2.935 $X2=2.84
+ $Y2=2.96
cc_244 N_A_27_115#_c_339_n N_Y_c_523_n 0.00250481f $X=3.055 $Y=3.01 $X2=2.84
+ $Y2=2.96
cc_245 N_A_27_115#_M1015_g N_Y_c_488_n 0.00231637f $X=3.485 $Y=1.075 $X2=3.7
+ $Y2=0.825
cc_246 N_A_27_115#_c_287_n N_Y_c_488_n 0.00280419f $X=3.84 $Y=1.845 $X2=3.7
+ $Y2=0.825
cc_247 N_A_27_115#_M1017_g N_Y_c_488_n 0.00231637f $X=3.915 $Y=1.075 $X2=3.7
+ $Y2=0.825
cc_248 N_A_27_115#_c_345_n N_Y_c_526_n 0.00250481f $X=3.485 $Y=3.01 $X2=3.7
+ $Y2=2.96
cc_249 N_A_27_115#_c_288_n N_Y_c_526_n 0.013404f $X=3.84 $Y=2.935 $X2=3.7
+ $Y2=2.96
cc_250 N_A_27_115#_c_350_n N_Y_c_526_n 0.00250481f $X=3.915 $Y=3.01 $X2=3.7
+ $Y2=2.96
cc_251 N_A_27_115#_M1001_g N_Y_c_492_n 0.00541983f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=1.595
cc_252 N_A_27_115#_M1003_g N_Y_c_492_n 0.00262362f $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=1.595
cc_253 N_A_27_115#_c_310_n N_Y_c_492_n 0.00278861f $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=1.595
cc_254 N_A_27_115#_c_311_n N_Y_c_495_n 0.00120715f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.845
cc_255 N_A_27_115#_c_246_n N_Y_c_495_n 0.00215118f $X=1.18 $Y=2.86 $X2=1.12
+ $Y2=2.845
cc_256 N_A_27_115#_c_315_n N_Y_c_495_n 0.00113627f $X=1.335 $Y=3.01 $X2=1.12
+ $Y2=2.845
cc_257 N_A_27_115#_c_255_n N_Y_c_495_n 0.00372325f $X=1.41 $Y=2.935 $X2=1.12
+ $Y2=2.845
cc_258 N_A_27_115#_M1001_g Y 0.00251111f $X=0.905 $Y=1.075 $X2=1.055 $Y2=2.27
cc_259 N_A_27_115#_c_246_n Y 0.0314621f $X=1.18 $Y=2.86 $X2=1.055 $Y2=2.27
cc_260 N_A_27_115#_M1003_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.055 $Y2=2.27
cc_261 N_A_27_115#_c_253_n Y 0.0166018f $X=1.41 $Y=1.845 $X2=1.055 $Y2=2.27
cc_262 N_A_27_115#_c_307_n Y 8.73078e-19 $X=0.88 $Y=1.935 $X2=1.055 $Y2=2.27
cc_263 N_A_27_115#_c_310_n Y 0.0121742f $X=0.965 $Y=1.935 $X2=1.055 $Y2=2.27
cc_264 N_A_27_115#_M1003_g N_Y_c_497_n 0.0133661f $X=1.335 $Y=1.075 $X2=1.835
+ $Y2=1.48
cc_265 N_A_27_115#_c_251_n N_Y_c_497_n 0.00213861f $X=1.69 $Y=1.845 $X2=1.835
+ $Y2=1.48
cc_266 N_A_27_115#_M1007_g N_Y_c_497_n 0.0130095f $X=1.765 $Y=1.075 $X2=1.835
+ $Y2=1.48
cc_267 N_A_27_115#_c_315_n N_Y_c_530_n 0.00639369f $X=1.335 $Y=3.01 $X2=1.835
+ $Y2=2.96
cc_268 N_A_27_115#_c_254_n N_Y_c_530_n 0.0125005f $X=1.69 $Y=2.935 $X2=1.835
+ $Y2=2.96
cc_269 N_A_27_115#_c_255_n N_Y_c_530_n 0.00627763f $X=1.41 $Y=2.935 $X2=1.835
+ $Y2=2.96
cc_270 N_A_27_115#_c_323_n N_Y_c_530_n 0.00639369f $X=1.765 $Y=3.01 $X2=1.835
+ $Y2=2.96
cc_271 N_A_27_115#_c_294_n N_Y_c_530_n 0.00580646f $X=1.765 $Y=2.935 $X2=1.835
+ $Y2=2.96
cc_272 N_A_27_115#_c_253_n N_Y_c_499_n 0.013329f $X=1.41 $Y=1.845 $X2=1.98
+ $Y2=2.845
cc_273 N_A_27_115#_M1007_g N_Y_c_499_n 0.00251111f $X=1.765 $Y=1.075 $X2=1.98
+ $Y2=2.845
cc_274 N_A_27_115#_c_260_n N_Y_c_499_n 0.0178059f $X=2.12 $Y=1.845 $X2=1.98
+ $Y2=2.845
cc_275 N_A_27_115#_M1010_g N_Y_c_499_n 0.00251111f $X=2.195 $Y=1.075 $X2=1.98
+ $Y2=2.845
cc_276 N_A_27_115#_c_273_n N_Y_c_499_n 0.0137936f $X=2.625 $Y=2.86 $X2=1.98
+ $Y2=2.845
cc_277 N_A_27_115#_M1010_g N_Y_c_500_n 0.0130095f $X=2.195 $Y=1.075 $X2=2.695
+ $Y2=1.48
cc_278 N_A_27_115#_c_266_n N_Y_c_500_n 0.00213861f $X=2.55 $Y=1.845 $X2=2.695
+ $Y2=1.48
cc_279 N_A_27_115#_M1011_g N_Y_c_500_n 0.0136594f $X=2.625 $Y=1.075 $X2=2.695
+ $Y2=1.48
cc_280 N_A_27_115#_M1007_g N_Y_c_502_n 0.00259902f $X=1.765 $Y=1.075 $X2=2.125
+ $Y2=1.48
cc_281 N_A_27_115#_M1010_g N_Y_c_502_n 0.00259902f $X=2.195 $Y=1.075 $X2=2.125
+ $Y2=1.48
cc_282 N_A_27_115#_c_328_n N_Y_c_532_n 0.00639369f $X=2.195 $Y=3.01 $X2=2.695
+ $Y2=2.96
cc_283 N_A_27_115#_c_268_n N_Y_c_532_n 0.0130313f $X=2.55 $Y=2.935 $X2=2.695
+ $Y2=2.96
cc_284 N_A_27_115#_c_334_n N_Y_c_532_n 0.00639369f $X=2.625 $Y=3.01 $X2=2.695
+ $Y2=2.96
cc_285 N_A_27_115#_c_296_n N_Y_c_532_n 0.00580646f $X=2.195 $Y=2.935 $X2=2.695
+ $Y2=2.96
cc_286 N_A_27_115#_c_298_n N_Y_c_532_n 0.00666531f $X=2.625 $Y=2.935 $X2=2.695
+ $Y2=2.96
cc_287 N_A_27_115#_c_323_n N_Y_c_505_n 0.00113627f $X=1.765 $Y=3.01 $X2=2.125
+ $Y2=2.96
cc_288 N_A_27_115#_c_261_n N_Y_c_505_n 0.00364679f $X=2.12 $Y=2.935 $X2=2.125
+ $Y2=2.96
cc_289 N_A_27_115#_c_328_n N_Y_c_505_n 0.00113627f $X=2.195 $Y=3.01 $X2=2.125
+ $Y2=2.96
cc_290 N_A_27_115#_c_294_n N_Y_c_505_n 6.99501e-19 $X=1.765 $Y=2.935 $X2=2.125
+ $Y2=2.96
cc_291 N_A_27_115#_c_296_n N_Y_c_505_n 6.99501e-19 $X=2.195 $Y=2.935 $X2=2.125
+ $Y2=2.96
cc_292 N_A_27_115#_M1011_g N_Y_c_506_n 0.00251111f $X=2.625 $Y=1.075 $X2=2.84
+ $Y2=2.845
cc_293 N_A_27_115#_c_273_n N_Y_c_506_n 0.017762f $X=2.625 $Y=2.86 $X2=2.84
+ $Y2=2.845
cc_294 N_A_27_115#_c_274_n N_Y_c_506_n 0.0178059f $X=2.98 $Y=1.845 $X2=2.84
+ $Y2=2.845
cc_295 N_A_27_115#_M1014_g N_Y_c_506_n 0.00251111f $X=3.055 $Y=1.075 $X2=2.84
+ $Y2=2.845
cc_296 N_A_27_115#_M1014_g N_Y_c_507_n 0.0130095f $X=3.055 $Y=1.075 $X2=3.555
+ $Y2=1.48
cc_297 N_A_27_115#_c_280_n N_Y_c_507_n 0.00213861f $X=3.41 $Y=1.845 $X2=3.555
+ $Y2=1.48
cc_298 N_A_27_115#_M1015_g N_Y_c_507_n 0.0130095f $X=3.485 $Y=1.075 $X2=3.555
+ $Y2=1.48
cc_299 N_A_27_115#_M1011_g N_Y_c_509_n 0.00262362f $X=2.625 $Y=1.075 $X2=2.985
+ $Y2=1.48
cc_300 N_A_27_115#_M1014_g N_Y_c_509_n 0.00259902f $X=3.055 $Y=1.075 $X2=2.985
+ $Y2=1.48
cc_301 N_A_27_115#_c_339_n N_Y_c_535_n 0.00639369f $X=3.055 $Y=3.01 $X2=3.555
+ $Y2=2.96
cc_302 N_A_27_115#_c_282_n N_Y_c_535_n 0.0125005f $X=3.41 $Y=2.935 $X2=3.555
+ $Y2=2.96
cc_303 N_A_27_115#_c_345_n N_Y_c_535_n 0.00639369f $X=3.485 $Y=3.01 $X2=3.555
+ $Y2=2.96
cc_304 N_A_27_115#_c_300_n N_Y_c_535_n 0.00580646f $X=3.055 $Y=2.935 $X2=3.555
+ $Y2=2.96
cc_305 N_A_27_115#_c_302_n N_Y_c_535_n 0.00580646f $X=3.485 $Y=2.935 $X2=3.555
+ $Y2=2.96
cc_306 N_A_27_115#_c_273_n N_Y_c_512_n 8.30534e-19 $X=2.625 $Y=2.86 $X2=2.985
+ $Y2=2.96
cc_307 N_A_27_115#_c_334_n N_Y_c_512_n 0.00113627f $X=2.625 $Y=3.01 $X2=2.985
+ $Y2=2.96
cc_308 N_A_27_115#_c_275_n N_Y_c_512_n 0.00364679f $X=2.98 $Y=2.935 $X2=2.985
+ $Y2=2.96
cc_309 N_A_27_115#_c_339_n N_Y_c_512_n 0.00113627f $X=3.055 $Y=3.01 $X2=2.985
+ $Y2=2.96
cc_310 N_A_27_115#_c_298_n N_Y_c_512_n 6.59375e-19 $X=2.625 $Y=2.935 $X2=2.985
+ $Y2=2.96
cc_311 N_A_27_115#_c_300_n N_Y_c_512_n 6.99501e-19 $X=3.055 $Y=2.935 $X2=2.985
+ $Y2=2.96
cc_312 N_A_27_115#_M1015_g N_Y_c_513_n 0.00259902f $X=3.485 $Y=1.075 $X2=3.7
+ $Y2=1.595
cc_313 N_A_27_115#_M1017_g N_Y_c_513_n 0.00939545f $X=3.915 $Y=1.075 $X2=3.7
+ $Y2=1.595
cc_314 N_A_27_115#_M1015_g N_Y_c_516_n 0.00251111f $X=3.485 $Y=1.075 $X2=3.7
+ $Y2=2.845
cc_315 N_A_27_115#_c_345_n N_Y_c_516_n 0.00113627f $X=3.485 $Y=3.01 $X2=3.7
+ $Y2=2.845
cc_316 N_A_27_115#_c_287_n N_Y_c_516_n 0.0170354f $X=3.84 $Y=1.845 $X2=3.7
+ $Y2=2.845
cc_317 N_A_27_115#_c_288_n N_Y_c_516_n 0.00966211f $X=3.84 $Y=2.935 $X2=3.7
+ $Y2=2.845
cc_318 N_A_27_115#_M1017_g N_Y_c_516_n 0.00251111f $X=3.915 $Y=1.075 $X2=3.7
+ $Y2=2.845
cc_319 N_A_27_115#_c_350_n N_Y_c_516_n 0.0031083f $X=3.915 $Y=3.01 $X2=3.7
+ $Y2=2.845
cc_320 N_A_27_115#_c_302_n N_Y_c_516_n 6.99501e-19 $X=3.485 $Y=2.935 $X2=3.7
+ $Y2=2.845
