* File: sky130_osu_sc_12T_ls__tielo.spice
* Created: Fri Nov 12 15:40:41 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__tielo.pex.spice"
.subckt sky130_osu_sc_12T_ls__tielo  GND VDD Y
* 
* Y	Y
* VDD	VDD
* GND	GND
MM1001 N_Y_M1001_d N_A_80_89#_M1001_g N_GND_M1001_s N_GND_M1001_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.1378 PD=1.57 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_A_80_89#_M1000_d N_A_80_89#_M1000_g N_VDD_M1000_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=2.1424 P=6.2
pX3_noxref noxref_5 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__tielo.pxi.spice"
*
.ends
*
*
