* File: sky130_osu_sc_15T_ms__mux2_1.pex.spice
* Created: Fri Nov 12 14:44:53 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%GND 1 29 33 54 56
r35 54 56 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r36 31 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r37 29 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r38 29 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r39 29 31 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r40 29 35 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r41 29 35 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r42 1 33 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%VDD 1 9 13 19 23
r30 23 26 0.00227273 $w=2.75e-06 $l=5e-08 $layer=MET1_cond $X=1.375 $Y=5.31
+ $X2=1.375 $Y2=5.36
r31 19 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.38 $Y=5.36
+ $X2=2.38 $Y2=5.36
r32 17 19 76.8925 $w=3.03e-07 $l=2.035e-06 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=2.38 $Y2=5.397
r33 13 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r34 11 17 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.345 $Y2=5.397
r35 11 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r36 9 19 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r37 1 16 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r38 1 13 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%A_110_115# 1 3 9 11 15 19 24 28 31 34 37
+ 44 49
c69 9 0 3.63536e-20 $X=1.35 $Y=1.53
r70 46 49 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=2.43
+ $X2=0.925 $Y2=2.43
r71 41 44 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.925 $Y2=1.59
r72 37 39 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r73 35 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.595
+ $X2=0.69 $Y2=2.43
r74 35 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.69 $Y=2.595
+ $X2=0.69 $Y2=3.205
r75 34 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.265
+ $X2=0.69 $Y2=2.43
r76 33 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.755
+ $X2=0.69 $Y2=1.59
r77 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.69 $Y=1.755
+ $X2=0.69 $Y2=2.265
r78 29 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.425
+ $X2=0.69 $Y2=1.59
r79 29 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.69 $Y=1.425
+ $X2=0.69 $Y2=0.865
r80 26 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.43 $X2=0.925 $Y2=2.43
r81 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.43
+ $X2=1.09 $Y2=2.43
r82 22 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.59 $X2=0.925 $Y2=1.59
r83 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.59
+ $X2=1.09 $Y2=1.59
r84 17 19 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=1.855 $Y=2.445
+ $X2=1.855 $Y2=3.825
r85 13 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.425 $Y=1.455
+ $X2=1.425 $Y2=0.945
r86 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.37
+ $X2=1.855 $Y2=2.445
r87 11 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.78 $Y=2.37
+ $X2=1.09 $Y2=2.37
r88 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=1.53
+ $X2=1.425 $Y2=1.455
r89 9 24 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.35 $Y=1.53 $X2=1.09
+ $Y2=1.53
r90 3 39 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r91 3 37 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r92 1 31 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%S0 3 8 9 11 12 13 15 18 24 26 32
c65 8 0 1.8854e-20 $X=0.475 $Y=3.825
r66 29 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.07
+ $X2=0.27 $Y2=3.07
r67 26 29 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.27 $Y=2.045
+ $X2=0.27 $Y2=3.07
r68 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.045
+ $X2=0.55 $Y2=2.045
r69 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.045 $X2=0.27 $Y2=2.045
r70 21 23 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.045
+ $X2=0.475 $Y2=2.045
r71 16 18 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=1.855 $Y=1.935
+ $X2=1.855 $Y2=0.945
r72 13 15 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.425 $Y=4.9
+ $X2=1.425 $Y2=3.825
r73 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=4.975
+ $X2=1.425 $Y2=4.9
r74 11 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.35 $Y=4.975 $X2=0.55
+ $Y2=4.975
r75 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.01
+ $X2=1.855 $Y2=1.935
r76 9 24 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.78 $Y=2.01
+ $X2=0.55 $Y2=2.01
r77 6 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=4.9
+ $X2=0.55 $Y2=4.975
r78 6 8 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.475 $Y=4.9
+ $X2=0.475 $Y2=3.825
r79 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.21
+ $X2=0.475 $Y2=2.045
r80 5 8 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=0.475 $Y=2.21
+ $X2=0.475 $Y2=3.825
r81 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.88
+ $X2=0.475 $Y2=2.045
r82 1 3 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.475 $Y=1.88
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%A0 1 3 11 15 22 24 26 28
c40 28 0 1.8854e-20 $X=1.265 $Y=2.7
r41 25 26 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=2.855
+ $X2=1.237 $Y2=3.025
r42 23 24 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=1.075
+ $X2=1.237 $Y2=1.245
r43 22 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.265 $Y=2.7
+ $X2=1.265 $Y2=2.7
r44 22 25 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.265 $Y=2.7
+ $X2=1.265 $Y2=2.855
r45 22 24 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=1.265 $Y=2.7
+ $X2=1.265 $Y2=1.245
r46 15 17 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.21 $Y=3.205
+ $X2=1.21 $Y2=4.565
r47 15 26 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.21 $Y=3.205
+ $X2=1.21 $Y2=3.025
r48 11 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.21 $Y=0.865
+ $X2=1.21 $Y2=1.075
r49 3 17 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.825 $X2=1.21 $Y2=4.565
r50 3 15 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.825 $X2=1.21 $Y2=3.205
r51 1 11 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%Y 1 3 10 16 24 26 29
c36 29 0 3.63536e-20 $X=1.64 $Y=1.96
r37 24 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=1.845
+ $X2=1.64 $Y2=1.96
r38 23 26 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=1.335
+ $X2=1.64 $Y2=1.22
r39 23 24 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=1.64 $Y=1.335
+ $X2=1.64 $Y2=1.845
r40 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.64 $Y=3.205
+ $X2=1.64 $Y2=4.565
r41 16 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.96
+ $X2=1.64 $Y2=1.96
r42 16 19 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=1.64 $Y=1.96
+ $X2=1.64 $Y2=3.205
r43 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.22
+ $X2=1.64 $Y2=1.22
r44 10 13 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.64 $Y=0.865
+ $X2=1.64 $Y2=1.22
r45 3 21 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.825 $X2=1.64 $Y2=4.565
r46 3 19 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.825 $X2=1.64 $Y2=3.205
r47 1 10 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__MUX2_1%A1 1 3 10 20
r17 15 17 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.07 $Y=3.205
+ $X2=2.07 $Y2=4.565
r18 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.33
+ $X2=2.07 $Y2=2.33
r19 13 15 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.07 $Y=2.33
+ $X2=2.07 $Y2=3.205
r20 10 13 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=2.07 $Y=0.865
+ $X2=2.07 $Y2=2.33
r21 3 17 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=2.825 $X2=2.07 $Y2=4.565
r22 3 15 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=2.825 $X2=2.07 $Y2=3.205
r23 1 10 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.865
.ends

