* File: sky130_osu_sc_15T_ls__xor2_l.pxi.spice
* Created: Fri Nov 12 15:00:53 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%GND N_GND_M1002_d N_GND_M1008_d N_GND_M1002_b
+ N_GND_c_9_p N_GND_c_2_p N_GND_c_3_p N_GND_c_39_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_15T_LS__XOR2_L%GND
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%VDD N_VDD_M1001_d N_VDD_M1009_d N_VDD_M1001_b
+ N_VDD_c_72_p N_VDD_c_77_p N_VDD_c_68_p N_VDD_c_99_p N_VDD_c_95_p VDD
+ N_VDD_c_69_p PM_SKY130_OSU_SC_15T_LS__XOR2_L%VDD
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_M1010_g
+ N_A_27_115#_c_116_n N_A_27_115#_c_118_n N_A_27_115#_c_119_n
+ N_A_27_115#_c_122_n N_A_27_115#_c_123_n N_A_27_115#_c_124_n
+ N_A_27_115#_c_125_n PM_SKY130_OSU_SC_15T_LS__XOR2_L%A_27_115#
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%A N_A_c_188_n N_A_M1002_g N_A_c_206_n
+ N_A_M1001_g N_A_c_189_n N_A_M1005_g N_A_M1007_g N_A_c_193_n N_A_c_194_n
+ N_A_c_195_n N_A_c_199_n N_A_c_200_n N_A_c_201_n N_A_c_213_n N_A_c_202_n
+ N_A_c_217_n N_A_c_203_n N_A_c_204_n N_A_c_220_n N_A_c_205_n N_A_c_246_n
+ N_A_c_248_n A N_A_c_249_n PM_SKY130_OSU_SC_15T_LS__XOR2_L%A
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%A_238_89# N_A_238_89#_M1003_d
+ N_A_238_89#_M1004_d N_A_238_89#_M1011_g N_A_238_89#_M1006_g
+ N_A_238_89#_c_311_n N_A_238_89#_c_312_n N_A_238_89#_c_315_n
+ N_A_238_89#_c_317_n N_A_238_89#_c_319_n N_A_238_89#_c_320_n
+ PM_SKY130_OSU_SC_15T_LS__XOR2_L%A_238_89#
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%B N_B_c_374_n N_B_M1008_g N_B_c_389_n
+ N_B_M1009_g N_B_c_378_n N_B_c_380_n N_B_c_381_n N_B_M1003_g N_B_c_384_n
+ N_B_c_393_n N_B_M1004_g N_B_c_385_n N_B_c_386_n N_B_c_387_n B
+ PM_SKY130_OSU_SC_15T_LS__XOR2_L%B
x_PM_SKY130_OSU_SC_15T_LS__XOR2_L%Y N_Y_M1011_d N_Y_M1006_d N_Y_c_432_n
+ N_Y_c_462_n N_Y_c_433_n N_Y_c_441_n N_Y_c_448_n Y N_Y_c_437_n N_Y_c_438_n
+ PM_SKY130_OSU_SC_15T_LS__XOR2_L%Y
cc_1 N_GND_M1002_b N_A_27_115#_M1000_g 0.0358816f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.945
cc_2 N_GND_c_2_p N_A_27_115#_M1000_g 0.00388248f $X=0.69 $Y=0.865 $X2=0.905
+ $Y2=0.945
cc_3 N_GND_c_3_p N_A_27_115#_M1000_g 0.00606474f $X=2.355 $Y=0.152 $X2=0.905
+ $Y2=0.945
cc_4 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.905
+ $Y2=0.945
cc_5 N_GND_M1002_b N_A_27_115#_c_116_n 0.0277843f $X=-0.045 $Y=0 $X2=0.845
+ $Y2=1.965
cc_6 N_GND_c_2_p N_A_27_115#_c_116_n 0.00172615f $X=0.69 $Y=0.865 $X2=0.845
+ $Y2=1.965
cc_7 N_GND_M1002_b N_A_27_115#_c_118_n 0.0287684f $X=-0.045 $Y=0 $X2=1.805
+ $Y2=2.505
cc_8 N_GND_M1002_b N_A_27_115#_c_119_n 0.028416f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_9 N_GND_c_9_p N_A_27_115#_c_119_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_10 N_GND_c_4_p N_A_27_115#_c_119_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_11 N_GND_M1002_b N_A_27_115#_c_122_n 0.0279827f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.205
cc_12 N_GND_M1002_b N_A_27_115#_c_123_n 0.0351362f $X=-0.045 $Y=0 $X2=1.72
+ $Y2=1.965
cc_13 N_GND_M1002_b N_A_27_115#_c_124_n 0.00402941f $X=-0.045 $Y=0 $X2=1.805
+ $Y2=2.505
cc_14 N_GND_M1002_b N_A_27_115#_c_125_n 0.00692367f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.965
cc_15 N_GND_M1002_b N_A_c_188_n 0.0619806f $X=-0.045 $Y=0 $X2=0.425 $Y2=2.6
cc_16 N_GND_M1002_b N_A_c_189_n 0.00178356f $X=-0.045 $Y=0 $X2=0.71 $Y2=2.675
cc_17 N_GND_M1002_b N_A_M1007_g 0.0361289f $X=-0.045 $Y=0 $X2=1.865 $Y2=0.945
cc_18 N_GND_c_3_p N_A_M1007_g 0.00606474f $X=2.355 $Y=0.152 $X2=1.865 $Y2=0.945
cc_19 N_GND_c_4_p N_A_M1007_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.865 $Y2=0.945
cc_20 N_GND_M1002_b N_A_c_193_n 0.0125853f $X=-0.045 $Y=0 $X2=2.1 $Y2=1.825
cc_21 N_GND_M1002_b N_A_c_194_n 0.00928792f $X=-0.045 $Y=0 $X2=1.94 $Y2=1.825
cc_22 N_GND_M1002_b N_A_c_195_n 0.0186719f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.39
cc_23 N_GND_c_9_p N_A_c_195_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.45 $Y2=1.39
cc_24 N_GND_c_2_p N_A_c_195_n 0.00388248f $X=0.69 $Y=0.865 $X2=0.45 $Y2=1.39
cc_25 N_GND_c_4_p N_A_c_195_n 0.00468827f $X=2.38 $Y=0.19 $X2=0.45 $Y2=1.39
cc_26 N_GND_M1002_b N_A_c_199_n 0.012055f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.515
cc_27 N_GND_M1002_b N_A_c_200_n 0.00205699f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.675
cc_28 N_GND_M1002_b N_A_c_201_n 0.0203167f $X=-0.045 $Y=0 $X2=0.845 $Y2=2.505
cc_29 N_GND_M1002_b N_A_c_202_n 0.0338763f $X=-0.045 $Y=0 $X2=2.235 $Y2=1.825
cc_30 N_GND_M1002_b N_A_c_203_n 0.00930883f $X=-0.045 $Y=0 $X2=2.145 $Y2=3.07
cc_31 N_GND_M1002_b N_A_c_204_n 0.00457153f $X=-0.045 $Y=0 $X2=0.845 $Y2=2.505
cc_32 N_GND_M1002_b N_A_c_205_n 0.00312742f $X=-0.045 $Y=0 $X2=2.235 $Y2=1.96
cc_33 N_GND_M1002_b N_A_238_89#_M1006_g 0.053375f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=3.825
cc_34 N_GND_M1002_b N_A_238_89#_c_311_n 0.0270758f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=1.59
cc_35 N_GND_M1002_b N_A_238_89#_c_312_n 0.0169421f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=1.425
cc_36 N_GND_c_3_p N_A_238_89#_c_312_n 0.00606474f $X=2.355 $Y=0.152 $X2=1.325
+ $Y2=1.425
cc_37 N_GND_c_4_p N_A_238_89#_c_312_n 0.00468827f $X=2.38 $Y=0.19 $X2=1.325
+ $Y2=1.425
cc_38 N_GND_M1002_b N_A_238_89#_c_315_n 0.026678f $X=-0.045 $Y=0 $X2=2.785
+ $Y2=1.59
cc_39 N_GND_c_39_p N_A_238_89#_c_315_n 0.00756829f $X=2.44 $Y=0.865 $X2=2.785
+ $Y2=1.59
cc_40 N_GND_M1002_b N_A_238_89#_c_317_n 0.0176967f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=0.865
cc_41 N_GND_c_4_p N_A_238_89#_c_317_n 0.00476261f $X=2.38 $Y=0.19 $X2=2.87
+ $Y2=0.865
cc_42 N_GND_M1002_b N_A_238_89#_c_319_n 0.045758f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=3.205
cc_43 N_GND_M1002_b N_A_238_89#_c_320_n 0.00720662f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=1.59
cc_44 N_GND_M1002_b N_B_c_374_n 0.0139689f $X=-0.045 $Y=0 $X2=2.225 $Y2=1.39
cc_45 N_GND_c_3_p N_B_c_374_n 0.00606474f $X=2.355 $Y=0.152 $X2=2.225 $Y2=1.39
cc_46 N_GND_c_39_p N_B_c_374_n 0.00388248f $X=2.44 $Y=0.865 $X2=2.225 $Y2=1.39
cc_47 N_GND_c_4_p N_B_c_374_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.225 $Y2=1.39
cc_48 N_GND_M1002_b N_B_c_378_n 0.0134223f $X=-0.045 $Y=0 $X2=2.58 $Y2=1.465
cc_49 N_GND_c_39_p N_B_c_378_n 0.00209358f $X=2.44 $Y=0.865 $X2=2.58 $Y2=1.465
cc_50 N_GND_M1002_b N_B_c_380_n 0.00622799f $X=-0.045 $Y=0 $X2=2.3 $Y2=1.465
cc_51 N_GND_M1002_b N_B_c_381_n 0.0243938f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.39
cc_52 N_GND_c_39_p N_B_c_381_n 0.00388248f $X=2.44 $Y=0.865 $X2=2.655 $Y2=1.39
cc_53 N_GND_c_4_p N_B_c_381_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.655 $Y2=1.39
cc_54 N_GND_M1002_b N_B_c_384_n 0.0434452f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.34
cc_55 N_GND_M1002_b N_B_c_385_n 0.0377483f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.545
cc_56 N_GND_M1002_b N_B_c_386_n 0.0061678f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.465
cc_57 N_GND_M1002_b N_B_c_387_n 0.00229251f $X=-0.045 $Y=0 $X2=2.53 $Y2=2.505
cc_58 N_GND_M1002_b B 2.21435e-19 $X=-0.045 $Y=0 $X2=2.53 $Y2=2.7
cc_59 N_GND_M1002_b N_Y_c_432_n 0.00910143f $X=-0.045 $Y=0 $X2=1.425 $Y2=2.33
cc_60 N_GND_M1002_b N_Y_c_433_n 0.00313521f $X=-0.045 $Y=0 $X2=1.565 $Y2=0.865
cc_61 N_GND_c_3_p N_Y_c_433_n 0.0148533f $X=2.355 $Y=0.152 $X2=1.565 $Y2=0.865
cc_62 N_GND_c_4_p N_Y_c_433_n 0.00955743f $X=2.38 $Y=0.19 $X2=1.565 $Y2=0.865
cc_63 N_GND_M1002_b Y 0.00678007f $X=-0.045 $Y=0 $X2=1.425 $Y2=2.17
cc_64 N_GND_M1002_b N_Y_c_437_n 0.00252706f $X=-0.045 $Y=0 $X2=1.425 $Y2=2.33
cc_65 N_GND_M1002_b N_Y_c_438_n 0.00176349f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.22
cc_66 N_GND_c_2_p N_Y_c_438_n 3.91112e-19 $X=0.69 $Y=0.865 $X2=1.425 $Y2=1.22
cc_67 N_VDD_M1001_b N_A_27_115#_M1010_g 0.0204171f $X=-0.045 $Y=2.645 $X2=1.865
+ $Y2=3.825
cc_68 N_VDD_c_68_p N_A_27_115#_M1010_g 0.00496961f $X=2.355 $Y=5.397 $X2=1.865
+ $Y2=3.825
cc_69 N_VDD_c_69_p N_A_27_115#_M1010_g 0.00429146f $X=2.38 $Y=5.36 $X2=1.865
+ $Y2=3.825
cc_70 N_VDD_M1001_b N_A_27_115#_c_118_n 0.00494544f $X=-0.045 $Y=2.645 $X2=1.805
+ $Y2=2.505
cc_71 N_VDD_M1001_b N_A_27_115#_c_122_n 0.010711f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.205
cc_72 N_VDD_c_72_p N_A_27_115#_c_122_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.205
cc_73 N_VDD_c_69_p N_A_27_115#_c_122_n 0.00435496f $X=2.38 $Y=5.36 $X2=0.26
+ $Y2=3.205
cc_74 N_VDD_M1001_b N_A_27_115#_c_124_n 9.80914e-19 $X=-0.045 $Y=2.645 $X2=1.805
+ $Y2=2.505
cc_75 N_VDD_M1001_b N_A_c_206_n 0.0187048f $X=-0.045 $Y=2.645 $X2=0.475 $Y2=2.75
cc_76 N_VDD_c_72_p N_A_c_206_n 0.00496961f $X=0.605 $Y=5.397 $X2=0.475 $Y2=2.75
cc_77 N_VDD_c_77_p N_A_c_206_n 0.00362996f $X=0.69 $Y=3.885 $X2=0.475 $Y2=2.75
cc_78 N_VDD_c_69_p N_A_c_206_n 0.00429146f $X=2.38 $Y=5.36 $X2=0.475 $Y2=2.75
cc_79 N_VDD_M1001_b N_A_c_189_n 0.00557443f $X=-0.045 $Y=2.645 $X2=0.71
+ $Y2=2.675
cc_80 N_VDD_M1001_b N_A_c_200_n 0.00756323f $X=-0.045 $Y=2.645 $X2=0.45
+ $Y2=2.675
cc_81 N_VDD_M1001_b N_A_c_201_n 0.00635728f $X=-0.045 $Y=2.645 $X2=0.845
+ $Y2=2.505
cc_82 N_VDD_M1001_b N_A_c_213_n 0.0140256f $X=-0.045 $Y=2.645 $X2=0.845 $Y2=2.75
cc_83 N_VDD_c_77_p N_A_c_213_n 0.00362996f $X=0.69 $Y=3.885 $X2=0.845 $Y2=2.75
cc_84 N_VDD_c_68_p N_A_c_213_n 0.00496961f $X=2.355 $Y=5.397 $X2=0.845 $Y2=2.75
cc_85 N_VDD_c_69_p N_A_c_213_n 0.00429146f $X=2.38 $Y=5.36 $X2=0.845 $Y2=2.75
cc_86 N_VDD_M1001_d N_A_c_217_n 0.00200838f $X=0.55 $Y=2.825 $X2=0.845 $Y2=2.985
cc_87 N_VDD_M1001_b N_A_c_217_n 6.29066e-19 $X=-0.045 $Y=2.645 $X2=0.845
+ $Y2=2.985
cc_88 N_VDD_M1001_b N_A_c_203_n 0.00153939f $X=-0.045 $Y=2.645 $X2=2.145
+ $Y2=3.07
cc_89 N_VDD_M1001_d N_A_c_220_n 0.00237538f $X=0.55 $Y=2.825 $X2=1.085 $Y2=3.07
cc_90 N_VDD_c_77_p N_A_c_220_n 4.80344e-19 $X=0.69 $Y=3.885 $X2=1.085 $Y2=3.07
cc_91 N_VDD_M1001_b N_A_238_89#_M1006_g 0.0217118f $X=-0.045 $Y=2.645 $X2=1.265
+ $Y2=3.825
cc_92 N_VDD_c_68_p N_A_238_89#_M1006_g 0.00496961f $X=2.355 $Y=5.397 $X2=1.265
+ $Y2=3.825
cc_93 N_VDD_c_69_p N_A_238_89#_M1006_g 0.00429146f $X=2.38 $Y=5.36 $X2=1.265
+ $Y2=3.825
cc_94 N_VDD_M1001_b N_A_238_89#_c_319_n 0.0101605f $X=-0.045 $Y=2.645 $X2=2.87
+ $Y2=3.205
cc_95 N_VDD_c_95_p N_A_238_89#_c_319_n 0.00477009f $X=2.38 $Y=5.36 $X2=2.87
+ $Y2=3.205
cc_96 N_VDD_c_69_p N_A_238_89#_c_319_n 0.00435496f $X=2.38 $Y=5.36 $X2=2.87
+ $Y2=3.205
cc_97 N_VDD_M1001_b N_B_c_389_n 0.0137488f $X=-0.045 $Y=2.645 $X2=2.225 $Y2=2.75
cc_98 N_VDD_c_68_p N_B_c_389_n 0.00496961f $X=2.355 $Y=5.397 $X2=2.225 $Y2=2.75
cc_99 N_VDD_c_99_p N_B_c_389_n 0.00362996f $X=2.44 $Y=3.885 $X2=2.225 $Y2=2.75
cc_100 N_VDD_c_69_p N_B_c_389_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.225 $Y2=2.75
cc_101 N_VDD_M1001_b N_B_c_393_n 0.0184556f $X=-0.045 $Y=2.645 $X2=2.655
+ $Y2=2.75
cc_102 N_VDD_c_99_p N_B_c_393_n 0.00362996f $X=2.44 $Y=3.885 $X2=2.655 $Y2=2.75
cc_103 N_VDD_c_95_p N_B_c_393_n 0.00496961f $X=2.38 $Y=5.36 $X2=2.655 $Y2=2.75
cc_104 N_VDD_c_69_p N_B_c_393_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.655 $Y2=2.75
cc_105 N_VDD_M1001_b N_B_c_385_n 0.0132516f $X=-0.045 $Y=2.645 $X2=2.655
+ $Y2=2.545
cc_106 N_VDD_M1001_b N_B_c_387_n 0.00187626f $X=-0.045 $Y=2.645 $X2=2.53
+ $Y2=2.505
cc_107 N_VDD_M1001_b B 0.0105467f $X=-0.045 $Y=2.645 $X2=2.53 $Y2=2.7
cc_108 N_VDD_M1001_b N_Y_c_432_n 0.00419006f $X=-0.045 $Y=2.645 $X2=1.425
+ $Y2=2.33
cc_109 N_VDD_M1001_b N_Y_c_441_n 0.00402069f $X=-0.045 $Y=2.645 $X2=1.565
+ $Y2=3.205
cc_110 N_VDD_c_68_p N_Y_c_441_n 0.00925108f $X=2.355 $Y=5.397 $X2=1.565
+ $Y2=3.205
cc_111 N_VDD_c_69_p N_Y_c_441_n 0.00876183f $X=2.38 $Y=5.36 $X2=1.565 $Y2=3.205
cc_112 N_A_27_115#_M1000_g N_A_c_188_n 0.010446f $X=0.905 $Y=0.945 $X2=0.425
+ $Y2=2.6
cc_113 N_A_27_115#_c_116_n N_A_c_188_n 0.0212638f $X=0.845 $Y=1.965 $X2=0.425
+ $Y2=2.6
cc_114 N_A_27_115#_c_122_n N_A_c_188_n 0.0250234f $X=0.26 $Y=3.205 $X2=0.425
+ $Y2=2.6
cc_115 N_A_27_115#_c_123_n N_A_c_188_n 0.0200248f $X=1.72 $Y=1.965 $X2=0.425
+ $Y2=2.6
cc_116 N_A_27_115#_c_122_n N_A_c_206_n 0.00665557f $X=0.26 $Y=3.205 $X2=0.475
+ $Y2=2.75
cc_117 N_A_27_115#_c_123_n N_A_c_189_n 8.37626e-19 $X=1.72 $Y=1.965 $X2=0.71
+ $Y2=2.675
cc_118 N_A_27_115#_c_118_n N_A_c_194_n 0.00428847f $X=1.805 $Y=2.505 $X2=1.94
+ $Y2=1.825
cc_119 N_A_27_115#_c_123_n N_A_c_194_n 0.00407778f $X=1.72 $Y=1.965 $X2=1.94
+ $Y2=1.825
cc_120 N_A_27_115#_M1000_g N_A_c_195_n 0.0279575f $X=0.905 $Y=0.945 $X2=0.45
+ $Y2=1.39
cc_121 N_A_27_115#_c_119_n N_A_c_195_n 0.00957633f $X=0.26 $Y=0.865 $X2=0.45
+ $Y2=1.39
cc_122 N_A_27_115#_c_119_n N_A_c_199_n 0.0202283f $X=0.26 $Y=0.865 $X2=0.45
+ $Y2=1.515
cc_123 N_A_27_115#_c_123_n N_A_c_199_n 0.00168707f $X=1.72 $Y=1.965 $X2=0.45
+ $Y2=1.515
cc_124 N_A_27_115#_c_116_n N_A_c_201_n 0.0184982f $X=0.845 $Y=1.965 $X2=0.845
+ $Y2=2.505
cc_125 N_A_27_115#_c_123_n N_A_c_201_n 9.97344e-19 $X=1.72 $Y=1.965 $X2=0.845
+ $Y2=2.505
cc_126 N_A_27_115#_c_123_n N_A_c_202_n 0.0010613f $X=1.72 $Y=1.965 $X2=2.235
+ $Y2=1.825
cc_127 N_A_27_115#_c_124_n N_A_c_202_n 4.73221e-19 $X=1.805 $Y=2.505 $X2=2.235
+ $Y2=1.825
cc_128 N_A_27_115#_c_122_n N_A_c_217_n 0.0118732f $X=0.26 $Y=3.205 $X2=0.845
+ $Y2=2.985
cc_129 N_A_27_115#_c_118_n N_A_c_203_n 0.00657692f $X=1.805 $Y=2.505 $X2=2.145
+ $Y2=3.07
cc_130 N_A_27_115#_c_123_n N_A_c_203_n 4.20036e-19 $X=1.72 $Y=1.965 $X2=2.145
+ $Y2=3.07
cc_131 N_A_27_115#_c_124_n N_A_c_203_n 0.0441291f $X=1.805 $Y=2.505 $X2=2.145
+ $Y2=3.07
cc_132 N_A_27_115#_c_116_n N_A_c_204_n 9.48646e-19 $X=0.845 $Y=1.965 $X2=0.845
+ $Y2=2.505
cc_133 N_A_27_115#_c_122_n N_A_c_204_n 0.00840379f $X=0.26 $Y=3.205 $X2=0.845
+ $Y2=2.505
cc_134 N_A_27_115#_c_123_n N_A_c_204_n 0.0130076f $X=1.72 $Y=1.965 $X2=0.845
+ $Y2=2.505
cc_135 N_A_27_115#_c_123_n N_A_c_205_n 0.0140397f $X=1.72 $Y=1.965 $X2=2.235
+ $Y2=1.96
cc_136 N_A_27_115#_M1010_g N_A_c_246_n 0.0126423f $X=1.865 $Y=3.825 $X2=2
+ $Y2=3.07
cc_137 N_A_27_115#_c_124_n N_A_c_246_n 0.00625535f $X=1.805 $Y=2.505 $X2=2
+ $Y2=3.07
cc_138 N_A_27_115#_c_122_n N_A_c_248_n 0.00186628f $X=0.26 $Y=3.205 $X2=1.23
+ $Y2=3.07
cc_139 N_A_27_115#_M1010_g N_A_c_249_n 9.56269e-19 $X=1.865 $Y=3.825 $X2=2.145
+ $Y2=3.07
cc_140 N_A_27_115#_M1010_g N_A_238_89#_M1006_g 0.0432496f $X=1.865 $Y=3.825
+ $X2=1.265 $Y2=3.825
cc_141 N_A_27_115#_c_118_n N_A_238_89#_M1006_g 0.0104023f $X=1.805 $Y=2.505
+ $X2=1.265 $Y2=3.825
cc_142 N_A_27_115#_c_123_n N_A_238_89#_M1006_g 0.0147853f $X=1.72 $Y=1.965
+ $X2=1.265 $Y2=3.825
cc_143 N_A_27_115#_c_124_n N_A_238_89#_M1006_g 0.00467915f $X=1.805 $Y=2.505
+ $X2=1.265 $Y2=3.825
cc_144 N_A_27_115#_c_116_n N_A_238_89#_c_311_n 0.052311f $X=0.845 $Y=1.965
+ $X2=1.325 $Y2=1.59
cc_145 N_A_27_115#_c_123_n N_A_238_89#_c_311_n 0.00220335f $X=1.72 $Y=1.965
+ $X2=1.325 $Y2=1.59
cc_146 N_A_27_115#_M1000_g N_A_238_89#_c_312_n 0.052311f $X=0.905 $Y=0.945
+ $X2=1.325 $Y2=1.425
cc_147 N_A_27_115#_M1000_g N_A_238_89#_c_315_n 0.00444529f $X=0.905 $Y=0.945
+ $X2=2.785 $Y2=1.59
cc_148 N_A_27_115#_c_118_n N_A_238_89#_c_315_n 5.57661e-19 $X=1.805 $Y=2.505
+ $X2=2.785 $Y2=1.59
cc_149 N_A_27_115#_c_123_n N_A_238_89#_c_315_n 0.0449127f $X=1.72 $Y=1.965
+ $X2=2.785 $Y2=1.59
cc_150 N_A_27_115#_M1010_g N_B_c_389_n 0.0706461f $X=1.865 $Y=3.825 $X2=2.225
+ $Y2=2.75
cc_151 N_A_27_115#_c_118_n N_B_c_385_n 0.0757008f $X=1.805 $Y=2.505 $X2=2.655
+ $Y2=2.545
cc_152 N_A_27_115#_M1010_g N_Y_c_432_n 0.00249536f $X=1.865 $Y=3.825 $X2=1.425
+ $Y2=2.33
cc_153 N_A_27_115#_c_118_n N_Y_c_432_n 0.00232323f $X=1.805 $Y=2.505 $X2=1.425
+ $Y2=2.33
cc_154 N_A_27_115#_c_123_n N_Y_c_432_n 0.0106304f $X=1.72 $Y=1.965 $X2=1.425
+ $Y2=2.33
cc_155 N_A_27_115#_c_124_n N_Y_c_432_n 0.0239314f $X=1.805 $Y=2.505 $X2=1.425
+ $Y2=2.33
cc_156 N_A_27_115#_M1010_g N_Y_c_448_n 0.0120844f $X=1.865 $Y=3.825 $X2=1.537
+ $Y2=3.115
cc_157 N_A_27_115#_c_118_n N_Y_c_448_n 0.00211862f $X=1.805 $Y=2.505 $X2=1.537
+ $Y2=3.115
cc_158 N_A_27_115#_c_124_n N_Y_c_448_n 6.46587e-19 $X=1.805 $Y=2.505 $X2=1.537
+ $Y2=3.115
cc_159 N_A_27_115#_M1000_g Y 0.00162478f $X=0.905 $Y=0.945 $X2=1.425 $Y2=2.17
cc_160 N_A_27_115#_c_123_n Y 0.0149378f $X=1.72 $Y=1.965 $X2=1.425 $Y2=2.17
cc_161 N_A_27_115#_c_124_n Y 0.00729051f $X=1.805 $Y=2.505 $X2=1.425 $Y2=2.17
cc_162 N_A_27_115#_c_118_n N_Y_c_437_n 0.00177801f $X=1.805 $Y=2.505 $X2=1.425
+ $Y2=2.33
cc_163 N_A_27_115#_c_123_n N_Y_c_437_n 0.00529564f $X=1.72 $Y=1.965 $X2=1.425
+ $Y2=2.33
cc_164 N_A_27_115#_c_124_n N_Y_c_437_n 0.00741445f $X=1.805 $Y=2.505 $X2=1.425
+ $Y2=2.33
cc_165 N_A_27_115#_M1000_g N_Y_c_438_n 0.00127075f $X=0.905 $Y=0.945 $X2=1.425
+ $Y2=1.22
cc_166 N_A_c_188_n N_A_238_89#_M1006_g 0.00462097f $X=0.425 $Y=2.6 $X2=1.265
+ $Y2=3.825
cc_167 N_A_c_194_n N_A_238_89#_M1006_g 0.00424093f $X=1.94 $Y=1.825 $X2=1.265
+ $Y2=3.825
cc_168 N_A_c_201_n N_A_238_89#_M1006_g 0.157467f $X=0.845 $Y=2.505 $X2=1.265
+ $Y2=3.825
cc_169 N_A_c_217_n N_A_238_89#_M1006_g 0.00122231f $X=0.845 $Y=2.985 $X2=1.265
+ $Y2=3.825
cc_170 N_A_c_204_n N_A_238_89#_M1006_g 0.00120277f $X=0.845 $Y=2.505 $X2=1.265
+ $Y2=3.825
cc_171 N_A_c_220_n N_A_238_89#_M1006_g 7.7948e-19 $X=1.085 $Y=3.07 $X2=1.265
+ $Y2=3.825
cc_172 N_A_c_246_n N_A_238_89#_M1006_g 0.00913315f $X=2 $Y=3.07 $X2=1.265
+ $Y2=3.825
cc_173 N_A_c_248_n N_A_238_89#_M1006_g 0.00504822f $X=1.23 $Y=3.07 $X2=1.265
+ $Y2=3.825
cc_174 N_A_M1007_g N_A_238_89#_c_311_n 0.0126897f $X=1.865 $Y=0.945 $X2=1.325
+ $Y2=1.59
cc_175 N_A_M1007_g N_A_238_89#_c_312_n 0.0210321f $X=1.865 $Y=0.945 $X2=1.325
+ $Y2=1.425
cc_176 N_A_M1007_g N_A_238_89#_c_315_n 0.0169961f $X=1.865 $Y=0.945 $X2=2.785
+ $Y2=1.59
cc_177 N_A_c_193_n N_A_238_89#_c_315_n 0.00822635f $X=2.1 $Y=1.825 $X2=2.785
+ $Y2=1.59
cc_178 N_A_c_205_n N_A_238_89#_c_315_n 0.0216132f $X=2.235 $Y=1.96 $X2=2.785
+ $Y2=1.59
cc_179 N_A_c_203_n N_A_238_89#_c_319_n 0.0129458f $X=2.145 $Y=3.07 $X2=2.87
+ $Y2=3.205
cc_180 N_A_c_205_n N_A_238_89#_c_319_n 0.00757462f $X=2.235 $Y=1.96 $X2=2.87
+ $Y2=3.205
cc_181 N_A_c_249_n N_A_238_89#_c_319_n 0.00547471f $X=2.145 $Y=3.07 $X2=2.87
+ $Y2=3.205
cc_182 N_A_M1007_g N_B_c_374_n 0.0673936f $X=1.865 $Y=0.945 $X2=2.225 $Y2=1.39
cc_183 N_A_c_203_n N_B_c_389_n 0.0110965f $X=2.145 $Y=3.07 $X2=2.225 $Y2=2.75
cc_184 N_A_c_249_n N_B_c_389_n 0.0108195f $X=2.145 $Y=3.07 $X2=2.225 $Y2=2.75
cc_185 N_A_c_202_n N_B_c_380_n 0.0137512f $X=2.235 $Y=1.825 $X2=2.3 $Y2=1.465
cc_186 N_A_M1007_g N_B_c_384_n 0.00230834f $X=1.865 $Y=0.945 $X2=2.655 $Y2=2.34
cc_187 N_A_c_202_n N_B_c_384_n 0.0234824f $X=2.235 $Y=1.825 $X2=2.655 $Y2=2.34
cc_188 N_A_c_203_n N_B_c_384_n 0.00252389f $X=2.145 $Y=3.07 $X2=2.655 $Y2=2.34
cc_189 N_A_c_205_n N_B_c_384_n 0.00130506f $X=2.235 $Y=1.96 $X2=2.655 $Y2=2.34
cc_190 N_A_c_203_n N_B_c_393_n 0.00146094f $X=2.145 $Y=3.07 $X2=2.655 $Y2=2.75
cc_191 N_A_c_249_n N_B_c_393_n 0.00122438f $X=2.145 $Y=3.07 $X2=2.655 $Y2=2.75
cc_192 N_A_c_202_n N_B_c_385_n 0.0057573f $X=2.235 $Y=1.825 $X2=2.655 $Y2=2.545
cc_193 N_A_c_203_n N_B_c_385_n 0.00757946f $X=2.145 $Y=3.07 $X2=2.655 $Y2=2.545
cc_194 N_A_c_205_n N_B_c_385_n 0.0016552f $X=2.235 $Y=1.96 $X2=2.655 $Y2=2.545
cc_195 N_A_c_203_n N_B_c_387_n 0.0237616f $X=2.145 $Y=3.07 $X2=2.53 $Y2=2.505
cc_196 N_A_c_202_n B 5.32411e-19 $X=2.235 $Y=1.825 $X2=2.53 $Y2=2.7
cc_197 N_A_c_203_n B 0.00707785f $X=2.145 $Y=3.07 $X2=2.53 $Y2=2.7
cc_198 N_A_c_205_n B 0.00327406f $X=2.235 $Y=1.96 $X2=2.53 $Y2=2.7
cc_199 N_A_c_249_n B 0.00136805f $X=2.145 $Y=3.07 $X2=2.53 $Y2=2.7
cc_200 N_A_c_220_n A_196_565# 0.00327132f $X=1.085 $Y=3.07 $X2=0.98 $Y2=2.825
cc_201 N_A_c_248_n A_196_565# 0.0158919f $X=1.23 $Y=3.07 $X2=0.98 $Y2=2.825
cc_202 N_A_c_246_n N_Y_M1006_d 0.00470028f $X=2 $Y=3.07 $X2=1.34 $Y2=2.825
cc_203 N_A_c_217_n N_Y_c_432_n 0.0110423f $X=0.845 $Y=2.985 $X2=1.425 $Y2=2.33
cc_204 N_A_c_203_n N_Y_c_432_n 0.00873529f $X=2.145 $Y=3.07 $X2=1.425 $Y2=2.33
cc_205 N_A_c_204_n N_Y_c_432_n 0.00811087f $X=0.845 $Y=2.505 $X2=1.425 $Y2=2.33
cc_206 N_A_M1007_g N_Y_c_462_n 0.00296624f $X=1.865 $Y=0.945 $X2=1.565 $Y2=0.985
cc_207 N_A_c_220_n N_Y_c_441_n 0.00106197f $X=1.085 $Y=3.07 $X2=1.565 $Y2=3.205
cc_208 N_A_c_246_n N_Y_c_441_n 0.020967f $X=2 $Y=3.07 $X2=1.565 $Y2=3.205
cc_209 N_A_c_248_n N_Y_c_441_n 0.00145646f $X=1.23 $Y=3.07 $X2=1.565 $Y2=3.205
cc_210 N_A_c_249_n N_Y_c_441_n 0.00142425f $X=2.145 $Y=3.07 $X2=1.565 $Y2=3.205
cc_211 N_A_c_203_n N_Y_c_448_n 0.00530707f $X=2.145 $Y=3.07 $X2=1.537 $Y2=3.115
cc_212 N_A_c_220_n N_Y_c_448_n 0.00470321f $X=1.085 $Y=3.07 $X2=1.537 $Y2=3.115
cc_213 N_A_c_246_n N_Y_c_448_n 0.0217901f $X=2 $Y=3.07 $X2=1.537 $Y2=3.115
cc_214 N_A_c_248_n N_Y_c_448_n 9.55407e-19 $X=1.23 $Y=3.07 $X2=1.537 $Y2=3.115
cc_215 N_A_c_249_n N_Y_c_448_n 8.57579e-19 $X=2.145 $Y=3.07 $X2=1.537 $Y2=3.115
cc_216 N_A_M1007_g Y 0.00504329f $X=1.865 $Y=0.945 $X2=1.425 $Y2=2.17
cc_217 N_A_c_203_n Y 2.67392e-19 $X=2.145 $Y=3.07 $X2=1.425 $Y2=2.17
cc_218 N_A_c_205_n Y 7.53753e-19 $X=2.235 $Y=1.96 $X2=1.425 $Y2=2.17
cc_219 N_A_c_201_n N_Y_c_437_n 3.98944e-19 $X=0.845 $Y=2.505 $X2=1.425 $Y2=2.33
cc_220 N_A_c_204_n N_Y_c_437_n 6.11977e-19 $X=0.845 $Y=2.505 $X2=1.425 $Y2=2.33
cc_221 N_A_c_246_n N_Y_c_437_n 0.0126696f $X=2 $Y=3.07 $X2=1.425 $Y2=2.33
cc_222 N_A_M1007_g N_Y_c_438_n 0.00334017f $X=1.865 $Y=0.945 $X2=1.425 $Y2=1.22
cc_223 N_A_c_203_n A_388_565# 0.003952f $X=2.145 $Y=3.07 $X2=1.94 $Y2=2.825
cc_224 N_A_c_246_n A_388_565# 0.00457146f $X=2 $Y=3.07 $X2=1.94 $Y2=2.825
cc_225 N_A_c_249_n A_388_565# 0.00897914f $X=2.145 $Y=3.07 $X2=1.94 $Y2=2.825
cc_226 N_A_238_89#_c_315_n N_B_c_378_n 0.0123371f $X=2.785 $Y=1.59 $X2=2.58
+ $Y2=1.465
cc_227 N_A_238_89#_c_315_n N_B_c_380_n 0.00821444f $X=2.785 $Y=1.59 $X2=2.3
+ $Y2=1.465
cc_228 N_A_238_89#_c_317_n N_B_c_381_n 0.0148161f $X=2.87 $Y=0.865 $X2=2.655
+ $Y2=1.39
cc_229 N_A_238_89#_c_315_n N_B_c_384_n 0.0113699f $X=2.785 $Y=1.59 $X2=2.655
+ $Y2=2.34
cc_230 N_A_238_89#_c_319_n N_B_c_384_n 0.0382539f $X=2.87 $Y=3.205 $X2=2.655
+ $Y2=2.34
cc_231 N_A_238_89#_c_315_n N_B_c_385_n 0.00171569f $X=2.785 $Y=1.59 $X2=2.655
+ $Y2=2.545
cc_232 N_A_238_89#_c_315_n N_B_c_386_n 0.00775577f $X=2.785 $Y=1.59 $X2=2.655
+ $Y2=1.465
cc_233 N_A_238_89#_c_315_n N_B_c_387_n 0.00443258f $X=2.785 $Y=1.59 $X2=2.53
+ $Y2=2.505
cc_234 N_A_238_89#_c_319_n N_B_c_387_n 0.0299635f $X=2.87 $Y=3.205 $X2=2.53
+ $Y2=2.505
cc_235 N_A_238_89#_c_319_n B 0.00657877f $X=2.87 $Y=3.205 $X2=2.53 $Y2=2.7
cc_236 N_A_238_89#_M1006_g N_Y_c_432_n 0.0124336f $X=1.265 $Y=3.825 $X2=1.425
+ $Y2=2.33
cc_237 N_A_238_89#_c_311_n N_Y_c_462_n 0.00100251f $X=1.325 $Y=1.59 $X2=1.565
+ $Y2=0.985
cc_238 N_A_238_89#_c_312_n N_Y_c_462_n 0.00394924f $X=1.325 $Y=1.425 $X2=1.565
+ $Y2=0.985
cc_239 N_A_238_89#_c_315_n N_Y_c_462_n 0.0151305f $X=2.785 $Y=1.59 $X2=1.565
+ $Y2=0.985
cc_240 N_A_238_89#_M1006_g N_Y_c_441_n 0.0108074f $X=1.265 $Y=3.825 $X2=1.565
+ $Y2=3.205
cc_241 N_A_238_89#_M1006_g Y 0.00604691f $X=1.265 $Y=3.825 $X2=1.425 $Y2=2.17
cc_242 N_A_238_89#_c_311_n Y 0.00612713f $X=1.325 $Y=1.59 $X2=1.425 $Y2=2.17
cc_243 N_A_238_89#_c_315_n Y 0.0165787f $X=2.785 $Y=1.59 $X2=1.425 $Y2=2.17
cc_244 N_A_238_89#_M1006_g N_Y_c_437_n 0.00966885f $X=1.265 $Y=3.825 $X2=1.425
+ $Y2=2.33
cc_245 N_A_238_89#_c_312_n N_Y_c_438_n 0.0053972f $X=1.325 $Y=1.425 $X2=1.425
+ $Y2=1.22
cc_246 N_A_238_89#_c_315_n N_Y_c_438_n 0.00572048f $X=2.785 $Y=1.59 $X2=1.425
+ $Y2=1.22
