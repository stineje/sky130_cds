magic
tech sky130A
magscale 1 2
timestamp 1612372068
<< nwell >>
rect -9 529 376 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 252 115 282 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 166 243
rect 110 131 121 215
rect 155 131 166 215
rect 110 115 166 131
rect 196 215 252 243
rect 196 131 207 215
rect 241 131 252 215
rect 196 115 252 131
rect 282 215 335 243
rect 282 131 293 215
rect 327 131 335 215
rect 282 115 335 131
<< pdiff >>
rect 27 949 80 965
rect 27 605 35 949
rect 69 605 80 949
rect 27 565 80 605
rect 110 949 166 965
rect 110 741 121 949
rect 155 741 166 949
rect 110 565 166 741
rect 196 949 252 965
rect 196 605 207 949
rect 241 605 252 949
rect 196 565 252 605
rect 282 949 335 965
rect 282 605 293 949
rect 327 605 335 949
rect 282 565 335 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 207 131 241 215
rect 293 131 327 215
<< pdiffc >>
rect 35 605 69 949
rect 121 741 155 949
rect 207 605 241 949
rect 293 605 327 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 992
rect 80 477 110 565
rect 166 550 196 565
rect 252 550 282 565
rect 166 520 282 550
rect 80 461 154 477
rect 80 427 110 461
rect 144 427 154 461
rect 80 411 154 427
rect 80 243 110 411
rect 221 368 251 520
rect 166 352 251 368
rect 166 318 176 352
rect 210 332 251 352
rect 210 318 282 332
rect 166 302 282 318
rect 166 243 196 302
rect 252 243 282 302
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
<< polycont >>
rect 110 427 144 461
rect 176 318 210 352
<< locali >>
rect 0 1089 374 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 374 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 725 155 741
rect 207 949 241 965
rect 35 352 69 605
rect 110 461 144 597
rect 207 557 241 605
rect 293 949 327 1049
rect 293 589 327 605
rect 110 411 144 427
rect 176 352 210 368
rect 35 318 176 352
rect 35 215 69 318
rect 176 302 210 318
rect 35 115 69 131
rect 121 215 155 231
rect 121 61 155 131
rect 207 215 241 227
rect 207 115 241 131
rect 293 215 327 231
rect 293 61 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 110 597 144 631
rect 207 523 241 557
rect 207 227 241 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 374 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 374 1089
rect 0 1049 374 1055
rect 98 631 156 637
rect 64 597 110 631
rect 144 597 156 631
rect 98 591 156 597
rect 195 557 253 563
rect 195 523 207 557
rect 241 523 253 557
rect 195 517 253 523
rect 207 267 241 517
rect 195 261 253 267
rect 195 227 207 261
rect 241 227 253 261
rect 195 221 253 227
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel viali 127 614 127 614 1 A
port 1 n
rlabel metal1 211 402 211 402 1 Y
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
