* File: sky130_osu_sc_15T_ms__inv_8.pxi.spice
* Created: Fri Nov 12 14:44:36 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__INV_8%GND N_GND_M1001_d N_GND_M1003_d N_GND_M1009_d
+ N_GND_M1011_d N_GND_M1013_d N_GND_M1001_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p
+ N_GND_c_17_p N_GND_c_23_p N_GND_c_30_p N_GND_c_37_p N_GND_c_44_p N_GND_c_50_p
+ GND N_GND_c_4_p PM_SKY130_OSU_SC_15T_MS__INV_8%GND
x_PM_SKY130_OSU_SC_15T_MS__INV_8%VDD N_VDD_M1000_d N_VDD_M1002_d N_VDD_M1005_d
+ N_VDD_M1008_d N_VDD_M1015_d N_VDD_M1000_b N_VDD_c_112_p N_VDD_c_113_p
+ N_VDD_c_118_p N_VDD_c_124_p N_VDD_c_129_p N_VDD_c_135_p N_VDD_c_140_p
+ N_VDD_c_146_p N_VDD_c_151_p VDD N_VDD_c_114_p
+ PM_SKY130_OSU_SC_15T_MS__INV_8%VDD
x_PM_SKY130_OSU_SC_15T_MS__INV_8%A N_A_c_188_n N_A_M1001_g N_A_c_192_n
+ N_A_c_258_n N_A_M1000_g N_A_c_193_n N_A_c_194_n N_A_c_195_n N_A_M1003_g
+ N_A_c_263_n N_A_M1002_g N_A_c_199_n N_A_c_201_n N_A_c_202_n N_A_M1007_g
+ N_A_c_269_n N_A_M1004_g N_A_c_206_n N_A_c_207_n N_A_c_208_n N_A_M1009_g
+ N_A_c_274_n N_A_M1005_g N_A_c_212_n N_A_c_214_n N_A_c_215_n N_A_M1010_g
+ N_A_c_219_n N_A_c_280_n N_A_M1006_g N_A_c_220_n N_A_c_221_n N_A_c_222_n
+ N_A_M1011_g N_A_c_285_n N_A_M1008_g N_A_c_226_n N_A_c_228_n N_A_c_229_n
+ N_A_M1012_g N_A_c_291_n N_A_M1014_g N_A_c_233_n N_A_c_234_n N_A_c_235_n
+ N_A_M1013_g N_A_c_296_n N_A_M1015_g N_A_c_239_n N_A_c_240_n N_A_c_241_n
+ N_A_c_242_n N_A_c_243_n N_A_c_244_n N_A_c_245_n N_A_c_246_n N_A_c_247_n
+ N_A_c_248_n N_A_c_249_n N_A_c_250_n N_A_c_251_n N_A_c_252_n N_A_c_253_n
+ N_A_c_254_n N_A_c_255_n N_A_c_256_n N_A_c_257_n A
+ PM_SKY130_OSU_SC_15T_MS__INV_8%A
x_PM_SKY130_OSU_SC_15T_MS__INV_8%Y N_Y_M1001_s N_Y_M1007_s N_Y_M1010_s
+ N_Y_M1012_s N_Y_M1000_s N_Y_M1004_s N_Y_M1006_s N_Y_M1014_s N_Y_c_422_n
+ N_Y_c_462_n N_Y_c_426_n N_Y_c_465_n N_Y_c_431_n N_Y_c_468_n N_Y_c_436_n
+ N_Y_c_471_n N_Y_c_440_n N_Y_c_474_n Y N_Y_c_444_n N_Y_c_475_n N_Y_c_446_n
+ N_Y_c_447_n N_Y_c_449_n N_Y_c_477_n N_Y_c_479_n N_Y_c_452_n N_Y_c_453_n
+ N_Y_c_455_n N_Y_c_480_n N_Y_c_482_n N_Y_c_458_n N_Y_c_461_n
+ PM_SKY130_OSU_SC_15T_MS__INV_8%Y
cc_1 N_GND_M1001_b N_A_c_188_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.44
cc_2 N_GND_c_2_p N_A_c_188_n 0.00866533f $X=0.26 $Y=0.865 $X2=0.475 $Y2=1.44
cc_3 N_GND_c_3_p N_A_c_188_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.44
cc_4 N_GND_c_4_p N_A_c_188_n 0.00468827f $X=3.06 $Y=0.19 $X2=0.475 $Y2=1.44
cc_5 N_GND_M1001_b N_A_c_192_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.55
cc_6 N_GND_M1001_b N_A_c_193_n 0.01476f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.515
cc_7 N_GND_M1001_b N_A_c_194_n 0.00981662f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.625
cc_8 N_GND_M1001_b N_A_c_195_n 0.0166526f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.44
cc_9 N_GND_c_3_p N_A_c_195_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.44
cc_10 N_GND_c_10_p N_A_c_195_n 0.00390533f $X=1.12 $Y=0.865 $X2=0.905 $Y2=1.44
cc_11 N_GND_c_4_p N_A_c_195_n 0.00468827f $X=3.06 $Y=0.19 $X2=0.905 $Y2=1.44
cc_12 N_GND_M1001_b N_A_c_199_n 0.0213783f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.515
cc_13 N_GND_c_10_p N_A_c_199_n 0.00283047f $X=1.12 $Y=0.865 $X2=1.26 $Y2=1.515
cc_14 N_GND_M1001_b N_A_c_201_n 0.0173499f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.625
cc_15 N_GND_M1001_b N_A_c_202_n 0.0166526f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.44
cc_16 N_GND_c_10_p N_A_c_202_n 0.00390533f $X=1.12 $Y=0.865 $X2=1.335 $Y2=1.44
cc_17 N_GND_c_17_p N_A_c_202_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.335 $Y2=1.44
cc_18 N_GND_c_4_p N_A_c_202_n 0.00468827f $X=3.06 $Y=0.19 $X2=1.335 $Y2=1.44
cc_19 N_GND_M1001_b N_A_c_206_n 0.0195339f $X=-0.045 $Y=0 $X2=1.69 $Y2=1.515
cc_20 N_GND_M1001_b N_A_c_207_n 0.0145324f $X=-0.045 $Y=0 $X2=1.69 $Y2=2.625
cc_21 N_GND_M1001_b N_A_c_208_n 0.0166526f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.44
cc_22 N_GND_c_17_p N_A_c_208_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.765 $Y2=1.44
cc_23 N_GND_c_23_p N_A_c_208_n 0.00390533f $X=1.98 $Y=0.865 $X2=1.765 $Y2=1.44
cc_24 N_GND_c_4_p N_A_c_208_n 0.00468827f $X=3.06 $Y=0.19 $X2=1.765 $Y2=1.44
cc_25 N_GND_M1001_b N_A_c_212_n 0.0164591f $X=-0.045 $Y=0 $X2=2.12 $Y2=1.515
cc_26 N_GND_c_23_p N_A_c_212_n 0.00283047f $X=1.98 $Y=0.865 $X2=2.12 $Y2=1.515
cc_27 N_GND_M1001_b N_A_c_214_n 0.0124307f $X=-0.045 $Y=0 $X2=2.12 $Y2=2.625
cc_28 N_GND_M1001_b N_A_c_215_n 0.0166526f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.44
cc_29 N_GND_c_23_p N_A_c_215_n 0.00390533f $X=1.98 $Y=0.865 $X2=2.195 $Y2=1.44
cc_30 N_GND_c_30_p N_A_c_215_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.195 $Y2=1.44
cc_31 N_GND_c_4_p N_A_c_215_n 0.00468827f $X=3.06 $Y=0.19 $X2=2.195 $Y2=1.44
cc_32 N_GND_M1001_b N_A_c_219_n 0.0685082f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.55
cc_33 N_GND_M1001_b N_A_c_220_n 0.0195339f $X=-0.045 $Y=0 $X2=2.55 $Y2=1.515
cc_34 N_GND_M1001_b N_A_c_221_n 0.0145324f $X=-0.045 $Y=0 $X2=2.55 $Y2=2.625
cc_35 N_GND_M1001_b N_A_c_222_n 0.0166526f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.44
cc_36 N_GND_c_30_p N_A_c_222_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.625 $Y2=1.44
cc_37 N_GND_c_37_p N_A_c_222_n 0.00390533f $X=2.84 $Y=0.865 $X2=2.625 $Y2=1.44
cc_38 N_GND_c_4_p N_A_c_222_n 0.00468827f $X=3.06 $Y=0.19 $X2=2.625 $Y2=1.44
cc_39 N_GND_M1001_b N_A_c_226_n 0.0213783f $X=-0.045 $Y=0 $X2=2.98 $Y2=1.515
cc_40 N_GND_c_37_p N_A_c_226_n 0.00283047f $X=2.84 $Y=0.865 $X2=2.98 $Y2=1.515
cc_41 N_GND_M1001_b N_A_c_228_n 0.0173499f $X=-0.045 $Y=0 $X2=2.98 $Y2=2.625
cc_42 N_GND_M1001_b N_A_c_229_n 0.0166526f $X=-0.045 $Y=0 $X2=3.055 $Y2=1.44
cc_43 N_GND_c_37_p N_A_c_229_n 0.00390533f $X=2.84 $Y=0.865 $X2=3.055 $Y2=1.44
cc_44 N_GND_c_44_p N_A_c_229_n 0.00606474f $X=3.615 $Y=0.152 $X2=3.055 $Y2=1.44
cc_45 N_GND_c_4_p N_A_c_229_n 0.00468827f $X=3.06 $Y=0.19 $X2=3.055 $Y2=1.44
cc_46 N_GND_M1001_b N_A_c_233_n 0.0385034f $X=-0.045 $Y=0 $X2=3.41 $Y2=1.515
cc_47 N_GND_M1001_b N_A_c_234_n 0.0295863f $X=-0.045 $Y=0 $X2=3.41 $Y2=2.625
cc_48 N_GND_M1001_b N_A_c_235_n 0.0208613f $X=-0.045 $Y=0 $X2=3.485 $Y2=1.44
cc_49 N_GND_c_44_p N_A_c_235_n 0.00606474f $X=3.615 $Y=0.152 $X2=3.485 $Y2=1.44
cc_50 N_GND_c_50_p N_A_c_235_n 0.00866533f $X=3.7 $Y=0.865 $X2=3.485 $Y2=1.44
cc_51 N_GND_c_4_p N_A_c_235_n 0.00468827f $X=3.06 $Y=0.19 $X2=3.485 $Y2=1.44
cc_52 N_GND_M1001_b N_A_c_239_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.515
cc_53 N_GND_M1001_b N_A_c_240_n 0.0382476f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.045
cc_54 N_GND_M1001_b N_A_c_241_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.88
cc_55 N_GND_M1001_b N_A_c_242_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.625
cc_56 N_GND_M1001_b N_A_c_243_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.515
cc_57 N_GND_M1001_b N_A_c_244_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.625
cc_58 N_GND_M1001_b N_A_c_245_n 0.0106787f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.515
cc_59 N_GND_M1001_b N_A_c_246_n 0.00980309f $X=-0.045 $Y=0 $X2=1.335 $Y2=2.625
cc_60 N_GND_M1001_b N_A_c_247_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.515
cc_61 N_GND_M1001_b N_A_c_248_n 0.00980309f $X=-0.045 $Y=0 $X2=1.765 $Y2=2.625
cc_62 N_GND_M1001_b N_A_c_249_n 0.0023879f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.515
cc_63 N_GND_M1001_b N_A_c_250_n 0.00151234f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.625
cc_64 N_GND_M1001_b N_A_c_251_n 0.0106787f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.515
cc_65 N_GND_M1001_b N_A_c_252_n 0.00980309f $X=-0.045 $Y=0 $X2=2.625 $Y2=2.625
cc_66 N_GND_M1001_b N_A_c_253_n 0.0106787f $X=-0.045 $Y=0 $X2=3.055 $Y2=1.515
cc_67 N_GND_M1001_b N_A_c_254_n 0.00980309f $X=-0.045 $Y=0 $X2=3.055 $Y2=2.625
cc_68 N_GND_M1001_b N_A_c_255_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.07
cc_69 N_GND_M1001_b N_A_c_256_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.045
cc_70 N_GND_M1001_b N_A_c_257_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.045
cc_71 N_GND_M1001_b N_Y_c_422_n 0.00155118f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.865
cc_72 N_GND_c_3_p N_Y_c_422_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.865
cc_73 N_GND_c_10_p N_Y_c_422_n 8.14297e-19 $X=1.12 $Y=0.865 $X2=0.69 $Y2=0.865
cc_74 N_GND_c_4_p N_Y_c_422_n 0.00475776f $X=3.06 $Y=0.19 $X2=0.69 $Y2=0.865
cc_75 N_GND_M1001_b N_Y_c_426_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.865
cc_76 N_GND_c_10_p N_Y_c_426_n 8.14297e-19 $X=1.12 $Y=0.865 $X2=1.55 $Y2=0.865
cc_77 N_GND_c_17_p N_Y_c_426_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.865
cc_78 N_GND_c_23_p N_Y_c_426_n 8.14297e-19 $X=1.98 $Y=0.865 $X2=1.55 $Y2=0.865
cc_79 N_GND_c_4_p N_Y_c_426_n 0.00475776f $X=3.06 $Y=0.19 $X2=1.55 $Y2=0.865
cc_80 N_GND_M1001_b N_Y_c_431_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.865
cc_81 N_GND_c_23_p N_Y_c_431_n 8.14297e-19 $X=1.98 $Y=0.865 $X2=2.41 $Y2=0.865
cc_82 N_GND_c_30_p N_Y_c_431_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.865
cc_83 N_GND_c_37_p N_Y_c_431_n 8.14297e-19 $X=2.84 $Y=0.865 $X2=2.41 $Y2=0.865
cc_84 N_GND_c_4_p N_Y_c_431_n 0.00475776f $X=3.06 $Y=0.19 $X2=2.41 $Y2=0.865
cc_85 N_GND_M1001_b N_Y_c_436_n 0.00155118f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.865
cc_86 N_GND_c_37_p N_Y_c_436_n 8.14297e-19 $X=2.84 $Y=0.865 $X2=3.27 $Y2=0.865
cc_87 N_GND_c_44_p N_Y_c_436_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.865
cc_88 N_GND_c_4_p N_Y_c_436_n 0.00475776f $X=3.06 $Y=0.19 $X2=3.27 $Y2=0.865
cc_89 N_GND_M1001_b N_Y_c_440_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.335
cc_90 N_GND_c_2_p N_Y_c_440_n 0.00134236f $X=0.26 $Y=0.865 $X2=0.69 $Y2=1.335
cc_91 N_GND_c_10_p N_Y_c_440_n 7.53951e-19 $X=1.12 $Y=0.865 $X2=0.69 $Y2=1.335
cc_92 N_GND_M1001_b Y 0.0456345f $X=-0.045 $Y=0 $X2=0.76 $Y2=1.94
cc_93 N_GND_M1003_d N_Y_c_444_n 0.0127699f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1.22
cc_94 N_GND_c_10_p N_Y_c_444_n 0.0142303f $X=1.12 $Y=0.865 $X2=1.405 $Y2=1.22
cc_95 N_GND_M1001_b N_Y_c_446_n 0.0591815f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.585
cc_96 N_GND_M1009_d N_Y_c_447_n 0.0127699f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.22
cc_97 N_GND_c_23_p N_Y_c_447_n 0.0142303f $X=1.98 $Y=0.865 $X2=2.265 $Y2=1.22
cc_98 N_GND_M1001_b N_Y_c_449_n 0.00409378f $X=-0.045 $Y=0 $X2=1.695 $Y2=1.22
cc_99 N_GND_c_10_p N_Y_c_449_n 7.53951e-19 $X=1.12 $Y=0.865 $X2=1.695 $Y2=1.22
cc_100 N_GND_c_23_p N_Y_c_449_n 7.53951e-19 $X=1.98 $Y=0.865 $X2=1.695 $Y2=1.22
cc_101 N_GND_M1001_b N_Y_c_452_n 0.0580131f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.585
cc_102 N_GND_M1011_d N_Y_c_453_n 0.0127699f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.22
cc_103 N_GND_c_37_p N_Y_c_453_n 0.0142303f $X=2.84 $Y=0.865 $X2=3.125 $Y2=1.22
cc_104 N_GND_M1001_b N_Y_c_455_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.22
cc_105 N_GND_c_23_p N_Y_c_455_n 7.53951e-19 $X=1.98 $Y=0.865 $X2=2.555 $Y2=1.22
cc_106 N_GND_c_37_p N_Y_c_455_n 7.53951e-19 $X=2.84 $Y=0.865 $X2=2.555 $Y2=1.22
cc_107 N_GND_M1001_b N_Y_c_458_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.335
cc_108 N_GND_c_37_p N_Y_c_458_n 7.53951e-19 $X=2.84 $Y=0.865 $X2=3.27 $Y2=1.335
cc_109 N_GND_c_50_p N_Y_c_458_n 0.00134236f $X=3.7 $Y=0.865 $X2=3.27 $Y2=1.335
cc_110 N_GND_M1001_b N_Y_c_461_n 0.0754129f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.585
cc_111 N_VDD_M1000_b N_A_c_258_n 0.0185527f $X=-0.045 $Y=2.645 $X2=0.475 $Y2=2.7
cc_112 N_VDD_c_112_p N_A_c_258_n 0.00751602f $X=0.26 $Y=3.885 $X2=0.475 $Y2=2.7
cc_113 N_VDD_c_113_p N_A_c_258_n 0.00496961f $X=1.035 $Y=5.397 $X2=0.475 $Y2=2.7
cc_114 N_VDD_c_114_p N_A_c_258_n 0.00429146f $X=3.06 $Y=5.36 $X2=0.475 $Y2=2.7
cc_115 N_VDD_M1000_b N_A_c_194_n 0.00448664f $X=-0.045 $Y=2.645 $X2=0.83
+ $Y2=2.625
cc_116 N_VDD_M1000_b N_A_c_263_n 0.0163194f $X=-0.045 $Y=2.645 $X2=0.905 $Y2=2.7
cc_117 N_VDD_c_113_p N_A_c_263_n 0.00496961f $X=1.035 $Y=5.397 $X2=0.905 $Y2=2.7
cc_118 N_VDD_c_118_p N_A_c_263_n 0.00362996f $X=1.12 $Y=3.205 $X2=0.905 $Y2=2.7
cc_119 N_VDD_c_114_p N_A_c_263_n 0.00429146f $X=3.06 $Y=5.36 $X2=0.905 $Y2=2.7
cc_120 N_VDD_M1000_b N_A_c_201_n 0.00500158f $X=-0.045 $Y=2.645 $X2=1.26
+ $Y2=2.625
cc_121 N_VDD_c_118_p N_A_c_201_n 0.00341318f $X=1.12 $Y=3.205 $X2=1.26 $Y2=2.625
cc_122 N_VDD_M1000_b N_A_c_269_n 0.0163194f $X=-0.045 $Y=2.645 $X2=1.335 $Y2=2.7
cc_123 N_VDD_c_118_p N_A_c_269_n 0.00362996f $X=1.12 $Y=3.205 $X2=1.335 $Y2=2.7
cc_124 N_VDD_c_124_p N_A_c_269_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335 $Y2=2.7
cc_125 N_VDD_c_114_p N_A_c_269_n 0.00429146f $X=3.06 $Y=5.36 $X2=1.335 $Y2=2.7
cc_126 N_VDD_M1000_b N_A_c_207_n 0.00448664f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_127 N_VDD_M1000_b N_A_c_274_n 0.0163194f $X=-0.045 $Y=2.645 $X2=1.765 $Y2=2.7
cc_128 N_VDD_c_124_p N_A_c_274_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.765 $Y2=2.7
cc_129 N_VDD_c_129_p N_A_c_274_n 0.00362996f $X=1.98 $Y=3.205 $X2=1.765 $Y2=2.7
cc_130 N_VDD_c_114_p N_A_c_274_n 0.00429146f $X=3.06 $Y=5.36 $X2=1.765 $Y2=2.7
cc_131 N_VDD_M1000_b N_A_c_214_n 0.00500158f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.625
cc_132 N_VDD_c_129_p N_A_c_214_n 0.00341318f $X=1.98 $Y=3.205 $X2=2.12 $Y2=2.625
cc_133 N_VDD_M1000_b N_A_c_280_n 0.0163194f $X=-0.045 $Y=2.645 $X2=2.195 $Y2=2.7
cc_134 N_VDD_c_129_p N_A_c_280_n 0.00362996f $X=1.98 $Y=3.205 $X2=2.195 $Y2=2.7
cc_135 N_VDD_c_135_p N_A_c_280_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.195 $Y2=2.7
cc_136 N_VDD_c_114_p N_A_c_280_n 0.00429146f $X=3.06 $Y=5.36 $X2=2.195 $Y2=2.7
cc_137 N_VDD_M1000_b N_A_c_221_n 0.00448664f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.625
cc_138 N_VDD_M1000_b N_A_c_285_n 0.0163194f $X=-0.045 $Y=2.645 $X2=2.625 $Y2=2.7
cc_139 N_VDD_c_135_p N_A_c_285_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.625 $Y2=2.7
cc_140 N_VDD_c_140_p N_A_c_285_n 0.00362996f $X=2.84 $Y=3.205 $X2=2.625 $Y2=2.7
cc_141 N_VDD_c_114_p N_A_c_285_n 0.00429146f $X=3.06 $Y=5.36 $X2=2.625 $Y2=2.7
cc_142 N_VDD_M1000_b N_A_c_228_n 0.00500158f $X=-0.045 $Y=2.645 $X2=2.98
+ $Y2=2.625
cc_143 N_VDD_c_140_p N_A_c_228_n 0.00341318f $X=2.84 $Y=3.205 $X2=2.98 $Y2=2.625
cc_144 N_VDD_M1000_b N_A_c_291_n 0.0163194f $X=-0.045 $Y=2.645 $X2=3.055 $Y2=2.7
cc_145 N_VDD_c_140_p N_A_c_291_n 0.00362996f $X=2.84 $Y=3.205 $X2=3.055 $Y2=2.7
cc_146 N_VDD_c_146_p N_A_c_291_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.055 $Y2=2.7
cc_147 N_VDD_c_114_p N_A_c_291_n 0.00429146f $X=3.06 $Y=5.36 $X2=3.055 $Y2=2.7
cc_148 N_VDD_M1000_b N_A_c_234_n 0.00840215f $X=-0.045 $Y=2.645 $X2=3.41
+ $Y2=2.625
cc_149 N_VDD_M1000_b N_A_c_296_n 0.0208694f $X=-0.045 $Y=2.645 $X2=3.485 $Y2=2.7
cc_150 N_VDD_c_146_p N_A_c_296_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.485 $Y2=2.7
cc_151 N_VDD_c_151_p N_A_c_296_n 0.00751602f $X=3.7 $Y=3.205 $X2=3.485 $Y2=2.7
cc_152 N_VDD_c_114_p N_A_c_296_n 0.00429146f $X=3.06 $Y=5.36 $X2=3.485 $Y2=2.7
cc_153 N_VDD_M1000_b N_A_c_242_n 0.00244521f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=2.625
cc_154 N_VDD_M1000_b N_A_c_244_n 8.75564e-19 $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=2.625
cc_155 N_VDD_M1000_b N_A_c_246_n 8.75564e-19 $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.625
cc_156 N_VDD_M1000_b N_A_c_248_n 8.75564e-19 $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.625
cc_157 N_VDD_M1000_b N_A_c_250_n 8.75564e-19 $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.625
cc_158 N_VDD_M1000_b N_A_c_252_n 8.75564e-19 $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.625
cc_159 N_VDD_M1000_b N_A_c_254_n 8.75564e-19 $X=-0.045 $Y=2.645 $X2=3.055
+ $Y2=2.625
cc_160 N_VDD_M1000_d N_A_c_255_n 0.00953431f $X=0.135 $Y=2.825 $X2=0.32 $Y2=3.07
cc_161 N_VDD_M1000_b N_A_c_255_n 0.00618364f $X=-0.045 $Y=2.645 $X2=0.32
+ $Y2=3.07
cc_162 N_VDD_c_112_p N_A_c_255_n 0.00252874f $X=0.26 $Y=3.885 $X2=0.32 $Y2=3.07
cc_163 N_VDD_M1000_d A 0.0162774f $X=0.135 $Y=2.825 $X2=0.32 $Y2=3.065
cc_164 N_VDD_c_112_p A 0.00522047f $X=0.26 $Y=3.885 $X2=0.32 $Y2=3.065
cc_165 N_VDD_c_118_p A 9.09141e-19 $X=1.12 $Y=3.205 $X2=0.32 $Y2=3.065
cc_166 N_VDD_M1000_b N_Y_c_462_n 0.00404956f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.7
cc_167 N_VDD_c_113_p N_Y_c_462_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69 $Y2=2.7
cc_168 N_VDD_c_114_p N_Y_c_462_n 0.00434939f $X=3.06 $Y=5.36 $X2=0.69 $Y2=2.7
cc_169 N_VDD_M1000_b N_Y_c_465_n 0.00509484f $X=-0.045 $Y=2.645 $X2=1.55 $Y2=2.7
cc_170 N_VDD_c_124_p N_Y_c_465_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.7
cc_171 N_VDD_c_114_p N_Y_c_465_n 0.00434939f $X=3.06 $Y=5.36 $X2=1.55 $Y2=2.7
cc_172 N_VDD_M1000_b N_Y_c_468_n 0.00509484f $X=-0.045 $Y=2.645 $X2=2.41 $Y2=2.7
cc_173 N_VDD_c_135_p N_Y_c_468_n 0.0045126f $X=2.755 $Y=5.397 $X2=2.41 $Y2=2.7
cc_174 N_VDD_c_114_p N_Y_c_468_n 0.00434939f $X=3.06 $Y=5.36 $X2=2.41 $Y2=2.7
cc_175 N_VDD_M1000_b N_Y_c_471_n 0.00509484f $X=-0.045 $Y=2.645 $X2=3.27 $Y2=2.7
cc_176 N_VDD_c_146_p N_Y_c_471_n 0.00464147f $X=3.615 $Y=5.397 $X2=3.27 $Y2=2.7
cc_177 N_VDD_c_114_p N_Y_c_471_n 0.00434939f $X=3.06 $Y=5.36 $X2=3.27 $Y2=2.7
cc_178 N_VDD_M1000_b N_Y_c_474_n 0.00248543f $X=-0.045 $Y=2.645 $X2=0.69
+ $Y2=2.585
cc_179 N_VDD_M1000_b N_Y_c_475_n 0.00520877f $X=-0.045 $Y=2.645 $X2=1.405
+ $Y2=2.7
cc_180 N_VDD_c_118_p N_Y_c_475_n 0.0090257f $X=1.12 $Y=3.205 $X2=1.405 $Y2=2.7
cc_181 N_VDD_M1000_b N_Y_c_477_n 0.00520877f $X=-0.045 $Y=2.645 $X2=2.265
+ $Y2=2.7
cc_182 N_VDD_c_129_p N_Y_c_477_n 0.0090257f $X=1.98 $Y=3.205 $X2=2.265 $Y2=2.7
cc_183 N_VDD_M1000_b N_Y_c_479_n 0.00409378f $X=-0.045 $Y=2.645 $X2=1.695
+ $Y2=2.7
cc_184 N_VDD_M1000_b N_Y_c_480_n 0.00520877f $X=-0.045 $Y=2.645 $X2=3.125
+ $Y2=2.7
cc_185 N_VDD_c_140_p N_Y_c_480_n 0.0090257f $X=2.84 $Y=3.205 $X2=3.125 $Y2=2.7
cc_186 N_VDD_M1000_b N_Y_c_482_n 0.00409378f $X=-0.045 $Y=2.645 $X2=2.555
+ $Y2=2.7
cc_187 N_VDD_M1000_b N_Y_c_461_n 0.00409378f $X=-0.045 $Y=2.645 $X2=3.27
+ $Y2=2.585
cc_188 A N_Y_M1000_s 0.00251573f $X=0.32 $Y=3.065 $X2=0.55 $Y2=2.825
cc_189 N_A_c_188_n N_Y_c_422_n 0.00265306f $X=0.475 $Y=1.44 $X2=0.69 $Y2=0.865
cc_190 N_A_c_193_n N_Y_c_422_n 0.00256118f $X=0.83 $Y=1.515 $X2=0.69 $Y2=0.865
cc_191 N_A_c_195_n N_Y_c_422_n 0.00265306f $X=0.905 $Y=1.44 $X2=0.69 $Y2=0.865
cc_192 N_A_c_240_n N_Y_c_422_n 3.64468e-19 $X=0.535 $Y=2.045 $X2=0.69 $Y2=0.865
cc_193 N_A_c_257_n N_Y_c_422_n 0.00110256f $X=0.535 $Y=2.045 $X2=0.69 $Y2=0.865
cc_194 N_A_c_258_n N_Y_c_462_n 0.00206894f $X=0.475 $Y=2.7 $X2=0.69 $Y2=2.7
cc_195 N_A_c_194_n N_Y_c_462_n 0.00899372f $X=0.83 $Y=2.625 $X2=0.69 $Y2=2.7
cc_196 N_A_c_263_n N_Y_c_462_n 0.00360548f $X=0.905 $Y=2.7 $X2=0.69 $Y2=2.7
cc_197 N_A_c_240_n N_Y_c_462_n 5.06602e-19 $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.7
cc_198 N_A_c_255_n N_Y_c_462_n 0.0226156f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.7
cc_199 N_A_c_257_n N_Y_c_462_n 0.00165526f $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.7
cc_200 A N_Y_c_462_n 0.00938699f $X=0.32 $Y=3.065 $X2=0.69 $Y2=2.7
cc_201 N_A_c_202_n N_Y_c_426_n 0.00265306f $X=1.335 $Y=1.44 $X2=1.55 $Y2=0.865
cc_202 N_A_c_206_n N_Y_c_426_n 0.00317228f $X=1.69 $Y=1.515 $X2=1.55 $Y2=0.865
cc_203 N_A_c_208_n N_Y_c_426_n 0.00265306f $X=1.765 $Y=1.44 $X2=1.55 $Y2=0.865
cc_204 N_A_c_269_n N_Y_c_465_n 0.00360548f $X=1.335 $Y=2.7 $X2=1.55 $Y2=2.7
cc_205 N_A_c_207_n N_Y_c_465_n 0.0108863f $X=1.69 $Y=2.625 $X2=1.55 $Y2=2.7
cc_206 N_A_c_274_n N_Y_c_465_n 0.00360548f $X=1.765 $Y=2.7 $X2=1.55 $Y2=2.7
cc_207 N_A_c_215_n N_Y_c_431_n 0.00265306f $X=2.195 $Y=1.44 $X2=2.41 $Y2=0.865
cc_208 N_A_c_220_n N_Y_c_431_n 0.00317228f $X=2.55 $Y=1.515 $X2=2.41 $Y2=0.865
cc_209 N_A_c_222_n N_Y_c_431_n 0.00265306f $X=2.625 $Y=1.44 $X2=2.41 $Y2=0.865
cc_210 N_A_c_280_n N_Y_c_468_n 0.00360548f $X=2.195 $Y=2.7 $X2=2.41 $Y2=2.7
cc_211 N_A_c_221_n N_Y_c_468_n 0.0108863f $X=2.55 $Y=2.625 $X2=2.41 $Y2=2.7
cc_212 N_A_c_285_n N_Y_c_468_n 0.00360548f $X=2.625 $Y=2.7 $X2=2.41 $Y2=2.7
cc_213 N_A_c_229_n N_Y_c_436_n 0.00265306f $X=3.055 $Y=1.44 $X2=3.27 $Y2=0.865
cc_214 N_A_c_233_n N_Y_c_436_n 0.00317228f $X=3.41 $Y=1.515 $X2=3.27 $Y2=0.865
cc_215 N_A_c_235_n N_Y_c_436_n 0.00265306f $X=3.485 $Y=1.44 $X2=3.27 $Y2=0.865
cc_216 N_A_c_291_n N_Y_c_471_n 0.00360548f $X=3.055 $Y=2.7 $X2=3.27 $Y2=2.7
cc_217 N_A_c_234_n N_Y_c_471_n 0.0105836f $X=3.41 $Y=2.625 $X2=3.27 $Y2=2.7
cc_218 N_A_c_296_n N_Y_c_471_n 0.00360548f $X=3.485 $Y=2.7 $X2=3.27 $Y2=2.7
cc_219 N_A_c_188_n N_Y_c_440_n 0.00942005f $X=0.475 $Y=1.44 $X2=0.69 $Y2=1.335
cc_220 N_A_c_195_n N_Y_c_440_n 0.00259753f $X=0.905 $Y=1.44 $X2=0.69 $Y2=1.335
cc_221 N_A_c_240_n N_Y_c_440_n 0.0011424f $X=0.535 $Y=2.045 $X2=0.69 $Y2=1.335
cc_222 N_A_c_258_n N_Y_c_474_n 0.00169643f $X=0.475 $Y=2.7 $X2=0.69 $Y2=2.585
cc_223 N_A_c_194_n N_Y_c_474_n 0.00270155f $X=0.83 $Y=2.625 $X2=0.69 $Y2=2.585
cc_224 N_A_c_263_n N_Y_c_474_n 0.00144225f $X=0.905 $Y=2.7 $X2=0.69 $Y2=2.585
cc_225 N_A_c_240_n N_Y_c_474_n 8.31386e-19 $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.585
cc_226 N_A_c_242_n N_Y_c_474_n 0.00102602f $X=0.475 $Y=2.625 $X2=0.69 $Y2=2.585
cc_227 N_A_c_244_n N_Y_c_474_n 0.00150284f $X=0.905 $Y=2.625 $X2=0.69 $Y2=2.585
cc_228 N_A_c_255_n N_Y_c_474_n 0.0071561f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.585
cc_229 N_A_c_257_n N_Y_c_474_n 0.00173027f $X=0.535 $Y=2.045 $X2=0.69 $Y2=2.585
cc_230 A N_Y_c_474_n 0.00815006f $X=0.32 $Y=3.065 $X2=0.69 $Y2=2.585
cc_231 N_A_c_188_n Y 0.00150089f $X=0.475 $Y=1.44 $X2=0.76 $Y2=1.94
cc_232 N_A_c_192_n Y 0.00792324f $X=0.475 $Y=2.55 $X2=0.76 $Y2=1.94
cc_233 N_A_c_193_n Y 0.0161013f $X=0.83 $Y=1.515 $X2=0.76 $Y2=1.94
cc_234 N_A_c_194_n Y 0.00363305f $X=0.83 $Y=2.625 $X2=0.76 $Y2=1.94
cc_235 N_A_c_195_n Y 0.00150089f $X=0.905 $Y=1.44 $X2=0.76 $Y2=1.94
cc_236 N_A_c_240_n Y 0.00668675f $X=0.535 $Y=2.045 $X2=0.76 $Y2=1.94
cc_237 N_A_c_241_n Y 0.00675469f $X=0.535 $Y=1.88 $X2=0.76 $Y2=1.94
cc_238 N_A_c_255_n Y 0.0182346f $X=0.32 $Y=3.07 $X2=0.76 $Y2=1.94
cc_239 N_A_c_257_n Y 0.0178517f $X=0.535 $Y=2.045 $X2=0.76 $Y2=1.94
cc_240 N_A_c_195_n N_Y_c_444_n 0.0129682f $X=0.905 $Y=1.44 $X2=1.405 $Y2=1.22
cc_241 N_A_c_199_n N_Y_c_444_n 0.0022289f $X=1.26 $Y=1.515 $X2=1.405 $Y2=1.22
cc_242 N_A_c_202_n N_Y_c_444_n 0.0129682f $X=1.335 $Y=1.44 $X2=1.405 $Y2=1.22
cc_243 N_A_c_263_n N_Y_c_475_n 0.00693713f $X=0.905 $Y=2.7 $X2=1.405 $Y2=2.7
cc_244 N_A_c_201_n N_Y_c_475_n 0.0120397f $X=1.26 $Y=2.625 $X2=1.405 $Y2=2.7
cc_245 N_A_c_269_n N_Y_c_475_n 0.00693713f $X=1.335 $Y=2.7 $X2=1.405 $Y2=2.7
cc_246 N_A_c_244_n N_Y_c_475_n 0.00560085f $X=0.905 $Y=2.625 $X2=1.405 $Y2=2.7
cc_247 N_A_c_246_n N_Y_c_475_n 0.00560085f $X=1.335 $Y=2.625 $X2=1.405 $Y2=2.7
cc_248 N_A_c_202_n N_Y_c_446_n 0.00150089f $X=1.335 $Y=1.44 $X2=1.55 $Y2=2.585
cc_249 N_A_c_206_n N_Y_c_446_n 0.0177499f $X=1.69 $Y=1.515 $X2=1.55 $Y2=2.585
cc_250 N_A_c_207_n N_Y_c_446_n 0.00562481f $X=1.69 $Y=2.625 $X2=1.55 $Y2=2.585
cc_251 N_A_c_208_n N_Y_c_446_n 0.00150089f $X=1.765 $Y=1.44 $X2=1.55 $Y2=2.585
cc_252 N_A_c_219_n N_Y_c_446_n 0.0141566f $X=2.195 $Y=2.55 $X2=1.55 $Y2=2.585
cc_253 N_A_c_208_n N_Y_c_447_n 0.0129682f $X=1.765 $Y=1.44 $X2=2.265 $Y2=1.22
cc_254 N_A_c_212_n N_Y_c_447_n 0.0022289f $X=2.12 $Y=1.515 $X2=2.265 $Y2=1.22
cc_255 N_A_c_215_n N_Y_c_447_n 0.0136594f $X=2.195 $Y=1.44 $X2=2.265 $Y2=1.22
cc_256 N_A_c_202_n N_Y_c_449_n 0.00259753f $X=1.335 $Y=1.44 $X2=1.695 $Y2=1.22
cc_257 N_A_c_208_n N_Y_c_449_n 0.00259753f $X=1.765 $Y=1.44 $X2=1.695 $Y2=1.22
cc_258 N_A_c_274_n N_Y_c_477_n 0.00693713f $X=1.765 $Y=2.7 $X2=2.265 $Y2=2.7
cc_259 N_A_c_214_n N_Y_c_477_n 0.0125508f $X=2.12 $Y=2.625 $X2=2.265 $Y2=2.7
cc_260 N_A_c_280_n N_Y_c_477_n 0.00693713f $X=2.195 $Y=2.7 $X2=2.265 $Y2=2.7
cc_261 N_A_c_248_n N_Y_c_477_n 0.00560085f $X=1.765 $Y=2.625 $X2=2.265 $Y2=2.7
cc_262 N_A_c_250_n N_Y_c_477_n 0.00642784f $X=2.195 $Y=2.625 $X2=2.265 $Y2=2.7
cc_263 N_A_c_269_n N_Y_c_479_n 0.00144225f $X=1.335 $Y=2.7 $X2=1.695 $Y2=2.7
cc_264 N_A_c_207_n N_Y_c_479_n 0.00397642f $X=1.69 $Y=2.625 $X2=1.695 $Y2=2.7
cc_265 N_A_c_274_n N_Y_c_479_n 0.00144225f $X=1.765 $Y=2.7 $X2=1.695 $Y2=2.7
cc_266 N_A_c_246_n N_Y_c_479_n 0.00150284f $X=1.335 $Y=2.625 $X2=1.695 $Y2=2.7
cc_267 N_A_c_248_n N_Y_c_479_n 0.00150284f $X=1.765 $Y=2.625 $X2=1.695 $Y2=2.7
cc_268 N_A_c_215_n N_Y_c_452_n 0.00150089f $X=2.195 $Y=1.44 $X2=2.41 $Y2=2.585
cc_269 N_A_c_219_n N_Y_c_452_n 0.0182294f $X=2.195 $Y=2.55 $X2=2.41 $Y2=2.585
cc_270 N_A_c_220_n N_Y_c_452_n 0.0177499f $X=2.55 $Y=1.515 $X2=2.41 $Y2=2.585
cc_271 N_A_c_221_n N_Y_c_452_n 0.00562481f $X=2.55 $Y=2.625 $X2=2.41 $Y2=2.585
cc_272 N_A_c_222_n N_Y_c_452_n 0.00150089f $X=2.625 $Y=1.44 $X2=2.41 $Y2=2.585
cc_273 N_A_c_222_n N_Y_c_453_n 0.0129682f $X=2.625 $Y=1.44 $X2=3.125 $Y2=1.22
cc_274 N_A_c_226_n N_Y_c_453_n 0.0022289f $X=2.98 $Y=1.515 $X2=3.125 $Y2=1.22
cc_275 N_A_c_229_n N_Y_c_453_n 0.0129682f $X=3.055 $Y=1.44 $X2=3.125 $Y2=1.22
cc_276 N_A_c_215_n N_Y_c_455_n 0.00262362f $X=2.195 $Y=1.44 $X2=2.555 $Y2=1.22
cc_277 N_A_c_222_n N_Y_c_455_n 0.00259753f $X=2.625 $Y=1.44 $X2=2.555 $Y2=1.22
cc_278 N_A_c_285_n N_Y_c_480_n 0.00693713f $X=2.625 $Y=2.7 $X2=3.125 $Y2=2.7
cc_279 N_A_c_228_n N_Y_c_480_n 0.0120397f $X=2.98 $Y=2.625 $X2=3.125 $Y2=2.7
cc_280 N_A_c_291_n N_Y_c_480_n 0.00693713f $X=3.055 $Y=2.7 $X2=3.125 $Y2=2.7
cc_281 N_A_c_252_n N_Y_c_480_n 0.00560085f $X=2.625 $Y=2.625 $X2=3.125 $Y2=2.7
cc_282 N_A_c_254_n N_Y_c_480_n 0.00560085f $X=3.055 $Y=2.625 $X2=3.125 $Y2=2.7
cc_283 N_A_c_280_n N_Y_c_482_n 0.00144225f $X=2.195 $Y=2.7 $X2=2.555 $Y2=2.7
cc_284 N_A_c_221_n N_Y_c_482_n 0.00397642f $X=2.55 $Y=2.625 $X2=2.555 $Y2=2.7
cc_285 N_A_c_285_n N_Y_c_482_n 0.00144225f $X=2.625 $Y=2.7 $X2=2.555 $Y2=2.7
cc_286 N_A_c_250_n N_Y_c_482_n 0.00153387f $X=2.195 $Y=2.625 $X2=2.555 $Y2=2.7
cc_287 N_A_c_252_n N_Y_c_482_n 0.00150284f $X=2.625 $Y=2.625 $X2=2.555 $Y2=2.7
cc_288 N_A_c_229_n N_Y_c_458_n 0.00259753f $X=3.055 $Y=1.44 $X2=3.27 $Y2=1.335
cc_289 N_A_c_235_n N_Y_c_458_n 0.00939395f $X=3.485 $Y=1.44 $X2=3.27 $Y2=1.335
cc_290 N_A_c_229_n N_Y_c_461_n 0.00150089f $X=3.055 $Y=1.44 $X2=3.27 $Y2=2.585
cc_291 N_A_c_291_n N_Y_c_461_n 0.00144225f $X=3.055 $Y=2.7 $X2=3.27 $Y2=2.585
cc_292 N_A_c_233_n N_Y_c_461_n 0.0169795f $X=3.41 $Y=1.515 $X2=3.27 $Y2=2.585
cc_293 N_A_c_234_n N_Y_c_461_n 0.0141541f $X=3.41 $Y=2.625 $X2=3.27 $Y2=2.585
cc_294 N_A_c_235_n N_Y_c_461_n 0.00150089f $X=3.485 $Y=1.44 $X2=3.27 $Y2=2.585
cc_295 N_A_c_296_n N_Y_c_461_n 0.00541616f $X=3.485 $Y=2.7 $X2=3.27 $Y2=2.585
cc_296 N_A_c_254_n N_Y_c_461_n 0.00150284f $X=3.055 $Y=2.625 $X2=3.27 $Y2=2.585
