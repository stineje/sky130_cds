* File: sky130_osu_sc_15T_ls__buf_4.pex.spice
* Created: Fri Nov 12 14:54:58 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__BUF_4%GND 1 2 3 31 35 39 41 42 49 63 65
r57 63 65 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r58 47 49 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.865
r59 41 47 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.325 $Y=0.152
+ $X2=2.41 $Y2=0.305
r60 37 42 3.38889 $w=3.06e-07 $l=8.6487e-08 $layer=LI1_cond $X=1.55 $Y=0.155
+ $X2=1.635 $Y2=0.152
r61 37 39 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.865
r62 33 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.865
r63 31 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r64 31 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r65 31 37 21.1307 $w=3.06e-07 $l=5.3e-07 $layer=LI1_cond $X=1.02 $Y=0.155
+ $X2=1.55 $Y2=0.155
r66 31 33 13.1569 $w=3.06e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=0.155
+ $X2=0.69 $Y2=0.155
r67 31 33 13.9542 $w=3.06e-07 $l=3.5e-07 $layer=LI1_cond $X=0.34 $Y=0.155
+ $X2=0.69 $Y2=0.155
r68 31 41 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r69 31 42 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r70 3 49 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.865
r71 2 39 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.865
r72 1 35 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_4%VDD 1 2 3 25 27 34 38 44 48 55 62 66
r44 62 66 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.7 $Y2=5.397
r45 55 58 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.205
+ $X2=2.41 $Y2=4.565
r46 53 58 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=5.245
+ $X2=2.41 $Y2=4.565
r47 51 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=5.36 $X2=1.7
+ $Y2=5.36
r48 49 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=5.397
+ $X2=1.55 $Y2=5.397
r49 49 51 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=5.397
+ $X2=1.7 $Y2=5.397
r50 48 53 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.325 $Y=5.397
+ $X2=2.41 $Y2=5.245
r51 48 51 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=5.397
+ $X2=1.7 $Y2=5.397
r52 44 47 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.205
+ $X2=1.55 $Y2=4.565
r53 42 60 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=5.245
+ $X2=1.55 $Y2=5.397
r54 42 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=5.245
+ $X2=1.55 $Y2=4.565
r55 39 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r56 39 41 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r57 38 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=5.397
+ $X2=1.55 $Y2=5.397
r58 38 41 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=5.397
+ $X2=1.02 $Y2=5.397
r59 34 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=3.885
+ $X2=0.69 $Y2=4.565
r60 32 59 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r61 32 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r62 29 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r63 27 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r64 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r65 25 51 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r66 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r67 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r68 3 58 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.565
r69 3 55 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.205
r70 2 47 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.565
r71 2 44 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.205
r72 1 37 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r73 1 34 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_4%A 3 7 10 14 20
r39 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.07
+ $X2=0.635 $Y2=3.07
r40 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2.22
+ $X2=0.635 $Y2=3.07
r41 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.22 $X2=0.635 $Y2=2.22
r42 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.22
+ $X2=0.585 $Y2=2.385
r43 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.22
+ $X2=0.585 $Y2=2.055
r44 7 12 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.385
r45 3 11 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_4%A_27_115# 1 3 11 13 15 17 20 22 24 25 26
+ 27 28 31 33 35 36 38 42 44 46 56 57 60 64 68 70 73
c118 33 0 1.33323e-19 $X=1.765 $Y=2.75
c119 31 0 1.33323e-19 $X=1.765 $Y=0.945
c120 22 0 1.33323e-19 $X=1.335 $Y=2.75
c121 20 0 1.33323e-19 $X=1.335 $Y=0.945
r122 69 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.675
+ $X2=0.26 $Y2=1.675
r123 68 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.675
+ $X2=0.965 $Y2=1.675
r124 68 69 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.675
+ $X2=0.345 $Y2=1.675
r125 64 66 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r126 62 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.76
+ $X2=0.26 $Y2=1.675
r127 62 64 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=0.26 $Y=1.76
+ $X2=0.26 $Y2=3.205
r128 58 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=1.675
r129 58 60 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.865
r130 53 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.675 $X2=0.965 $Y2=1.675
r131 53 54 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=1.18 $Y2=1.675
r132 51 53 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.965 $Y2=1.675
r133 49 50 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.675
+ $X2=1.335 $Y2=2.675
r134 47 49 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.675
+ $X2=1.18 $Y2=2.675
r135 44 46 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.195 $Y=2.75
+ $X2=2.195 $Y2=3.825
r136 40 42 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=0.945
r137 39 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.675
+ $X2=1.765 $Y2=2.675
r138 38 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=2.675
+ $X2=2.195 $Y2=2.75
r139 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.675
+ $X2=1.84 $Y2=2.675
r140 37 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.585
+ $X2=1.765 $Y2=1.585
r141 36 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=2.195 $Y2=1.51
r142 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=1.84 $Y2=1.585
r143 33 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.75
+ $X2=1.765 $Y2=2.675
r144 33 35 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.765 $Y=2.75
+ $X2=1.765 $Y2=3.825
r145 29 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=1.585
r146 29 31 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=0.945
r147 28 50 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.675
+ $X2=1.335 $Y2=2.675
r148 27 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.675
+ $X2=1.765 $Y2=2.675
r149 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.675
+ $X2=1.41 $Y2=2.675
r150 25 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.585
+ $X2=1.765 $Y2=1.585
r151 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.585
+ $X2=1.41 $Y2=1.585
r152 22 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.75
+ $X2=1.335 $Y2=2.675
r153 22 24 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.335 $Y=2.75
+ $X2=1.335 $Y2=3.825
r154 18 26 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.41 $Y2=1.585
r155 18 54 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.18 $Y2=1.675
r156 18 20 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.945
r157 17 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.6
+ $X2=1.18 $Y2=2.675
r158 16 54 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.84
+ $X2=1.18 $Y2=1.675
r159 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.84
+ $X2=1.18 $Y2=2.6
r160 13 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=2.675
r161 13 15 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=3.825
r162 9 51 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.905 $Y2=1.675
r163 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.905 $Y2=0.945
r164 3 66 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r165 3 64 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r166 1 60 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__BUF_4%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c80 55 0 1.33323e-19 $X=1.98 $Y=2.585
c81 54 0 1.33323e-19 $X=1.98 $Y=1.335
c82 46 0 1.33323e-19 $X=1.12 $Y=2.585
c83 45 0 1.33323e-19 $X=1.12 $Y=1.335
r84 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.585
+ $X2=1.98 $Y2=2.7
r85 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.335
+ $X2=1.98 $Y2=1.22
r86 54 55 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.335
+ $X2=1.98 $Y2=2.585
r87 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.7
+ $X2=1.12 $Y2=2.7
r88 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.7
+ $X2=1.98 $Y2=2.7
r89 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.7
+ $X2=1.265 $Y2=2.7
r90 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1.22
+ $X2=1.12 $Y2=1.22
r91 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1.22
+ $X2=1.98 $Y2=1.22
r92 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1.22
+ $X2=1.265 $Y2=1.22
r93 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.585
+ $X2=1.12 $Y2=2.7
r94 46 48 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.585
+ $X2=1.12 $Y2=2.01
r95 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=1.22
r96 45 48 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=2.01
r97 41 43 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.205
+ $X2=1.98 $Y2=4.565
r98 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.7 $X2=1.98
+ $Y2=2.7
r99 38 41 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.98 $Y=2.7
+ $X2=1.98 $Y2=3.205
r100 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1.22
+ $X2=1.98 $Y2=1.22
r101 32 35 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.98 $Y=0.865
+ $X2=1.98 $Y2=1.22
r102 27 29 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=3.205
+ $X2=1.12 $Y2=4.565
r103 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.7
+ $X2=1.12 $Y2=2.7
r104 24 27 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.12 $Y=2.7
+ $X2=1.12 $Y2=3.205
r105 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.22
+ $X2=1.12 $Y2=1.22
r106 18 21 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.12 $Y=0.865
+ $X2=1.12 $Y2=1.22
r107 6 43 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.565
r108 6 41 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.205
r109 5 29 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r110 5 27 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.205
r111 2 32 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.865
r112 1 18 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
.ends

