* File: sky130_osu_sc_18T_ms__inv_10.pxi.spice
* Created: Fri Nov 12 14:03:57 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__INV_10%GND N_GND_M1000_d N_GND_M1002_d N_GND_M1005_d
+ N_GND_M1010_d N_GND_M1014_d N_GND_M1018_d N_GND_M1000_b N_GND_c_2_p
+ N_GND_c_3_p N_GND_c_10_p N_GND_c_17_p N_GND_c_23_p N_GND_c_30_p N_GND_c_37_p
+ N_GND_c_44_p N_GND_c_50_p N_GND_c_57_p N_GND_c_63_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_MS__INV_10%GND
x_PM_SKY130_OSU_SC_18T_MS__INV_10%VDD N_VDD_M1001_d N_VDD_M1003_d N_VDD_M1007_d
+ N_VDD_M1011_d N_VDD_M1015_d N_VDD_M1019_d N_VDD_M1001_b N_VDD_c_140_p
+ N_VDD_c_141_p N_VDD_c_146_p N_VDD_c_152_p N_VDD_c_157_p N_VDD_c_163_p
+ N_VDD_c_168_p N_VDD_c_174_p N_VDD_c_179_p N_VDD_c_185_p N_VDD_c_190_p VDD
+ N_VDD_c_142_p PM_SKY130_OSU_SC_18T_MS__INV_10%VDD
x_PM_SKY130_OSU_SC_18T_MS__INV_10%A N_A_c_235_n N_A_M1000_g N_A_c_239_n
+ N_A_c_322_n N_A_M1001_g N_A_c_240_n N_A_c_241_n N_A_c_242_n N_A_M1002_g
+ N_A_c_327_n N_A_M1003_g N_A_c_246_n N_A_c_248_n N_A_c_249_n N_A_M1004_g
+ N_A_c_333_n N_A_M1006_g N_A_c_253_n N_A_c_254_n N_A_c_255_n N_A_M1005_g
+ N_A_c_338_n N_A_M1007_g N_A_c_259_n N_A_c_261_n N_A_c_262_n N_A_M1008_g
+ N_A_c_266_n N_A_c_344_n N_A_M1009_g N_A_c_267_n N_A_c_268_n N_A_c_269_n
+ N_A_M1010_g N_A_c_349_n N_A_M1011_g N_A_c_273_n N_A_c_275_n N_A_c_276_n
+ N_A_M1012_g N_A_c_355_n N_A_M1013_g N_A_c_280_n N_A_c_281_n N_A_c_282_n
+ N_A_M1014_g N_A_c_360_n N_A_M1015_g N_A_c_286_n N_A_c_288_n N_A_c_289_n
+ N_A_M1016_g N_A_c_366_n N_A_M1017_g N_A_c_293_n N_A_c_294_n N_A_c_295_n
+ N_A_M1018_g N_A_c_371_n N_A_M1019_g N_A_c_299_n N_A_c_300_n N_A_c_301_n
+ N_A_c_302_n N_A_c_303_n N_A_c_304_n N_A_c_305_n N_A_c_306_n N_A_c_307_n
+ N_A_c_308_n N_A_c_309_n N_A_c_310_n N_A_c_311_n N_A_c_312_n N_A_c_313_n
+ N_A_c_314_n N_A_c_315_n N_A_c_316_n N_A_c_317_n N_A_c_318_n N_A_c_319_n
+ N_A_c_320_n N_A_c_321_n A PM_SKY130_OSU_SC_18T_MS__INV_10%A
x_PM_SKY130_OSU_SC_18T_MS__INV_10%Y N_Y_M1000_s N_Y_M1004_s N_Y_M1008_s
+ N_Y_M1012_s N_Y_M1016_s N_Y_M1001_s N_Y_M1006_s N_Y_M1009_s N_Y_M1013_s
+ N_Y_M1017_s N_Y_c_524_n N_Y_c_575_n N_Y_c_528_n N_Y_c_578_n N_Y_c_533_n
+ N_Y_c_581_n N_Y_c_538_n N_Y_c_584_n N_Y_c_543_n N_Y_c_587_n N_Y_c_547_n
+ N_Y_c_590_n Y N_Y_c_551_n N_Y_c_591_n N_Y_c_553_n N_Y_c_554_n N_Y_c_556_n
+ N_Y_c_593_n N_Y_c_595_n N_Y_c_559_n N_Y_c_560_n N_Y_c_562_n N_Y_c_596_n
+ N_Y_c_598_n N_Y_c_565_n N_Y_c_566_n N_Y_c_568_n N_Y_c_599_n N_Y_c_601_n
+ N_Y_c_571_n N_Y_c_574_n PM_SKY130_OSU_SC_18T_MS__INV_10%Y
cc_1 N_GND_M1000_b N_A_c_235_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.7
cc_2 N_GND_c_2_p N_A_c_235_n 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.7
cc_3 N_GND_c_3_p N_A_c_235_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.7
cc_4 N_GND_c_4_p N_A_c_235_n 0.00468827f $X=4.42 $Y=0.19 $X2=0.475 $Y2=1.7
cc_5 N_GND_M1000_b N_A_c_239_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.81
cc_6 N_GND_M1000_b N_A_c_240_n 0.01476f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.775
cc_7 N_GND_M1000_b N_A_c_241_n 0.00981662f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.885
cc_8 N_GND_M1000_b N_A_c_242_n 0.0166526f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.7
cc_9 N_GND_c_3_p N_A_c_242_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.7
cc_10 N_GND_c_10_p N_A_c_242_n 0.00356864f $X=1.12 $Y=0.825 $X2=0.905 $Y2=1.7
cc_11 N_GND_c_4_p N_A_c_242_n 0.00468827f $X=4.42 $Y=0.19 $X2=0.905 $Y2=1.7
cc_12 N_GND_M1000_b N_A_c_246_n 0.0213783f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.775
cc_13 N_GND_c_10_p N_A_c_246_n 0.00283047f $X=1.12 $Y=0.825 $X2=1.26 $Y2=1.775
cc_14 N_GND_M1000_b N_A_c_248_n 0.0173499f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.885
cc_15 N_GND_M1000_b N_A_c_249_n 0.0166526f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.7
cc_16 N_GND_c_10_p N_A_c_249_n 0.00356864f $X=1.12 $Y=0.825 $X2=1.335 $Y2=1.7
cc_17 N_GND_c_17_p N_A_c_249_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.335 $Y2=1.7
cc_18 N_GND_c_4_p N_A_c_249_n 0.00468827f $X=4.42 $Y=0.19 $X2=1.335 $Y2=1.7
cc_19 N_GND_M1000_b N_A_c_253_n 0.0195339f $X=-0.045 $Y=0 $X2=1.69 $Y2=1.775
cc_20 N_GND_M1000_b N_A_c_254_n 0.0145324f $X=-0.045 $Y=0 $X2=1.69 $Y2=2.885
cc_21 N_GND_M1000_b N_A_c_255_n 0.0166526f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.7
cc_22 N_GND_c_17_p N_A_c_255_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.765 $Y2=1.7
cc_23 N_GND_c_23_p N_A_c_255_n 0.00356864f $X=1.98 $Y=0.825 $X2=1.765 $Y2=1.7
cc_24 N_GND_c_4_p N_A_c_255_n 0.00468827f $X=4.42 $Y=0.19 $X2=1.765 $Y2=1.7
cc_25 N_GND_M1000_b N_A_c_259_n 0.0164591f $X=-0.045 $Y=0 $X2=2.12 $Y2=1.775
cc_26 N_GND_c_23_p N_A_c_259_n 0.00283047f $X=1.98 $Y=0.825 $X2=2.12 $Y2=1.775
cc_27 N_GND_M1000_b N_A_c_261_n 0.0124307f $X=-0.045 $Y=0 $X2=2.12 $Y2=2.885
cc_28 N_GND_M1000_b N_A_c_262_n 0.0166526f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.7
cc_29 N_GND_c_23_p N_A_c_262_n 0.00356864f $X=1.98 $Y=0.825 $X2=2.195 $Y2=1.7
cc_30 N_GND_c_30_p N_A_c_262_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.195 $Y2=1.7
cc_31 N_GND_c_4_p N_A_c_262_n 0.00468827f $X=4.42 $Y=0.19 $X2=2.195 $Y2=1.7
cc_32 N_GND_M1000_b N_A_c_266_n 0.0685082f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.81
cc_33 N_GND_M1000_b N_A_c_267_n 0.0195339f $X=-0.045 $Y=0 $X2=2.55 $Y2=1.775
cc_34 N_GND_M1000_b N_A_c_268_n 0.0145324f $X=-0.045 $Y=0 $X2=2.55 $Y2=2.885
cc_35 N_GND_M1000_b N_A_c_269_n 0.0166526f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.7
cc_36 N_GND_c_30_p N_A_c_269_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.625 $Y2=1.7
cc_37 N_GND_c_37_p N_A_c_269_n 0.00356864f $X=2.84 $Y=0.825 $X2=2.625 $Y2=1.7
cc_38 N_GND_c_4_p N_A_c_269_n 0.00468827f $X=4.42 $Y=0.19 $X2=2.625 $Y2=1.7
cc_39 N_GND_M1000_b N_A_c_273_n 0.0213783f $X=-0.045 $Y=0 $X2=2.98 $Y2=1.775
cc_40 N_GND_c_37_p N_A_c_273_n 0.00283047f $X=2.84 $Y=0.825 $X2=2.98 $Y2=1.775
cc_41 N_GND_M1000_b N_A_c_275_n 0.0173499f $X=-0.045 $Y=0 $X2=2.98 $Y2=2.885
cc_42 N_GND_M1000_b N_A_c_276_n 0.0166526f $X=-0.045 $Y=0 $X2=3.055 $Y2=1.7
cc_43 N_GND_c_37_p N_A_c_276_n 0.00356864f $X=2.84 $Y=0.825 $X2=3.055 $Y2=1.7
cc_44 N_GND_c_44_p N_A_c_276_n 0.00606474f $X=3.615 $Y=0.152 $X2=3.055 $Y2=1.7
cc_45 N_GND_c_4_p N_A_c_276_n 0.00468827f $X=4.42 $Y=0.19 $X2=3.055 $Y2=1.7
cc_46 N_GND_M1000_b N_A_c_280_n 0.0195339f $X=-0.045 $Y=0 $X2=3.41 $Y2=1.775
cc_47 N_GND_M1000_b N_A_c_281_n 0.0145324f $X=-0.045 $Y=0 $X2=3.41 $Y2=2.885
cc_48 N_GND_M1000_b N_A_c_282_n 0.0166526f $X=-0.045 $Y=0 $X2=3.485 $Y2=1.7
cc_49 N_GND_c_44_p N_A_c_282_n 0.00606474f $X=3.615 $Y=0.152 $X2=3.485 $Y2=1.7
cc_50 N_GND_c_50_p N_A_c_282_n 0.00356864f $X=3.7 $Y=0.825 $X2=3.485 $Y2=1.7
cc_51 N_GND_c_4_p N_A_c_282_n 0.00468827f $X=4.42 $Y=0.19 $X2=3.485 $Y2=1.7
cc_52 N_GND_M1000_b N_A_c_286_n 0.0213783f $X=-0.045 $Y=0 $X2=3.84 $Y2=1.775
cc_53 N_GND_c_50_p N_A_c_286_n 0.00283047f $X=3.7 $Y=0.825 $X2=3.84 $Y2=1.775
cc_54 N_GND_M1000_b N_A_c_288_n 0.0173499f $X=-0.045 $Y=0 $X2=3.84 $Y2=2.885
cc_55 N_GND_M1000_b N_A_c_289_n 0.0166526f $X=-0.045 $Y=0 $X2=3.915 $Y2=1.7
cc_56 N_GND_c_50_p N_A_c_289_n 0.00356864f $X=3.7 $Y=0.825 $X2=3.915 $Y2=1.7
cc_57 N_GND_c_57_p N_A_c_289_n 0.00606474f $X=4.475 $Y=0.152 $X2=3.915 $Y2=1.7
cc_58 N_GND_c_4_p N_A_c_289_n 0.00468827f $X=4.42 $Y=0.19 $X2=3.915 $Y2=1.7
cc_59 N_GND_M1000_b N_A_c_293_n 0.0385034f $X=-0.045 $Y=0 $X2=4.27 $Y2=1.775
cc_60 N_GND_M1000_b N_A_c_294_n 0.0295863f $X=-0.045 $Y=0 $X2=4.27 $Y2=2.885
cc_61 N_GND_M1000_b N_A_c_295_n 0.0208613f $X=-0.045 $Y=0 $X2=4.345 $Y2=1.7
cc_62 N_GND_c_57_p N_A_c_295_n 0.00606474f $X=4.475 $Y=0.152 $X2=4.345 $Y2=1.7
cc_63 N_GND_c_63_p N_A_c_295_n 0.00713292f $X=4.56 $Y=0.825 $X2=4.345 $Y2=1.7
cc_64 N_GND_c_4_p N_A_c_295_n 0.00468827f $X=4.42 $Y=0.19 $X2=4.345 $Y2=1.7
cc_65 N_GND_M1000_b N_A_c_299_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.775
cc_66 N_GND_M1000_b N_A_c_300_n 0.0382476f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_67 N_GND_M1000_b N_A_c_301_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.14
cc_68 N_GND_M1000_b N_A_c_302_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.885
cc_69 N_GND_M1000_b N_A_c_303_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.775
cc_70 N_GND_M1000_b N_A_c_304_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.885
cc_71 N_GND_M1000_b N_A_c_305_n 0.0106787f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.775
cc_72 N_GND_M1000_b N_A_c_306_n 0.00980309f $X=-0.045 $Y=0 $X2=1.335 $Y2=2.885
cc_73 N_GND_M1000_b N_A_c_307_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.775
cc_74 N_GND_M1000_b N_A_c_308_n 0.00980309f $X=-0.045 $Y=0 $X2=1.765 $Y2=2.885
cc_75 N_GND_M1000_b N_A_c_309_n 0.0023879f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.775
cc_76 N_GND_M1000_b N_A_c_310_n 0.00151234f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.885
cc_77 N_GND_M1000_b N_A_c_311_n 0.0106787f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.775
cc_78 N_GND_M1000_b N_A_c_312_n 0.00980309f $X=-0.045 $Y=0 $X2=2.625 $Y2=2.885
cc_79 N_GND_M1000_b N_A_c_313_n 0.0106787f $X=-0.045 $Y=0 $X2=3.055 $Y2=1.775
cc_80 N_GND_M1000_b N_A_c_314_n 0.00980309f $X=-0.045 $Y=0 $X2=3.055 $Y2=2.885
cc_81 N_GND_M1000_b N_A_c_315_n 0.0106787f $X=-0.045 $Y=0 $X2=3.485 $Y2=1.775
cc_82 N_GND_M1000_b N_A_c_316_n 0.00980309f $X=-0.045 $Y=0 $X2=3.485 $Y2=2.885
cc_83 N_GND_M1000_b N_A_c_317_n 0.0106787f $X=-0.045 $Y=0 $X2=3.915 $Y2=1.775
cc_84 N_GND_M1000_b N_A_c_318_n 0.00980309f $X=-0.045 $Y=0 $X2=3.915 $Y2=2.885
cc_85 N_GND_M1000_b N_A_c_319_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.33
cc_86 N_GND_M1000_b N_A_c_320_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.305
cc_87 N_GND_M1000_b N_A_c_321_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_88 N_GND_M1000_b N_Y_c_524_n 0.00155118f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_89 N_GND_c_3_p N_Y_c_524_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.825
cc_90 N_GND_c_10_p N_Y_c_524_n 8.14297e-19 $X=1.12 $Y=0.825 $X2=0.69 $Y2=0.825
cc_91 N_GND_c_4_p N_Y_c_524_n 0.00475776f $X=4.42 $Y=0.19 $X2=0.69 $Y2=0.825
cc_92 N_GND_M1000_b N_Y_c_528_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_93 N_GND_c_10_p N_Y_c_528_n 8.14297e-19 $X=1.12 $Y=0.825 $X2=1.55 $Y2=0.825
cc_94 N_GND_c_17_p N_Y_c_528_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.825
cc_95 N_GND_c_23_p N_Y_c_528_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=0.825
cc_96 N_GND_c_4_p N_Y_c_528_n 0.00475776f $X=4.42 $Y=0.19 $X2=1.55 $Y2=0.825
cc_97 N_GND_M1000_b N_Y_c_533_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.825
cc_98 N_GND_c_23_p N_Y_c_533_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=0.825
cc_99 N_GND_c_30_p N_Y_c_533_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.825
cc_100 N_GND_c_37_p N_Y_c_533_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=2.41 $Y2=0.825
cc_101 N_GND_c_4_p N_Y_c_533_n 0.00475776f $X=4.42 $Y=0.19 $X2=2.41 $Y2=0.825
cc_102 N_GND_M1000_b N_Y_c_538_n 0.00155118f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.825
cc_103 N_GND_c_37_p N_Y_c_538_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=3.27 $Y2=0.825
cc_104 N_GND_c_44_p N_Y_c_538_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.825
cc_105 N_GND_c_50_p N_Y_c_538_n 8.14297e-19 $X=3.7 $Y=0.825 $X2=3.27 $Y2=0.825
cc_106 N_GND_c_4_p N_Y_c_538_n 0.00475776f $X=4.42 $Y=0.19 $X2=3.27 $Y2=0.825
cc_107 N_GND_M1000_b N_Y_c_543_n 0.00155118f $X=-0.045 $Y=0 $X2=4.13 $Y2=0.825
cc_108 N_GND_c_50_p N_Y_c_543_n 8.14297e-19 $X=3.7 $Y=0.825 $X2=4.13 $Y2=0.825
cc_109 N_GND_c_57_p N_Y_c_543_n 0.0075556f $X=4.475 $Y=0.152 $X2=4.13 $Y2=0.825
cc_110 N_GND_c_4_p N_Y_c_543_n 0.00475776f $X=4.42 $Y=0.19 $X2=4.13 $Y2=0.825
cc_111 N_GND_M1000_b N_Y_c_547_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.595
cc_112 N_GND_c_2_p N_Y_c_547_n 0.00134236f $X=0.26 $Y=0.825 $X2=0.69 $Y2=1.595
cc_113 N_GND_c_10_p N_Y_c_547_n 7.53951e-19 $X=1.12 $Y=0.825 $X2=0.69 $Y2=1.595
cc_114 N_GND_M1000_b Y 0.0456345f $X=-0.045 $Y=0 $X2=0.76 $Y2=2.2
cc_115 N_GND_M1002_d N_Y_c_551_n 0.0127699f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1.48
cc_116 N_GND_c_10_p N_Y_c_551_n 0.0142303f $X=1.12 $Y=0.825 $X2=1.405 $Y2=1.48
cc_117 N_GND_M1000_b N_Y_c_553_n 0.0591815f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.845
cc_118 N_GND_M1005_d N_Y_c_554_n 0.0127699f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.48
cc_119 N_GND_c_23_p N_Y_c_554_n 0.0142303f $X=1.98 $Y=0.825 $X2=2.265 $Y2=1.48
cc_120 N_GND_M1000_b N_Y_c_556_n 0.00409378f $X=-0.045 $Y=0 $X2=1.695 $Y2=1.48
cc_121 N_GND_c_10_p N_Y_c_556_n 7.53951e-19 $X=1.12 $Y=0.825 $X2=1.695 $Y2=1.48
cc_122 N_GND_c_23_p N_Y_c_556_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=1.695 $Y2=1.48
cc_123 N_GND_M1000_b N_Y_c_559_n 0.0580131f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.845
cc_124 N_GND_M1010_d N_Y_c_560_n 0.0127699f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.48
cc_125 N_GND_c_37_p N_Y_c_560_n 0.0142303f $X=2.84 $Y=0.825 $X2=3.125 $Y2=1.48
cc_126 N_GND_M1000_b N_Y_c_562_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.48
cc_127 N_GND_c_23_p N_Y_c_562_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=2.555 $Y2=1.48
cc_128 N_GND_c_37_p N_Y_c_562_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=2.555 $Y2=1.48
cc_129 N_GND_M1000_b N_Y_c_565_n 0.0752458f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.845
cc_130 N_GND_M1014_d N_Y_c_566_n 0.0127699f $X=3.56 $Y=0.575 $X2=3.985 $Y2=1.48
cc_131 N_GND_c_50_p N_Y_c_566_n 0.0142303f $X=3.7 $Y=0.825 $X2=3.985 $Y2=1.48
cc_132 N_GND_M1000_b N_Y_c_568_n 0.00409378f $X=-0.045 $Y=0 $X2=3.415 $Y2=1.48
cc_133 N_GND_c_37_p N_Y_c_568_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=3.415 $Y2=1.48
cc_134 N_GND_c_50_p N_Y_c_568_n 7.53951e-19 $X=3.7 $Y=0.825 $X2=3.415 $Y2=1.48
cc_135 N_GND_M1000_b N_Y_c_571_n 0.00409378f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.595
cc_136 N_GND_c_50_p N_Y_c_571_n 7.53951e-19 $X=3.7 $Y=0.825 $X2=4.13 $Y2=1.595
cc_137 N_GND_c_63_p N_Y_c_571_n 0.00134236f $X=4.56 $Y=0.825 $X2=4.13 $Y2=1.595
cc_138 N_GND_M1000_b N_Y_c_574_n 0.0754129f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.845
cc_139 N_VDD_M1001_b N_A_c_322_n 0.0181616f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.96
cc_140 N_VDD_c_140_p N_A_c_322_n 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=2.96
cc_141 N_VDD_c_141_p N_A_c_322_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.475
+ $Y2=2.96
cc_142 N_VDD_c_142_p N_A_c_322_n 0.00468827f $X=4.42 $Y=6.47 $X2=0.475 $Y2=2.96
cc_143 N_VDD_M1001_b N_A_c_241_n 0.00448664f $X=-0.045 $Y=2.905 $X2=0.83
+ $Y2=2.885
cc_144 N_VDD_M1001_b N_A_c_327_n 0.0159283f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=2.96
cc_145 N_VDD_c_141_p N_A_c_327_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.905
+ $Y2=2.96
cc_146 N_VDD_c_146_p N_A_c_327_n 0.00354579f $X=1.12 $Y=3.455 $X2=0.905 $Y2=2.96
cc_147 N_VDD_c_142_p N_A_c_327_n 0.00468827f $X=4.42 $Y=6.47 $X2=0.905 $Y2=2.96
cc_148 N_VDD_M1001_b N_A_c_248_n 0.00500158f $X=-0.045 $Y=2.905 $X2=1.26
+ $Y2=2.885
cc_149 N_VDD_c_146_p N_A_c_248_n 0.00341318f $X=1.12 $Y=3.455 $X2=1.26 $Y2=2.885
cc_150 N_VDD_M1001_b N_A_c_333_n 0.0159283f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.96
cc_151 N_VDD_c_146_p N_A_c_333_n 0.00354579f $X=1.12 $Y=3.455 $X2=1.335 $Y2=2.96
cc_152 N_VDD_c_152_p N_A_c_333_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.335
+ $Y2=2.96
cc_153 N_VDD_c_142_p N_A_c_333_n 0.00468827f $X=4.42 $Y=6.47 $X2=1.335 $Y2=2.96
cc_154 N_VDD_M1001_b N_A_c_254_n 0.00448664f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.885
cc_155 N_VDD_M1001_b N_A_c_338_n 0.0159283f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.96
cc_156 N_VDD_c_152_p N_A_c_338_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.765
+ $Y2=2.96
cc_157 N_VDD_c_157_p N_A_c_338_n 0.00354579f $X=1.98 $Y=3.455 $X2=1.765 $Y2=2.96
cc_158 N_VDD_c_142_p N_A_c_338_n 0.00468827f $X=4.42 $Y=6.47 $X2=1.765 $Y2=2.96
cc_159 N_VDD_M1001_b N_A_c_261_n 0.00500158f $X=-0.045 $Y=2.905 $X2=2.12
+ $Y2=2.885
cc_160 N_VDD_c_157_p N_A_c_261_n 0.00341318f $X=1.98 $Y=3.455 $X2=2.12 $Y2=2.885
cc_161 N_VDD_M1001_b N_A_c_344_n 0.0159283f $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.96
cc_162 N_VDD_c_157_p N_A_c_344_n 0.00354579f $X=1.98 $Y=3.455 $X2=2.195 $Y2=2.96
cc_163 N_VDD_c_163_p N_A_c_344_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.195
+ $Y2=2.96
cc_164 N_VDD_c_142_p N_A_c_344_n 0.00468827f $X=4.42 $Y=6.47 $X2=2.195 $Y2=2.96
cc_165 N_VDD_M1001_b N_A_c_268_n 0.00448664f $X=-0.045 $Y=2.905 $X2=2.55
+ $Y2=2.885
cc_166 N_VDD_M1001_b N_A_c_349_n 0.0159283f $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=2.96
cc_167 N_VDD_c_163_p N_A_c_349_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.625
+ $Y2=2.96
cc_168 N_VDD_c_168_p N_A_c_349_n 0.00354579f $X=2.84 $Y=3.455 $X2=2.625 $Y2=2.96
cc_169 N_VDD_c_142_p N_A_c_349_n 0.00468827f $X=4.42 $Y=6.47 $X2=2.625 $Y2=2.96
cc_170 N_VDD_M1001_b N_A_c_275_n 0.00500158f $X=-0.045 $Y=2.905 $X2=2.98
+ $Y2=2.885
cc_171 N_VDD_c_168_p N_A_c_275_n 0.00341318f $X=2.84 $Y=3.455 $X2=2.98 $Y2=2.885
cc_172 N_VDD_M1001_b N_A_c_355_n 0.0159283f $X=-0.045 $Y=2.905 $X2=3.055
+ $Y2=2.96
cc_173 N_VDD_c_168_p N_A_c_355_n 0.00354579f $X=2.84 $Y=3.455 $X2=3.055 $Y2=2.96
cc_174 N_VDD_c_174_p N_A_c_355_n 0.00606474f $X=3.615 $Y=6.507 $X2=3.055
+ $Y2=2.96
cc_175 N_VDD_c_142_p N_A_c_355_n 0.00468827f $X=4.42 $Y=6.47 $X2=3.055 $Y2=2.96
cc_176 N_VDD_M1001_b N_A_c_281_n 0.00448664f $X=-0.045 $Y=2.905 $X2=3.41
+ $Y2=2.885
cc_177 N_VDD_M1001_b N_A_c_360_n 0.0159283f $X=-0.045 $Y=2.905 $X2=3.485
+ $Y2=2.96
cc_178 N_VDD_c_174_p N_A_c_360_n 0.00606474f $X=3.615 $Y=6.507 $X2=3.485
+ $Y2=2.96
cc_179 N_VDD_c_179_p N_A_c_360_n 0.00354579f $X=3.7 $Y=3.455 $X2=3.485 $Y2=2.96
cc_180 N_VDD_c_142_p N_A_c_360_n 0.00468827f $X=4.42 $Y=6.47 $X2=3.485 $Y2=2.96
cc_181 N_VDD_M1001_b N_A_c_288_n 0.00500158f $X=-0.045 $Y=2.905 $X2=3.84
+ $Y2=2.885
cc_182 N_VDD_c_179_p N_A_c_288_n 0.00341318f $X=3.7 $Y=3.455 $X2=3.84 $Y2=2.885
cc_183 N_VDD_M1001_b N_A_c_366_n 0.0159283f $X=-0.045 $Y=2.905 $X2=3.915
+ $Y2=2.96
cc_184 N_VDD_c_179_p N_A_c_366_n 0.00354579f $X=3.7 $Y=3.455 $X2=3.915 $Y2=2.96
cc_185 N_VDD_c_185_p N_A_c_366_n 0.00606474f $X=4.475 $Y=6.507 $X2=3.915
+ $Y2=2.96
cc_186 N_VDD_c_142_p N_A_c_366_n 0.00468827f $X=4.42 $Y=6.47 $X2=3.915 $Y2=2.96
cc_187 N_VDD_M1001_b N_A_c_294_n 0.00840215f $X=-0.045 $Y=2.905 $X2=4.27
+ $Y2=2.885
cc_188 N_VDD_M1001_b N_A_c_371_n 0.0204783f $X=-0.045 $Y=2.905 $X2=4.345
+ $Y2=2.96
cc_189 N_VDD_c_185_p N_A_c_371_n 0.00606474f $X=4.475 $Y=6.507 $X2=4.345
+ $Y2=2.96
cc_190 N_VDD_c_190_p N_A_c_371_n 0.00713292f $X=4.56 $Y=3.455 $X2=4.345 $Y2=2.96
cc_191 N_VDD_c_142_p N_A_c_371_n 0.00468827f $X=4.42 $Y=6.47 $X2=4.345 $Y2=2.96
cc_192 N_VDD_M1001_b N_A_c_302_n 0.00244521f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.885
cc_193 N_VDD_M1001_b N_A_c_304_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=2.885
cc_194 N_VDD_M1001_b N_A_c_306_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.885
cc_195 N_VDD_M1001_b N_A_c_308_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.885
cc_196 N_VDD_M1001_b N_A_c_310_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.885
cc_197 N_VDD_M1001_b N_A_c_312_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=2.885
cc_198 N_VDD_M1001_b N_A_c_314_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=3.055
+ $Y2=2.885
cc_199 N_VDD_M1001_b N_A_c_316_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=3.485
+ $Y2=2.885
cc_200 N_VDD_M1001_b N_A_c_318_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=3.915
+ $Y2=2.885
cc_201 N_VDD_M1001_d N_A_c_319_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_202 N_VDD_M1001_b N_A_c_319_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.32
+ $Y2=3.33
cc_203 N_VDD_c_140_p N_A_c_319_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_204 N_VDD_M1001_d A 0.0162774f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.325
cc_205 N_VDD_c_140_p A 0.00522047f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.325
cc_206 N_VDD_c_146_p A 9.09141e-19 $X=1.12 $Y=3.455 $X2=0.32 $Y2=3.325
cc_207 N_VDD_M1001_b N_Y_c_575_n 0.00361433f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.96
cc_208 N_VDD_c_141_p N_Y_c_575_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69 $Y2=2.96
cc_209 N_VDD_c_142_p N_Y_c_575_n 0.00475776f $X=4.42 $Y=6.47 $X2=0.69 $Y2=2.96
cc_210 N_VDD_M1001_b N_Y_c_578_n 0.00465961f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=2.96
cc_211 N_VDD_c_152_p N_Y_c_578_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55 $Y2=2.96
cc_212 N_VDD_c_142_p N_Y_c_578_n 0.00475776f $X=4.42 $Y=6.47 $X2=1.55 $Y2=2.96
cc_213 N_VDD_M1001_b N_Y_c_581_n 0.00465961f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.96
cc_214 N_VDD_c_163_p N_Y_c_581_n 0.00734006f $X=2.755 $Y=6.507 $X2=2.41 $Y2=2.96
cc_215 N_VDD_c_142_p N_Y_c_581_n 0.00475776f $X=4.42 $Y=6.47 $X2=2.41 $Y2=2.96
cc_216 N_VDD_M1001_b N_Y_c_584_n 0.00465961f $X=-0.045 $Y=2.905 $X2=3.27
+ $Y2=2.96
cc_217 N_VDD_c_174_p N_Y_c_584_n 0.00745425f $X=3.615 $Y=6.507 $X2=3.27 $Y2=2.96
cc_218 N_VDD_c_142_p N_Y_c_584_n 0.00475776f $X=4.42 $Y=6.47 $X2=3.27 $Y2=2.96
cc_219 N_VDD_M1001_b N_Y_c_587_n 0.00465961f $X=-0.045 $Y=2.905 $X2=4.13
+ $Y2=2.96
cc_220 N_VDD_c_185_p N_Y_c_587_n 0.0075556f $X=4.475 $Y=6.507 $X2=4.13 $Y2=2.96
cc_221 N_VDD_c_142_p N_Y_c_587_n 0.00475776f $X=4.42 $Y=6.47 $X2=4.13 $Y2=2.96
cc_222 N_VDD_M1001_b N_Y_c_590_n 0.00248543f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.845
cc_223 N_VDD_M1001_b N_Y_c_591_n 0.00520877f $X=-0.045 $Y=2.905 $X2=1.405
+ $Y2=2.96
cc_224 N_VDD_c_146_p N_Y_c_591_n 0.0090257f $X=1.12 $Y=3.455 $X2=1.405 $Y2=2.96
cc_225 N_VDD_M1001_b N_Y_c_593_n 0.00520877f $X=-0.045 $Y=2.905 $X2=2.265
+ $Y2=2.96
cc_226 N_VDD_c_157_p N_Y_c_593_n 0.0090257f $X=1.98 $Y=3.455 $X2=2.265 $Y2=2.96
cc_227 N_VDD_M1001_b N_Y_c_595_n 0.00409378f $X=-0.045 $Y=2.905 $X2=1.695
+ $Y2=2.96
cc_228 N_VDD_M1001_b N_Y_c_596_n 0.00520877f $X=-0.045 $Y=2.905 $X2=3.125
+ $Y2=2.96
cc_229 N_VDD_c_168_p N_Y_c_596_n 0.0090257f $X=2.84 $Y=3.455 $X2=3.125 $Y2=2.96
cc_230 N_VDD_M1001_b N_Y_c_598_n 0.00409378f $X=-0.045 $Y=2.905 $X2=2.555
+ $Y2=2.96
cc_231 N_VDD_M1001_b N_Y_c_599_n 0.00520877f $X=-0.045 $Y=2.905 $X2=3.985
+ $Y2=2.96
cc_232 N_VDD_c_179_p N_Y_c_599_n 0.0090257f $X=3.7 $Y=3.455 $X2=3.985 $Y2=2.96
cc_233 N_VDD_M1001_b N_Y_c_601_n 0.00409378f $X=-0.045 $Y=2.905 $X2=3.415
+ $Y2=2.96
cc_234 N_VDD_M1001_b N_Y_c_574_n 0.00409378f $X=-0.045 $Y=2.905 $X2=4.13
+ $Y2=2.845
cc_235 A N_Y_M1001_s 0.00251573f $X=0.32 $Y=3.325 $X2=0.55 $Y2=3.085
cc_236 N_A_c_235_n N_Y_c_524_n 0.00231637f $X=0.475 $Y=1.7 $X2=0.69 $Y2=0.825
cc_237 N_A_c_240_n N_Y_c_524_n 0.00256118f $X=0.83 $Y=1.775 $X2=0.69 $Y2=0.825
cc_238 N_A_c_242_n N_Y_c_524_n 0.00231637f $X=0.905 $Y=1.7 $X2=0.69 $Y2=0.825
cc_239 N_A_c_300_n N_Y_c_524_n 3.64468e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_240 N_A_c_321_n N_Y_c_524_n 0.00110256f $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_241 N_A_c_322_n N_Y_c_575_n 0.00199065f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.96
cc_242 N_A_c_241_n N_Y_c_575_n 0.00899372f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.96
cc_243 N_A_c_327_n N_Y_c_575_n 0.0035213f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.96
cc_244 N_A_c_300_n N_Y_c_575_n 5.06602e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_245 N_A_c_319_n N_Y_c_575_n 0.0226156f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_246 N_A_c_321_n N_Y_c_575_n 0.00165526f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_247 A N_Y_c_575_n 0.00938699f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.96
cc_248 N_A_c_249_n N_Y_c_528_n 0.00231637f $X=1.335 $Y=1.7 $X2=1.55 $Y2=0.825
cc_249 N_A_c_253_n N_Y_c_528_n 0.00317228f $X=1.69 $Y=1.775 $X2=1.55 $Y2=0.825
cc_250 N_A_c_255_n N_Y_c_528_n 0.00231637f $X=1.765 $Y=1.7 $X2=1.55 $Y2=0.825
cc_251 N_A_c_333_n N_Y_c_578_n 0.0035213f $X=1.335 $Y=2.96 $X2=1.55 $Y2=2.96
cc_252 N_A_c_254_n N_Y_c_578_n 0.0108863f $X=1.69 $Y=2.885 $X2=1.55 $Y2=2.96
cc_253 N_A_c_338_n N_Y_c_578_n 0.0035213f $X=1.765 $Y=2.96 $X2=1.55 $Y2=2.96
cc_254 N_A_c_262_n N_Y_c_533_n 0.00231637f $X=2.195 $Y=1.7 $X2=2.41 $Y2=0.825
cc_255 N_A_c_267_n N_Y_c_533_n 0.00317228f $X=2.55 $Y=1.775 $X2=2.41 $Y2=0.825
cc_256 N_A_c_269_n N_Y_c_533_n 0.00231637f $X=2.625 $Y=1.7 $X2=2.41 $Y2=0.825
cc_257 N_A_c_344_n N_Y_c_581_n 0.0035213f $X=2.195 $Y=2.96 $X2=2.41 $Y2=2.96
cc_258 N_A_c_268_n N_Y_c_581_n 0.0108863f $X=2.55 $Y=2.885 $X2=2.41 $Y2=2.96
cc_259 N_A_c_349_n N_Y_c_581_n 0.0035213f $X=2.625 $Y=2.96 $X2=2.41 $Y2=2.96
cc_260 N_A_c_276_n N_Y_c_538_n 0.00231637f $X=3.055 $Y=1.7 $X2=3.27 $Y2=0.825
cc_261 N_A_c_280_n N_Y_c_538_n 0.00317228f $X=3.41 $Y=1.775 $X2=3.27 $Y2=0.825
cc_262 N_A_c_282_n N_Y_c_538_n 0.00231637f $X=3.485 $Y=1.7 $X2=3.27 $Y2=0.825
cc_263 N_A_c_355_n N_Y_c_584_n 0.0035213f $X=3.055 $Y=2.96 $X2=3.27 $Y2=2.96
cc_264 N_A_c_281_n N_Y_c_584_n 0.0108863f $X=3.41 $Y=2.885 $X2=3.27 $Y2=2.96
cc_265 N_A_c_360_n N_Y_c_584_n 0.0035213f $X=3.485 $Y=2.96 $X2=3.27 $Y2=2.96
cc_266 N_A_c_289_n N_Y_c_543_n 0.00231637f $X=3.915 $Y=1.7 $X2=4.13 $Y2=0.825
cc_267 N_A_c_293_n N_Y_c_543_n 0.00317228f $X=4.27 $Y=1.775 $X2=4.13 $Y2=0.825
cc_268 N_A_c_295_n N_Y_c_543_n 0.00231637f $X=4.345 $Y=1.7 $X2=4.13 $Y2=0.825
cc_269 N_A_c_366_n N_Y_c_587_n 0.0035213f $X=3.915 $Y=2.96 $X2=4.13 $Y2=2.96
cc_270 N_A_c_294_n N_Y_c_587_n 0.0105836f $X=4.27 $Y=2.885 $X2=4.13 $Y2=2.96
cc_271 N_A_c_371_n N_Y_c_587_n 0.0035213f $X=4.345 $Y=2.96 $X2=4.13 $Y2=2.96
cc_272 N_A_c_235_n N_Y_c_547_n 0.00942005f $X=0.475 $Y=1.7 $X2=0.69 $Y2=1.595
cc_273 N_A_c_242_n N_Y_c_547_n 0.00259753f $X=0.905 $Y=1.7 $X2=0.69 $Y2=1.595
cc_274 N_A_c_300_n N_Y_c_547_n 0.0011424f $X=0.535 $Y=2.305 $X2=0.69 $Y2=1.595
cc_275 N_A_c_322_n N_Y_c_590_n 0.00169643f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.845
cc_276 N_A_c_241_n N_Y_c_590_n 0.00270155f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.845
cc_277 N_A_c_327_n N_Y_c_590_n 0.00144225f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.845
cc_278 N_A_c_300_n N_Y_c_590_n 8.31386e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.845
cc_279 N_A_c_302_n N_Y_c_590_n 0.00102602f $X=0.475 $Y=2.885 $X2=0.69 $Y2=2.845
cc_280 N_A_c_304_n N_Y_c_590_n 0.00150284f $X=0.905 $Y=2.885 $X2=0.69 $Y2=2.845
cc_281 N_A_c_319_n N_Y_c_590_n 0.0071561f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.845
cc_282 N_A_c_321_n N_Y_c_590_n 0.00173027f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.845
cc_283 A N_Y_c_590_n 0.00815006f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.845
cc_284 N_A_c_235_n Y 0.00150089f $X=0.475 $Y=1.7 $X2=0.76 $Y2=2.2
cc_285 N_A_c_239_n Y 0.00792324f $X=0.475 $Y=2.81 $X2=0.76 $Y2=2.2
cc_286 N_A_c_240_n Y 0.0161013f $X=0.83 $Y=1.775 $X2=0.76 $Y2=2.2
cc_287 N_A_c_241_n Y 0.00363305f $X=0.83 $Y=2.885 $X2=0.76 $Y2=2.2
cc_288 N_A_c_242_n Y 0.00150089f $X=0.905 $Y=1.7 $X2=0.76 $Y2=2.2
cc_289 N_A_c_300_n Y 0.00668675f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_290 N_A_c_301_n Y 0.00675469f $X=0.535 $Y=2.14 $X2=0.76 $Y2=2.2
cc_291 N_A_c_319_n Y 0.0182346f $X=0.32 $Y=3.33 $X2=0.76 $Y2=2.2
cc_292 N_A_c_321_n Y 0.0178517f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_293 N_A_c_242_n N_Y_c_551_n 0.0129682f $X=0.905 $Y=1.7 $X2=1.405 $Y2=1.48
cc_294 N_A_c_246_n N_Y_c_551_n 0.0022289f $X=1.26 $Y=1.775 $X2=1.405 $Y2=1.48
cc_295 N_A_c_249_n N_Y_c_551_n 0.0129682f $X=1.335 $Y=1.7 $X2=1.405 $Y2=1.48
cc_296 N_A_c_327_n N_Y_c_591_n 0.00693713f $X=0.905 $Y=2.96 $X2=1.405 $Y2=2.96
cc_297 N_A_c_248_n N_Y_c_591_n 0.0120397f $X=1.26 $Y=2.885 $X2=1.405 $Y2=2.96
cc_298 N_A_c_333_n N_Y_c_591_n 0.00693713f $X=1.335 $Y=2.96 $X2=1.405 $Y2=2.96
cc_299 N_A_c_304_n N_Y_c_591_n 0.00560085f $X=0.905 $Y=2.885 $X2=1.405 $Y2=2.96
cc_300 N_A_c_306_n N_Y_c_591_n 0.00560085f $X=1.335 $Y=2.885 $X2=1.405 $Y2=2.96
cc_301 N_A_c_249_n N_Y_c_553_n 0.00150089f $X=1.335 $Y=1.7 $X2=1.55 $Y2=2.845
cc_302 N_A_c_253_n N_Y_c_553_n 0.0177499f $X=1.69 $Y=1.775 $X2=1.55 $Y2=2.845
cc_303 N_A_c_254_n N_Y_c_553_n 0.00562481f $X=1.69 $Y=2.885 $X2=1.55 $Y2=2.845
cc_304 N_A_c_255_n N_Y_c_553_n 0.00150089f $X=1.765 $Y=1.7 $X2=1.55 $Y2=2.845
cc_305 N_A_c_266_n N_Y_c_553_n 0.0141566f $X=2.195 $Y=2.81 $X2=1.55 $Y2=2.845
cc_306 N_A_c_255_n N_Y_c_554_n 0.0129682f $X=1.765 $Y=1.7 $X2=2.265 $Y2=1.48
cc_307 N_A_c_259_n N_Y_c_554_n 0.0022289f $X=2.12 $Y=1.775 $X2=2.265 $Y2=1.48
cc_308 N_A_c_262_n N_Y_c_554_n 0.0136594f $X=2.195 $Y=1.7 $X2=2.265 $Y2=1.48
cc_309 N_A_c_249_n N_Y_c_556_n 0.00259753f $X=1.335 $Y=1.7 $X2=1.695 $Y2=1.48
cc_310 N_A_c_255_n N_Y_c_556_n 0.00259753f $X=1.765 $Y=1.7 $X2=1.695 $Y2=1.48
cc_311 N_A_c_338_n N_Y_c_593_n 0.00693713f $X=1.765 $Y=2.96 $X2=2.265 $Y2=2.96
cc_312 N_A_c_261_n N_Y_c_593_n 0.0125508f $X=2.12 $Y=2.885 $X2=2.265 $Y2=2.96
cc_313 N_A_c_344_n N_Y_c_593_n 0.00693713f $X=2.195 $Y=2.96 $X2=2.265 $Y2=2.96
cc_314 N_A_c_308_n N_Y_c_593_n 0.00560085f $X=1.765 $Y=2.885 $X2=2.265 $Y2=2.96
cc_315 N_A_c_310_n N_Y_c_593_n 0.00642784f $X=2.195 $Y=2.885 $X2=2.265 $Y2=2.96
cc_316 N_A_c_333_n N_Y_c_595_n 0.00144225f $X=1.335 $Y=2.96 $X2=1.695 $Y2=2.96
cc_317 N_A_c_254_n N_Y_c_595_n 0.00397642f $X=1.69 $Y=2.885 $X2=1.695 $Y2=2.96
cc_318 N_A_c_338_n N_Y_c_595_n 0.00144225f $X=1.765 $Y=2.96 $X2=1.695 $Y2=2.96
cc_319 N_A_c_306_n N_Y_c_595_n 0.00150284f $X=1.335 $Y=2.885 $X2=1.695 $Y2=2.96
cc_320 N_A_c_308_n N_Y_c_595_n 0.00150284f $X=1.765 $Y=2.885 $X2=1.695 $Y2=2.96
cc_321 N_A_c_262_n N_Y_c_559_n 0.00150089f $X=2.195 $Y=1.7 $X2=2.41 $Y2=2.845
cc_322 N_A_c_266_n N_Y_c_559_n 0.0182294f $X=2.195 $Y=2.81 $X2=2.41 $Y2=2.845
cc_323 N_A_c_267_n N_Y_c_559_n 0.0177499f $X=2.55 $Y=1.775 $X2=2.41 $Y2=2.845
cc_324 N_A_c_268_n N_Y_c_559_n 0.00562481f $X=2.55 $Y=2.885 $X2=2.41 $Y2=2.845
cc_325 N_A_c_269_n N_Y_c_559_n 0.00150089f $X=2.625 $Y=1.7 $X2=2.41 $Y2=2.845
cc_326 N_A_c_269_n N_Y_c_560_n 0.0129682f $X=2.625 $Y=1.7 $X2=3.125 $Y2=1.48
cc_327 N_A_c_273_n N_Y_c_560_n 0.0022289f $X=2.98 $Y=1.775 $X2=3.125 $Y2=1.48
cc_328 N_A_c_276_n N_Y_c_560_n 0.0129682f $X=3.055 $Y=1.7 $X2=3.125 $Y2=1.48
cc_329 N_A_c_262_n N_Y_c_562_n 0.00262362f $X=2.195 $Y=1.7 $X2=2.555 $Y2=1.48
cc_330 N_A_c_269_n N_Y_c_562_n 0.00259753f $X=2.625 $Y=1.7 $X2=2.555 $Y2=1.48
cc_331 N_A_c_349_n N_Y_c_596_n 0.00693713f $X=2.625 $Y=2.96 $X2=3.125 $Y2=2.96
cc_332 N_A_c_275_n N_Y_c_596_n 0.0120397f $X=2.98 $Y=2.885 $X2=3.125 $Y2=2.96
cc_333 N_A_c_355_n N_Y_c_596_n 0.00693713f $X=3.055 $Y=2.96 $X2=3.125 $Y2=2.96
cc_334 N_A_c_312_n N_Y_c_596_n 0.00560085f $X=2.625 $Y=2.885 $X2=3.125 $Y2=2.96
cc_335 N_A_c_314_n N_Y_c_596_n 0.00560085f $X=3.055 $Y=2.885 $X2=3.125 $Y2=2.96
cc_336 N_A_c_344_n N_Y_c_598_n 0.00144225f $X=2.195 $Y=2.96 $X2=2.555 $Y2=2.96
cc_337 N_A_c_268_n N_Y_c_598_n 0.00397642f $X=2.55 $Y=2.885 $X2=2.555 $Y2=2.96
cc_338 N_A_c_349_n N_Y_c_598_n 0.00144225f $X=2.625 $Y=2.96 $X2=2.555 $Y2=2.96
cc_339 N_A_c_310_n N_Y_c_598_n 0.00153387f $X=2.195 $Y=2.885 $X2=2.555 $Y2=2.96
cc_340 N_A_c_312_n N_Y_c_598_n 0.00150284f $X=2.625 $Y=2.885 $X2=2.555 $Y2=2.96
cc_341 N_A_c_276_n N_Y_c_565_n 0.00150089f $X=3.055 $Y=1.7 $X2=3.27 $Y2=2.845
cc_342 N_A_c_280_n N_Y_c_565_n 0.0177499f $X=3.41 $Y=1.775 $X2=3.27 $Y2=2.845
cc_343 N_A_c_281_n N_Y_c_565_n 0.00562481f $X=3.41 $Y=2.885 $X2=3.27 $Y2=2.845
cc_344 N_A_c_282_n N_Y_c_565_n 0.00150089f $X=3.485 $Y=1.7 $X2=3.27 $Y2=2.845
cc_345 N_A_c_282_n N_Y_c_566_n 0.0129682f $X=3.485 $Y=1.7 $X2=3.985 $Y2=1.48
cc_346 N_A_c_286_n N_Y_c_566_n 0.0022289f $X=3.84 $Y=1.775 $X2=3.985 $Y2=1.48
cc_347 N_A_c_289_n N_Y_c_566_n 0.0129682f $X=3.915 $Y=1.7 $X2=3.985 $Y2=1.48
cc_348 N_A_c_276_n N_Y_c_568_n 0.00259753f $X=3.055 $Y=1.7 $X2=3.415 $Y2=1.48
cc_349 N_A_c_282_n N_Y_c_568_n 0.00259753f $X=3.485 $Y=1.7 $X2=3.415 $Y2=1.48
cc_350 N_A_c_360_n N_Y_c_599_n 0.00693713f $X=3.485 $Y=2.96 $X2=3.985 $Y2=2.96
cc_351 N_A_c_288_n N_Y_c_599_n 0.0120397f $X=3.84 $Y=2.885 $X2=3.985 $Y2=2.96
cc_352 N_A_c_366_n N_Y_c_599_n 0.00693713f $X=3.915 $Y=2.96 $X2=3.985 $Y2=2.96
cc_353 N_A_c_316_n N_Y_c_599_n 0.00560085f $X=3.485 $Y=2.885 $X2=3.985 $Y2=2.96
cc_354 N_A_c_318_n N_Y_c_599_n 0.00560085f $X=3.915 $Y=2.885 $X2=3.985 $Y2=2.96
cc_355 N_A_c_355_n N_Y_c_601_n 0.00144225f $X=3.055 $Y=2.96 $X2=3.415 $Y2=2.96
cc_356 N_A_c_281_n N_Y_c_601_n 0.00397642f $X=3.41 $Y=2.885 $X2=3.415 $Y2=2.96
cc_357 N_A_c_360_n N_Y_c_601_n 0.00144225f $X=3.485 $Y=2.96 $X2=3.415 $Y2=2.96
cc_358 N_A_c_314_n N_Y_c_601_n 0.00150284f $X=3.055 $Y=2.885 $X2=3.415 $Y2=2.96
cc_359 N_A_c_316_n N_Y_c_601_n 0.00150284f $X=3.485 $Y=2.885 $X2=3.415 $Y2=2.96
cc_360 N_A_c_289_n N_Y_c_571_n 0.00259753f $X=3.915 $Y=1.7 $X2=4.13 $Y2=1.595
cc_361 N_A_c_295_n N_Y_c_571_n 0.00939395f $X=4.345 $Y=1.7 $X2=4.13 $Y2=1.595
cc_362 N_A_c_289_n N_Y_c_574_n 0.00150089f $X=3.915 $Y=1.7 $X2=4.13 $Y2=2.845
cc_363 N_A_c_366_n N_Y_c_574_n 0.00144225f $X=3.915 $Y=2.96 $X2=4.13 $Y2=2.845
cc_364 N_A_c_293_n N_Y_c_574_n 0.0169795f $X=4.27 $Y=1.775 $X2=4.13 $Y2=2.845
cc_365 N_A_c_294_n N_Y_c_574_n 0.0141541f $X=4.27 $Y=2.885 $X2=4.13 $Y2=2.845
cc_366 N_A_c_295_n N_Y_c_574_n 0.00150089f $X=4.345 $Y=1.7 $X2=4.13 $Y2=2.845
cc_367 N_A_c_371_n N_Y_c_574_n 0.00541616f $X=4.345 $Y=2.96 $X2=4.13 $Y2=2.845
cc_368 N_A_c_318_n N_Y_c_574_n 0.00150284f $X=3.915 $Y=2.885 $X2=4.13 $Y2=2.845
