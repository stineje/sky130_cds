* File: sky130_osu_sc_18T_ls__and2_6.pxi.spice
* Created: Fri Nov 12 13:39:22 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__AND2_6%GND N_GND_M1001_d N_GND_M1009_s N_GND_M1012_s
+ N_GND_M1015_s N_GND_M1006_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p N_GND_c_23_p
+ N_GND_c_30_p N_GND_c_36_p N_GND_c_43_p N_GND_c_50_p GND N_GND_c_3_p
+ PM_SKY130_OSU_SC_18T_LS__AND2_6%GND
x_PM_SKY130_OSU_SC_18T_LS__AND2_6%VDD N_VDD_M1005_s N_VDD_M1014_d N_VDD_M1003_d
+ N_VDD_M1007_d N_VDD_M1011_d N_VDD_M1005_b N_VDD_c_107_p N_VDD_c_108_p
+ N_VDD_c_119_p N_VDD_c_126_p N_VDD_c_132_p N_VDD_c_138_p N_VDD_c_143_p
+ N_VDD_c_149_p N_VDD_c_154_p VDD N_VDD_c_109_p
+ PM_SKY130_OSU_SC_18T_LS__AND2_6%VDD
x_PM_SKY130_OSU_SC_18T_LS__AND2_6%A N_A_M1006_g N_A_M1005_g N_A_c_179_n
+ N_A_c_180_n A PM_SKY130_OSU_SC_18T_LS__AND2_6%A
x_PM_SKY130_OSU_SC_18T_LS__AND2_6%B N_B_M1001_g N_B_M1014_g N_B_c_210_n
+ N_B_c_211_n B PM_SKY130_OSU_SC_18T_LS__AND2_6%B
x_PM_SKY130_OSU_SC_18T_LS__AND2_6%A_27_115# N_A_27_115#_M1006_s
+ N_A_27_115#_M1005_d N_A_27_115#_M1000_g N_A_27_115#_c_247_n
+ N_A_27_115#_c_298_n N_A_27_115#_M1002_g N_A_27_115#_c_248_n
+ N_A_27_115#_c_249_n N_A_27_115#_M1009_g N_A_27_115#_c_303_n
+ N_A_27_115#_M1003_g N_A_27_115#_c_254_n N_A_27_115#_c_256_n
+ N_A_27_115#_M1010_g N_A_27_115#_c_310_n N_A_27_115#_M1004_g
+ N_A_27_115#_c_261_n N_A_27_115#_c_262_n N_A_27_115#_M1012_g
+ N_A_27_115#_c_315_n N_A_27_115#_M1007_g N_A_27_115#_c_267_n
+ N_A_27_115#_c_269_n N_A_27_115#_M1013_g N_A_27_115#_c_274_n
+ N_A_27_115#_c_321_n N_A_27_115#_M1008_g N_A_27_115#_c_275_n
+ N_A_27_115#_c_276_n N_A_27_115#_M1015_g N_A_27_115#_c_326_n
+ N_A_27_115#_M1011_g N_A_27_115#_c_281_n N_A_27_115#_c_282_n
+ N_A_27_115#_c_283_n N_A_27_115#_c_284_n N_A_27_115#_c_285_n
+ N_A_27_115#_c_286_n N_A_27_115#_c_287_n N_A_27_115#_c_288_n
+ N_A_27_115#_c_289_n N_A_27_115#_c_290_n N_A_27_115#_c_291_n
+ N_A_27_115#_c_294_n N_A_27_115#_c_336_n N_A_27_115#_c_295_n
+ N_A_27_115#_c_296_n N_A_27_115#_c_348_n
+ PM_SKY130_OSU_SC_18T_LS__AND2_6%A_27_115#
x_PM_SKY130_OSU_SC_18T_LS__AND2_6%Y N_Y_M1000_d N_Y_M1010_d N_Y_M1013_d
+ N_Y_M1002_s N_Y_M1004_s N_Y_M1008_s N_Y_c_431_n N_Y_c_436_n N_Y_c_437_n
+ N_Y_c_442_n N_Y_c_443_n N_Y_c_447_n N_Y_c_448_n N_Y_c_451_n Y N_Y_c_453_n
+ N_Y_c_455_n N_Y_c_456_n N_Y_c_457_n N_Y_c_459_n N_Y_c_462_n N_Y_c_463_n
+ N_Y_c_464_n N_Y_c_467_n PM_SKY130_OSU_SC_18T_LS__AND2_6%Y
cc_1 N_GND_M1006_b N_A_M1006_g 0.0805447f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1006_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1006_g 0.00468827f $X=3.06 $Y=0.19 $X2=0.475 $Y2=1.075
cc_4 N_GND_M1006_b N_A_c_179_n 0.0447183f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_5 N_GND_M1006_b N_A_c_180_n 0.00329519f $X=-0.045 $Y=0 $X2=0.235 $Y2=2.765
cc_6 N_GND_M1006_b N_B_M1001_g 0.0456699f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_7 N_GND_c_2_p N_B_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=1.075
cc_8 N_GND_c_8_p N_B_M1001_g 0.00376152f $X=1.05 $Y=0.825 $X2=0.835 $Y2=1.075
cc_9 N_GND_c_3_p N_B_M1001_g 0.00468827f $X=3.06 $Y=0.19 $X2=0.835 $Y2=1.075
cc_10 N_GND_M1006_b N_B_M1014_g 0.0145087f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_11 N_GND_M1006_b N_B_c_210_n 0.0304191f $X=-0.045 $Y=0 $X2=0.915 $Y2=2.425
cc_12 N_GND_M1006_b N_B_c_211_n 0.00352155f $X=-0.045 $Y=0 $X2=0.915 $Y2=2.425
cc_13 N_GND_M1006_b B 0.00685421f $X=-0.045 $Y=0 $X2=0.92 $Y2=2.96
cc_14 N_GND_M1006_b N_A_27_115#_M1000_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_15 N_GND_c_8_p N_A_27_115#_M1000_g 0.0103278f $X=1.05 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_16 N_GND_c_16_p N_A_27_115#_M1000_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=3.06 $Y=0.19 $X2=1.335
+ $Y2=1.075
cc_18 N_GND_M1006_b N_A_27_115#_c_247_n 0.0465667f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=2.81
cc_19 N_GND_M1006_b N_A_27_115#_c_248_n 0.00863342f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.885
cc_20 N_GND_M1006_b N_A_27_115#_c_249_n 0.0104564f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.845
cc_21 N_GND_M1006_b N_A_27_115#_M1009_g 0.0202142f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_22 N_GND_c_16_p N_A_27_115#_M1009_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=1.075
cc_23 N_GND_c_23_p N_A_27_115#_M1009_g 0.00356864f $X=1.98 $Y=0.825 $X2=1.765
+ $Y2=1.075
cc_24 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=3.06 $Y=0.19 $X2=1.765
+ $Y2=1.075
cc_25 N_GND_M1006_b N_A_27_115#_c_254_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.845
cc_26 N_GND_c_23_p N_A_27_115#_c_254_n 0.00256938f $X=1.98 $Y=0.825 $X2=2.12
+ $Y2=1.845
cc_27 N_GND_M1006_b N_A_27_115#_c_256_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.885
cc_28 N_GND_M1006_b N_A_27_115#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.075
cc_29 N_GND_c_23_p N_A_27_115#_M1010_g 0.00356864f $X=1.98 $Y=0.825 $X2=2.195
+ $Y2=1.075
cc_30 N_GND_c_30_p N_A_27_115#_M1010_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=1.075
cc_31 N_GND_c_3_p N_A_27_115#_M1010_g 0.00468827f $X=3.06 $Y=0.19 $X2=2.195
+ $Y2=1.075
cc_32 N_GND_M1006_b N_A_27_115#_c_261_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.845
cc_33 N_GND_M1006_b N_A_27_115#_c_262_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.885
cc_34 N_GND_M1006_b N_A_27_115#_M1012_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.075
cc_35 N_GND_c_30_p N_A_27_115#_M1012_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=1.075
cc_36 N_GND_c_36_p N_A_27_115#_M1012_g 0.00356864f $X=2.84 $Y=0.825 $X2=2.625
+ $Y2=1.075
cc_37 N_GND_c_3_p N_A_27_115#_M1012_g 0.00468827f $X=3.06 $Y=0.19 $X2=2.625
+ $Y2=1.075
cc_38 N_GND_M1006_b N_A_27_115#_c_267_n 0.0181078f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.845
cc_39 N_GND_c_36_p N_A_27_115#_c_267_n 0.00256938f $X=2.84 $Y=0.825 $X2=2.98
+ $Y2=1.845
cc_40 N_GND_M1006_b N_A_27_115#_c_269_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.885
cc_41 N_GND_M1006_b N_A_27_115#_M1013_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.075
cc_42 N_GND_c_36_p N_A_27_115#_M1013_g 0.00356864f $X=2.84 $Y=0.825 $X2=3.055
+ $Y2=1.075
cc_43 N_GND_c_43_p N_A_27_115#_M1013_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.055
+ $Y2=1.075
cc_44 N_GND_c_3_p N_A_27_115#_M1013_g 0.00468827f $X=3.06 $Y=0.19 $X2=3.055
+ $Y2=1.075
cc_45 N_GND_M1006_b N_A_27_115#_c_274_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.81
cc_46 N_GND_M1006_b N_A_27_115#_c_275_n 0.0369419f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.845
cc_47 N_GND_M1006_b N_A_27_115#_c_276_n 0.0268552f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.885
cc_48 N_GND_M1006_b N_A_27_115#_M1015_g 0.0264941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.075
cc_49 N_GND_c_43_p N_A_27_115#_M1015_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.485
+ $Y2=1.075
cc_50 N_GND_c_50_p N_A_27_115#_M1015_g 0.00713292f $X=3.7 $Y=0.825 $X2=3.485
+ $Y2=1.075
cc_51 N_GND_c_3_p N_A_27_115#_M1015_g 0.00468827f $X=3.06 $Y=0.19 $X2=3.485
+ $Y2=1.075
cc_52 N_GND_M1006_b N_A_27_115#_c_281_n 0.0264756f $X=-0.045 $Y=0 $X2=1.395
+ $Y2=1.845
cc_53 N_GND_M1006_b N_A_27_115#_c_282_n 0.00339913f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=2.885
cc_54 N_GND_M1006_b N_A_27_115#_c_283_n 0.00873941f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.845
cc_55 N_GND_M1006_b N_A_27_115#_c_284_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.885
cc_56 N_GND_M1006_b N_A_27_115#_c_285_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.845
cc_57 N_GND_M1006_b N_A_27_115#_c_286_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.885
cc_58 N_GND_M1006_b N_A_27_115#_c_287_n 0.00873941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.845
cc_59 N_GND_M1006_b N_A_27_115#_c_288_n 0.00735657f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.885
cc_60 N_GND_M1006_b N_A_27_115#_c_289_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.845
cc_61 N_GND_M1006_b N_A_27_115#_c_290_n 0.00151234f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.885
cc_62 N_GND_M1006_b N_A_27_115#_c_291_n 0.0148636f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_63 N_GND_c_2_p N_A_27_115#_c_291_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_64 N_GND_c_3_p N_A_27_115#_c_291_n 0.00476261f $X=3.06 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_65 N_GND_M1006_b N_A_27_115#_c_294_n 0.00626966f $X=-0.045 $Y=0 $X2=0.575
+ $Y2=3.545
cc_66 N_GND_M1006_b N_A_27_115#_c_295_n 0.0164401f $X=-0.045 $Y=0 $X2=0.66
+ $Y2=1.935
cc_67 N_GND_M1006_b N_A_27_115#_c_296_n 0.0251886f $X=-0.045 $Y=0 $X2=1.395
+ $Y2=1.935
cc_68 N_GND_c_8_p N_A_27_115#_c_296_n 0.00704977f $X=1.05 $Y=0.825 $X2=1.395
+ $Y2=1.935
cc_69 N_GND_M1006_b N_Y_c_431_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_70 N_GND_c_8_p N_Y_c_431_n 0.0187614f $X=1.05 $Y=0.825 $X2=1.55 $Y2=0.825
cc_71 N_GND_c_16_p N_Y_c_431_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.825
cc_72 N_GND_c_23_p N_Y_c_431_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=0.825
cc_73 N_GND_c_3_p N_Y_c_431_n 0.00475776f $X=3.06 $Y=0.19 $X2=1.55 $Y2=0.825
cc_74 N_GND_M1006_b N_Y_c_436_n 0.0110121f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_75 N_GND_M1006_b N_Y_c_437_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.825
cc_76 N_GND_c_23_p N_Y_c_437_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=0.825
cc_77 N_GND_c_30_p N_Y_c_437_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.825
cc_78 N_GND_c_36_p N_Y_c_437_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=2.41 $Y2=0.825
cc_79 N_GND_c_3_p N_Y_c_437_n 0.00475776f $X=3.06 $Y=0.19 $X2=2.41 $Y2=0.825
cc_80 N_GND_M1006_b N_Y_c_442_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.59
cc_81 N_GND_M1006_b N_Y_c_443_n 0.00155118f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.825
cc_82 N_GND_c_36_p N_Y_c_443_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=3.27 $Y2=0.825
cc_83 N_GND_c_43_p N_Y_c_443_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.825
cc_84 N_GND_c_3_p N_Y_c_443_n 0.00475776f $X=3.06 $Y=0.19 $X2=3.27 $Y2=0.825
cc_85 N_GND_M1006_b N_Y_c_447_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.59
cc_86 N_GND_M1006_b N_Y_c_448_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.595
cc_87 N_GND_c_8_p N_Y_c_448_n 0.00127231f $X=1.05 $Y=0.825 $X2=1.55 $Y2=1.595
cc_88 N_GND_c_23_p N_Y_c_448_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=1.595
cc_89 N_GND_M1006_b N_Y_c_451_n 0.00675046f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.475
cc_90 N_GND_M1006_b Y 0.030773f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_91 N_GND_M1009_s N_Y_c_453_n 0.0127884f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.48
cc_92 N_GND_c_23_p N_Y_c_453_n 0.0142303f $X=1.98 $Y=0.825 $X2=2.265 $Y2=1.48
cc_93 N_GND_M1006_b N_Y_c_455_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.59
cc_94 N_GND_M1006_b N_Y_c_456_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.475
cc_95 N_GND_M1012_s N_Y_c_457_n 0.0127884f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.48
cc_96 N_GND_c_36_p N_Y_c_457_n 0.0142303f $X=2.84 $Y=0.825 $X2=3.125 $Y2=1.48
cc_97 N_GND_M1006_b N_Y_c_459_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.48
cc_98 N_GND_c_23_p N_Y_c_459_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=2.555 $Y2=1.48
cc_99 N_GND_c_36_p N_Y_c_459_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=2.555 $Y2=1.48
cc_100 N_GND_M1006_b N_Y_c_462_n 0.0144211f $X=-0.045 $Y=0 $X2=3.125 $Y2=2.59
cc_101 N_GND_M1006_b N_Y_c_463_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.59
cc_102 N_GND_M1006_b N_Y_c_464_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.595
cc_103 N_GND_c_36_p N_Y_c_464_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=3.27 $Y2=1.595
cc_104 N_GND_c_50_p N_Y_c_464_n 0.00134236f $X=3.7 $Y=0.825 $X2=3.27 $Y2=1.595
cc_105 N_GND_M1006_b N_Y_c_467_n 0.0485933f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.475
cc_106 N_VDD_M1005_b N_A_M1005_g 0.0189715f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_107 N_VDD_c_107_p N_A_M1005_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_108 N_VDD_c_108_p N_A_M1005_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_109 N_VDD_c_109_p N_A_M1005_g 0.00468827f $X=3.06 $Y=6.47 $X2=0.475 $Y2=4.585
cc_110 N_VDD_M1005_b N_A_c_179_n 0.0124943f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.765
cc_111 N_VDD_M1005_s N_A_c_180_n 0.0150633f $X=0.135 $Y=3.085 $X2=0.235
+ $Y2=2.765
cc_112 N_VDD_M1005_b N_A_c_180_n 0.00613107f $X=-0.045 $Y=2.905 $X2=0.235
+ $Y2=2.765
cc_113 N_VDD_c_107_p N_A_c_180_n 0.00337102f $X=0.26 $Y=4.135 $X2=0.235
+ $Y2=2.765
cc_114 N_VDD_M1005_s A 0.00790556f $X=0.135 $Y=3.085 $X2=0.24 $Y2=3.33
cc_115 N_VDD_M1005_b A 0.0115315f $X=-0.045 $Y=2.905 $X2=0.24 $Y2=3.33
cc_116 N_VDD_c_107_p A 0.00459217f $X=0.26 $Y=4.135 $X2=0.24 $Y2=3.33
cc_117 N_VDD_M1005_b N_B_M1014_g 0.0187479f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_118 N_VDD_c_108_p N_B_M1014_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905
+ $Y2=4.585
cc_119 N_VDD_c_119_p N_B_M1014_g 0.00354579f $X=1.12 $Y=3.795 $X2=0.905
+ $Y2=4.585
cc_120 N_VDD_c_109_p N_B_M1014_g 0.00468827f $X=3.06 $Y=6.47 $X2=0.905 $Y2=4.585
cc_121 N_VDD_M1005_b N_B_c_211_n 0.00130234f $X=-0.045 $Y=2.905 $X2=0.915
+ $Y2=2.425
cc_122 N_VDD_M1005_b B 0.00872506f $X=-0.045 $Y=2.905 $X2=0.92 $Y2=2.96
cc_123 N_VDD_c_119_p B 9.65504e-19 $X=1.12 $Y=3.795 $X2=0.92 $Y2=2.96
cc_124 N_VDD_M1005_b N_A_27_115#_c_298_n 0.0171069f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.96
cc_125 N_VDD_c_119_p N_A_27_115#_c_298_n 0.00354579f $X=1.12 $Y=3.795 $X2=1.335
+ $Y2=2.96
cc_126 N_VDD_c_126_p N_A_27_115#_c_298_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.335
+ $Y2=2.96
cc_127 N_VDD_c_109_p N_A_27_115#_c_298_n 0.00468827f $X=3.06 $Y=6.47 $X2=1.335
+ $Y2=2.96
cc_128 N_VDD_M1005_b N_A_27_115#_c_248_n 0.00448664f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.885
cc_129 N_VDD_M1005_b N_A_27_115#_c_303_n 0.017006f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.96
cc_130 N_VDD_c_119_p N_A_27_115#_c_303_n 3.67508e-19 $X=1.12 $Y=3.795 $X2=1.765
+ $Y2=2.96
cc_131 N_VDD_c_126_p N_A_27_115#_c_303_n 0.00610567f $X=1.895 $Y=6.507 $X2=1.765
+ $Y2=2.96
cc_132 N_VDD_c_132_p N_A_27_115#_c_303_n 0.00373985f $X=1.98 $Y=3.455 $X2=1.765
+ $Y2=2.96
cc_133 N_VDD_c_109_p N_A_27_115#_c_303_n 0.00470215f $X=3.06 $Y=6.47 $X2=1.765
+ $Y2=2.96
cc_134 N_VDD_M1005_b N_A_27_115#_c_256_n 0.00396043f $X=-0.045 $Y=2.905 $X2=2.12
+ $Y2=2.885
cc_135 N_VDD_c_132_p N_A_27_115#_c_256_n 0.00379272f $X=1.98 $Y=3.455 $X2=2.12
+ $Y2=2.885
cc_136 N_VDD_M1005_b N_A_27_115#_c_310_n 0.0166898f $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.96
cc_137 N_VDD_c_132_p N_A_27_115#_c_310_n 0.00354579f $X=1.98 $Y=3.455 $X2=2.195
+ $Y2=2.96
cc_138 N_VDD_c_138_p N_A_27_115#_c_310_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.195
+ $Y2=2.96
cc_139 N_VDD_c_109_p N_A_27_115#_c_310_n 0.00468827f $X=3.06 $Y=6.47 $X2=2.195
+ $Y2=2.96
cc_140 N_VDD_M1005_b N_A_27_115#_c_262_n 0.00448664f $X=-0.045 $Y=2.905 $X2=2.55
+ $Y2=2.885
cc_141 N_VDD_M1005_b N_A_27_115#_c_315_n 0.0166898f $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=2.96
cc_142 N_VDD_c_138_p N_A_27_115#_c_315_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.625
+ $Y2=2.96
cc_143 N_VDD_c_143_p N_A_27_115#_c_315_n 0.00354579f $X=2.84 $Y=3.455 $X2=2.625
+ $Y2=2.96
cc_144 N_VDD_c_109_p N_A_27_115#_c_315_n 0.00468827f $X=3.06 $Y=6.47 $X2=2.625
+ $Y2=2.96
cc_145 N_VDD_M1005_b N_A_27_115#_c_269_n 0.00396043f $X=-0.045 $Y=2.905 $X2=2.98
+ $Y2=2.885
cc_146 N_VDD_c_143_p N_A_27_115#_c_269_n 0.00379272f $X=2.84 $Y=3.455 $X2=2.98
+ $Y2=2.885
cc_147 N_VDD_M1005_b N_A_27_115#_c_321_n 0.0166898f $X=-0.045 $Y=2.905 $X2=3.055
+ $Y2=2.96
cc_148 N_VDD_c_143_p N_A_27_115#_c_321_n 0.00354579f $X=2.84 $Y=3.455 $X2=3.055
+ $Y2=2.96
cc_149 N_VDD_c_149_p N_A_27_115#_c_321_n 0.00606474f $X=3.615 $Y=6.507 $X2=3.055
+ $Y2=2.96
cc_150 N_VDD_c_109_p N_A_27_115#_c_321_n 0.00468827f $X=3.06 $Y=6.47 $X2=3.055
+ $Y2=2.96
cc_151 N_VDD_M1005_b N_A_27_115#_c_276_n 0.00840215f $X=-0.045 $Y=2.905 $X2=3.41
+ $Y2=2.885
cc_152 N_VDD_M1005_b N_A_27_115#_c_326_n 0.0209036f $X=-0.045 $Y=2.905 $X2=3.485
+ $Y2=2.96
cc_153 N_VDD_c_149_p N_A_27_115#_c_326_n 0.00606474f $X=3.615 $Y=6.507 $X2=3.485
+ $Y2=2.96
cc_154 N_VDD_c_154_p N_A_27_115#_c_326_n 0.00713292f $X=3.7 $Y=3.455 $X2=3.485
+ $Y2=2.96
cc_155 N_VDD_c_109_p N_A_27_115#_c_326_n 0.00468827f $X=3.06 $Y=6.47 $X2=3.485
+ $Y2=2.96
cc_156 N_VDD_M1005_b N_A_27_115#_c_282_n 0.00196792f $X=-0.045 $Y=2.905
+ $X2=1.335 $Y2=2.885
cc_157 N_VDD_M1005_b N_A_27_115#_c_284_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.885
cc_158 N_VDD_M1005_b N_A_27_115#_c_286_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.885
cc_159 N_VDD_M1005_b N_A_27_115#_c_288_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=2.885
cc_160 N_VDD_M1005_b N_A_27_115#_c_290_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=3.055 $Y2=2.885
cc_161 N_VDD_M1005_b N_A_27_115#_c_294_n 8.35397e-19 $X=-0.045 $Y=2.905
+ $X2=0.575 $Y2=3.545
cc_162 N_VDD_M1005_b N_A_27_115#_c_336_n 0.00155118f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=3.795
cc_163 N_VDD_c_108_p N_A_27_115#_c_336_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69
+ $Y2=3.795
cc_164 N_VDD_c_109_p N_A_27_115#_c_336_n 0.00475776f $X=3.06 $Y=6.47 $X2=0.69
+ $Y2=3.795
cc_165 N_VDD_M1005_b N_Y_c_436_n 0.00347838f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=2.59
cc_166 N_VDD_c_126_p N_Y_c_436_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55 $Y2=2.59
cc_167 N_VDD_c_109_p N_Y_c_436_n 0.00475776f $X=3.06 $Y=6.47 $X2=1.55 $Y2=2.59
cc_168 N_VDD_M1005_b N_Y_c_442_n 0.00380347f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.59
cc_169 N_VDD_c_138_p N_Y_c_442_n 0.00734006f $X=2.755 $Y=6.507 $X2=2.41 $Y2=2.59
cc_170 N_VDD_c_109_p N_Y_c_442_n 0.00475776f $X=3.06 $Y=6.47 $X2=2.41 $Y2=2.59
cc_171 N_VDD_M1005_b N_Y_c_447_n 0.00380347f $X=-0.045 $Y=2.905 $X2=3.27
+ $Y2=2.59
cc_172 N_VDD_c_149_p N_Y_c_447_n 0.00745425f $X=3.615 $Y=6.507 $X2=3.27 $Y2=2.59
cc_173 N_VDD_c_109_p N_Y_c_447_n 0.00475776f $X=3.06 $Y=6.47 $X2=3.27 $Y2=2.59
cc_174 N_VDD_c_132_p N_Y_c_455_n 0.00634153f $X=1.98 $Y=3.455 $X2=2.265 $Y2=2.59
cc_175 N_VDD_c_143_p N_Y_c_462_n 0.00634153f $X=2.84 $Y=3.455 $X2=3.125 $Y2=2.59
cc_176 N_A_M1006_g N_B_M1001_g 0.129389f $X=0.475 $Y=1.075 $X2=0.835 $Y2=1.075
cc_177 N_A_M1006_g N_B_M1014_g 0.0497852f $X=0.475 $Y=1.075 $X2=0.905 $Y2=4.585
cc_178 N_A_M1006_g N_B_c_211_n 8.69605e-19 $X=0.475 $Y=1.075 $X2=0.915 $Y2=2.425
cc_179 N_A_M1006_g N_A_27_115#_c_291_n 0.0158254f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_180 N_A_M1006_g N_A_27_115#_c_294_n 0.0278506f $X=0.475 $Y=1.075 $X2=0.575
+ $Y2=3.545
cc_181 N_A_M1005_g N_A_27_115#_c_294_n 0.0152191f $X=0.475 $Y=4.585 $X2=0.575
+ $Y2=3.545
cc_182 N_A_c_179_n N_A_27_115#_c_294_n 0.00844699f $X=0.475 $Y=2.765 $X2=0.575
+ $Y2=3.545
cc_183 N_A_c_180_n N_A_27_115#_c_294_n 0.053763f $X=0.235 $Y=2.765 $X2=0.575
+ $Y2=3.545
cc_184 A N_A_27_115#_c_294_n 0.00781918f $X=0.24 $Y=3.33 $X2=0.575 $Y2=3.545
cc_185 N_A_M1006_g N_A_27_115#_c_295_n 0.0178909f $X=0.475 $Y=1.075 $X2=0.66
+ $Y2=1.935
cc_186 N_A_c_179_n N_A_27_115#_c_295_n 0.00272689f $X=0.475 $Y=2.765 $X2=0.66
+ $Y2=1.935
cc_187 N_A_c_180_n N_A_27_115#_c_295_n 0.00451097f $X=0.235 $Y=2.765 $X2=0.66
+ $Y2=1.935
cc_188 N_A_M1005_g N_A_27_115#_c_348_n 0.0109054f $X=0.475 $Y=4.585 $X2=0.69
+ $Y2=3.63
cc_189 N_B_M1001_g N_A_27_115#_M1000_g 0.0468623f $X=0.835 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_190 N_B_M1014_g N_A_27_115#_c_247_n 0.0492452f $X=0.905 $Y=4.585 $X2=1.335
+ $Y2=2.81
cc_191 N_B_c_210_n N_A_27_115#_c_247_n 0.0207593f $X=0.915 $Y=2.425 $X2=1.335
+ $Y2=2.81
cc_192 N_B_c_211_n N_A_27_115#_c_247_n 0.00498982f $X=0.915 $Y=2.425 $X2=1.335
+ $Y2=2.81
cc_193 B N_A_27_115#_c_282_n 0.00380362f $X=0.92 $Y=2.96 $X2=1.335 $Y2=2.885
cc_194 N_B_M1001_g N_A_27_115#_c_294_n 0.00719886f $X=0.835 $Y=1.075 $X2=0.575
+ $Y2=3.545
cc_195 N_B_M1014_g N_A_27_115#_c_294_n 0.01267f $X=0.905 $Y=4.585 $X2=0.575
+ $Y2=3.545
cc_196 N_B_c_211_n N_A_27_115#_c_294_n 0.0541394f $X=0.915 $Y=2.425 $X2=0.575
+ $Y2=3.545
cc_197 B N_A_27_115#_c_294_n 0.00871807f $X=0.92 $Y=2.96 $X2=0.575 $Y2=3.545
cc_198 N_B_M1001_g N_A_27_115#_c_296_n 0.0171085f $X=0.835 $Y=1.075 $X2=1.395
+ $Y2=1.935
cc_199 N_B_c_210_n N_A_27_115#_c_296_n 0.00235847f $X=0.915 $Y=2.425 $X2=1.395
+ $Y2=1.935
cc_200 N_B_c_211_n N_A_27_115#_c_296_n 0.0100447f $X=0.915 $Y=2.425 $X2=1.395
+ $Y2=1.935
cc_201 B N_A_27_115#_c_348_n 0.00385574f $X=0.92 $Y=2.96 $X2=0.69 $Y2=3.63
cc_202 N_B_c_211_n N_Y_c_436_n 0.0138653f $X=0.915 $Y=2.425 $X2=1.55 $Y2=2.59
cc_203 B N_Y_c_436_n 0.00632423f $X=0.92 $Y=2.96 $X2=1.55 $Y2=2.59
cc_204 N_B_M1001_g N_Y_c_448_n 8.18972e-19 $X=0.835 $Y=1.075 $X2=1.55 $Y2=1.595
cc_205 N_B_c_210_n N_Y_c_451_n 5.80618e-19 $X=0.915 $Y=2.425 $X2=1.55 $Y2=2.475
cc_206 N_B_c_211_n N_Y_c_451_n 0.00573285f $X=0.915 $Y=2.425 $X2=1.55 $Y2=2.475
cc_207 N_B_M1001_g Y 6.5988e-19 $X=0.835 $Y=1.075 $X2=1.555 $Y2=2.22
cc_208 N_B_c_211_n Y 0.00671947f $X=0.915 $Y=2.425 $X2=1.555 $Y2=2.22
cc_209 N_A_27_115#_M1000_g N_Y_c_431_n 0.00233629f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_210 N_A_27_115#_M1009_g N_Y_c_431_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_211 N_A_27_115#_c_281_n N_Y_c_431_n 0.00208849f $X=1.395 $Y=1.845 $X2=1.55
+ $Y2=0.825
cc_212 N_A_27_115#_c_296_n N_Y_c_431_n 0.00364905f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_213 N_A_27_115#_c_247_n N_Y_c_436_n 0.00711959f $X=1.335 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_214 N_A_27_115#_c_298_n N_Y_c_436_n 0.00282264f $X=1.335 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_215 N_A_27_115#_c_248_n N_Y_c_436_n 0.0163883f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.59
cc_216 N_A_27_115#_c_249_n N_Y_c_436_n 0.00122399f $X=1.69 $Y=1.845 $X2=1.55
+ $Y2=2.59
cc_217 N_A_27_115#_c_303_n N_Y_c_436_n 0.00392729f $X=1.765 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_218 N_A_27_115#_c_281_n N_Y_c_436_n 6.59752e-19 $X=1.395 $Y=1.845 $X2=1.55
+ $Y2=2.59
cc_219 N_A_27_115#_c_296_n N_Y_c_436_n 0.00202105f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_220 N_A_27_115#_M1010_g N_Y_c_437_n 0.00231637f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_221 N_A_27_115#_c_261_n N_Y_c_437_n 0.00280419f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=0.825
cc_222 N_A_27_115#_M1012_g N_Y_c_437_n 0.00231637f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_223 N_A_27_115#_c_310_n N_Y_c_442_n 0.00392729f $X=2.195 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_224 N_A_27_115#_c_261_n N_Y_c_442_n 0.00250559f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.59
cc_225 N_A_27_115#_c_262_n N_Y_c_442_n 0.021445f $X=2.55 $Y=2.885 $X2=2.41
+ $Y2=2.59
cc_226 N_A_27_115#_c_315_n N_Y_c_442_n 0.00392729f $X=2.625 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_227 N_A_27_115#_c_274_n N_Y_c_442_n 0.00361281f $X=3.055 $Y=2.81 $X2=2.41
+ $Y2=2.59
cc_228 N_A_27_115#_M1013_g N_Y_c_443_n 0.00231637f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=0.825
cc_229 N_A_27_115#_c_275_n N_Y_c_443_n 0.00280419f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=0.825
cc_230 N_A_27_115#_M1015_g N_Y_c_443_n 0.00231637f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=0.825
cc_231 N_A_27_115#_c_274_n N_Y_c_447_n 0.00721971f $X=3.055 $Y=2.81 $X2=3.27
+ $Y2=2.59
cc_232 N_A_27_115#_c_321_n N_Y_c_447_n 0.00392729f $X=3.055 $Y=2.96 $X2=3.27
+ $Y2=2.59
cc_233 N_A_27_115#_c_275_n N_Y_c_447_n 0.00250559f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=2.59
cc_234 N_A_27_115#_c_276_n N_Y_c_447_n 0.0206674f $X=3.41 $Y=2.885 $X2=3.27
+ $Y2=2.59
cc_235 N_A_27_115#_c_326_n N_Y_c_447_n 0.00392729f $X=3.485 $Y=2.96 $X2=3.27
+ $Y2=2.59
cc_236 N_A_27_115#_M1000_g N_Y_c_448_n 0.00554705f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_237 N_A_27_115#_M1009_g N_Y_c_448_n 0.00259902f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_238 N_A_27_115#_c_296_n N_Y_c_448_n 0.00238892f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=1.595
cc_239 N_A_27_115#_c_247_n N_Y_c_451_n 0.00638728f $X=1.335 $Y=2.81 $X2=1.55
+ $Y2=2.475
cc_240 N_A_27_115#_c_248_n N_Y_c_451_n 0.00186325f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.475
cc_241 N_A_27_115#_c_249_n N_Y_c_451_n 0.00140336f $X=1.69 $Y=1.845 $X2=1.55
+ $Y2=2.475
cc_242 N_A_27_115#_c_281_n N_Y_c_451_n 0.00144278f $X=1.395 $Y=1.845 $X2=1.55
+ $Y2=2.475
cc_243 N_A_27_115#_c_296_n N_Y_c_451_n 0.00194461f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=2.475
cc_244 N_A_27_115#_M1000_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_245 N_A_27_115#_c_247_n Y 0.00874077f $X=1.335 $Y=2.81 $X2=1.555 $Y2=2.22
cc_246 N_A_27_115#_c_249_n Y 0.00840707f $X=1.69 $Y=1.845 $X2=1.555 $Y2=2.22
cc_247 N_A_27_115#_M1009_g Y 0.00251111f $X=1.765 $Y=1.075 $X2=1.555 $Y2=2.22
cc_248 N_A_27_115#_c_281_n Y 0.00487273f $X=1.395 $Y=1.845 $X2=1.555 $Y2=2.22
cc_249 N_A_27_115#_c_296_n Y 0.0132141f $X=1.395 $Y=1.935 $X2=1.555 $Y2=2.22
cc_250 N_A_27_115#_M1009_g N_Y_c_453_n 0.0130095f $X=1.765 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_251 N_A_27_115#_c_254_n N_Y_c_453_n 0.00213861f $X=2.12 $Y=1.845 $X2=2.265
+ $Y2=1.48
cc_252 N_A_27_115#_M1010_g N_Y_c_453_n 0.0130095f $X=2.195 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_253 N_A_27_115#_c_283_n N_Y_c_455_n 0.0121767f $X=1.765 $Y=1.845 $X2=2.265
+ $Y2=2.59
cc_254 N_A_27_115#_c_284_n N_Y_c_455_n 0.0158479f $X=1.765 $Y=2.885 $X2=2.265
+ $Y2=2.59
cc_255 N_A_27_115#_M1010_g N_Y_c_456_n 0.00251111f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_256 N_A_27_115#_c_261_n N_Y_c_456_n 0.0177725f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.475
cc_257 N_A_27_115#_M1012_g N_Y_c_456_n 0.00251111f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_258 N_A_27_115#_c_274_n N_Y_c_456_n 0.00843025f $X=3.055 $Y=2.81 $X2=2.41
+ $Y2=2.475
cc_259 N_A_27_115#_M1012_g N_Y_c_457_n 0.0130095f $X=2.625 $Y=1.075 $X2=3.125
+ $Y2=1.48
cc_260 N_A_27_115#_c_267_n N_Y_c_457_n 0.00213861f $X=2.98 $Y=1.845 $X2=3.125
+ $Y2=1.48
cc_261 N_A_27_115#_M1013_g N_Y_c_457_n 0.0136594f $X=3.055 $Y=1.075 $X2=3.125
+ $Y2=1.48
cc_262 N_A_27_115#_M1010_g N_Y_c_459_n 0.00259902f $X=2.195 $Y=1.075 $X2=2.555
+ $Y2=1.48
cc_263 N_A_27_115#_M1012_g N_Y_c_459_n 0.00259902f $X=2.625 $Y=1.075 $X2=2.555
+ $Y2=1.48
cc_264 N_A_27_115#_c_274_n N_Y_c_462_n 0.0155956f $X=3.055 $Y=2.81 $X2=3.125
+ $Y2=2.59
cc_265 N_A_27_115#_c_287_n N_Y_c_462_n 0.00894336f $X=2.625 $Y=1.845 $X2=3.125
+ $Y2=2.59
cc_266 N_A_27_115#_c_288_n N_Y_c_462_n 0.00903839f $X=2.625 $Y=2.885 $X2=3.125
+ $Y2=2.59
cc_267 N_A_27_115#_c_261_n N_Y_c_463_n 0.00140336f $X=2.55 $Y=1.845 $X2=2.555
+ $Y2=2.59
cc_268 N_A_27_115#_c_274_n N_Y_c_463_n 0.0012308f $X=3.055 $Y=2.81 $X2=2.555
+ $Y2=2.59
cc_269 N_A_27_115#_c_285_n N_Y_c_463_n 0.00140336f $X=2.195 $Y=1.845 $X2=2.555
+ $Y2=2.59
cc_270 N_A_27_115#_c_286_n N_Y_c_463_n 0.00372651f $X=2.195 $Y=2.885 $X2=2.555
+ $Y2=2.59
cc_271 N_A_27_115#_M1013_g N_Y_c_464_n 0.00262362f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_272 N_A_27_115#_M1015_g N_Y_c_464_n 0.00939545f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_273 N_A_27_115#_M1013_g N_Y_c_467_n 0.00251111f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=2.475
cc_274 N_A_27_115#_c_274_n N_Y_c_467_n 0.0163934f $X=3.055 $Y=2.81 $X2=3.27
+ $Y2=2.475
cc_275 N_A_27_115#_c_275_n N_Y_c_467_n 0.0196907f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=2.475
cc_276 N_A_27_115#_c_276_n N_Y_c_467_n 0.00357274f $X=3.41 $Y=2.885 $X2=3.27
+ $Y2=2.475
cc_277 N_A_27_115#_M1015_g N_Y_c_467_n 0.00251111f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=2.475
