* File: sky130_osu_sc_15T_hs__tnbufi_l.pex.spice
* Created: Fri Nov 12 14:33:55 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%GND 1 17 19 26 35 38
r31 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r32 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r33 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r34 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r35 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r36 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r37 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r38 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r39 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%VDD 1 13 15 21 25 29 32
r22 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r23 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r24 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r25 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397 $X2=1.02
+ $Y2=5.397
r26 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r27 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.225
r28 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r29 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r30 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r31 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r32 1 21 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.565 $X2=0.69 $Y2=4.225
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%A_27_115# 1 3 11 16 20 24 26 28 31
r43 27 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.915
+ $X2=0.26 $Y2=1.915
r44 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=1.915
+ $X2=0.69 $Y2=1.915
r45 26 27 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.915
+ $X2=0.345 $Y2=1.915
r46 22 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2 $X2=0.26
+ $Y2=1.915
r47 22 24 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=0.26 $Y=2 $X2=0.26
+ $Y2=4.225
r48 18 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.83 $X2=0.26
+ $Y2=1.915
r49 18 20 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.26 $Y=1.83
+ $X2=0.26 $Y2=0.74
r50 14 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.915 $X2=0.69 $Y2=1.915
r51 14 16 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=1.915
+ $X2=0.905 $Y2=1.915
r52 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.75
+ $X2=0.905 $Y2=1.915
r53 9 11 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.905 $Y=1.75 $X2=0.905
+ $Y2=0.85
r54 3 24 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.225
r55 1 20 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%OE 5 7 9 13 17 22 28
r46 25 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.7 $X2=0.69
+ $Y2=2.7
r47 22 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.69 $Y=2.505
+ $X2=0.69 $Y2=2.7
r48 20 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.505 $X2=0.69 $Y2=2.505
r49 15 17 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.475 $Y2=1.465
r50 7 20 49.2914 $w=4.58e-07 $l=4.23124e-07 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.587 $Y2=2.505
r51 7 13 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=4.195
r52 7 9 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=4.195
r53 3 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.475 $Y2=1.465
r54 3 5 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.475 $Y2=0.85
r55 1 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=1.54 $X2=0.27
+ $Y2=1.465
r56 1 7 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.54 $X2=0.27
+ $Y2=2.6
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%A 3 7 10 15 20 23
r47 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.83
+ $X2=1.325 $Y2=1.83
r48 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=3.07
+ $X2=1.14 $Y2=3.07
r49 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.915
+ $X2=1.14 $Y2=1.83
r50 13 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=1.915
+ $X2=1.14 $Y2=3.07
r51 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.83 $X2=1.325 $Y2=1.83
r52 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.83
+ $X2=1.325 $Y2=1.995
r53 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.83
+ $X2=1.325 $Y2=1.665
r54 7 12 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=1.265 $Y=4.195
+ $X2=1.265 $Y2=1.995
r55 3 11 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.265 $Y=0.85
+ $X2=1.265 $Y2=1.665
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%Y 1 3 10 16 24 27 30
r31 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.215
+ $X2=1.48 $Y2=2.33
r32 22 24 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.215
+ $X2=1.48 $Y2=1.56
r33 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.335
+ $X2=1.48 $Y2=1.22
r34 21 24 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.335
+ $X2=1.48 $Y2=1.56
r35 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.33
+ $X2=1.48 $Y2=2.33
r36 16 19 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=1.48 $Y=2.33
+ $X2=1.48 $Y2=4.225
r37 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.22
+ $X2=1.48 $Y2=1.22
r38 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.48 $Y=0.74
+ $X2=1.48 $Y2=1.22
r39 3 19 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=3.565 $X2=1.48 $Y2=4.225
r40 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.74
.ends

