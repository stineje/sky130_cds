* File: sky130_osu_sc_15T_ls__aoi21_l.spice
* Created: Fri Nov 12 14:54:25 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__aoi21_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__aoi21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A0_M1003_g N_GND_M1003_s N_GND_M1003_b NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A1_M1002_g A_110_115# N_GND_M1003_b NSHORT L=0.15 W=0.74
+ AD=0.138075 AS=0.0777 PD=1.26857 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75000.6 SB=75000.5 A=0.111 P=1.78 MULT=1
MM1005 N_GND_M1005_d N_B0_M1005_g N_Y_M1002_d N_GND_M1003_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0970254 PD=1.57 PS=0.891429 NRD=0 NRS=14.412 M=1 R=3.46667
+ SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_VDD_M1000_d N_A0_M1000_g N_A_27_565#_M1000_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1004 N_A_27_565#_M1004_d N_A1_M1004_g N_VDD_M1000_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1001 N_Y_M1001_d N_B0_M1001_g N_A_27_565#_M1004_d N_VDD_M1000_b PHIGHVT L=0.15
+ W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=5.64925 P=9.73
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__aoi21_l.pxi.spice"
*
.ends
*
*
