* File: sky130_osu_sc_12T_hs__dff_1.pxi.spice
* Created: Fri Nov 12 15:08:56 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%GND N_GND_M1008_d N_GND_M1013_d N_GND_M1000_d
+ N_GND_M1009_s N_GND_M1010_d N_GND_M1008_b N_GND_c_2_p N_GND_c_3_p N_GND_c_16_p
+ N_GND_c_59_p N_GND_c_35_p N_GND_c_39_p N_GND_c_40_p N_GND_c_41_p N_GND_c_117_p
+ N_GND_c_118_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_HS__DFF_1%GND
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%VDD N_VDD_M1022_d N_VDD_M1004_d N_VDD_M1016_d
+ N_VDD_M1023_s N_VDD_M1024_d N_VDD_M1022_b N_VDD_c_184_p N_VDD_c_185_p
+ N_VDD_c_194_p N_VDD_c_220_p N_VDD_c_205_p N_VDD_c_209_p N_VDD_c_210_p
+ N_VDD_c_211_p N_VDD_c_251_p N_VDD_c_252_p N_VDD_c_273_p VDD N_VDD_c_186_p
+ PM_SKY130_OSU_SC_12T_HS__DFF_1%VDD
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%A_75_248# N_A_75_248#_M1025_d
+ N_A_75_248#_M1014_d N_A_75_248#_M1008_g N_A_75_248#_M1022_g
+ N_A_75_248#_c_284_n N_A_75_248#_c_288_n N_A_75_248#_c_289_n
+ N_A_75_248#_c_290_n N_A_75_248#_c_306_n N_A_75_248#_c_291_n
+ N_A_75_248#_c_293_n N_A_75_248#_c_307_n N_A_75_248#_c_309_n
+ N_A_75_248#_c_295_n N_A_75_248#_c_311_n N_A_75_248#_c_296_n
+ N_A_75_248#_c_297_n N_A_75_248#_c_298_n
+ PM_SKY130_OSU_SC_12T_HS__DFF_1%A_75_248#
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%D N_D_M1007_g N_D_M1021_g N_D_c_378_n
+ N_D_c_379_n D PM_SKY130_OSU_SC_12T_HS__DFF_1%D
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%CK N_CK_M1014_g N_CK_M1020_g N_CK_M1012_g
+ N_CK_M1019_g N_CK_M1001_g N_CK_c_416_n N_CK_M1017_g N_CK_c_417_n N_CK_c_418_n
+ N_CK_c_419_n N_CK_c_420_n N_CK_c_423_n N_CK_c_424_n N_CK_c_427_n N_CK_c_428_n
+ N_CK_c_433_n N_CK_c_434_n N_CK_c_435_n N_CK_c_436_n N_CK_c_437_n N_CK_c_438_n
+ N_CK_c_439_n N_CK_c_440_n N_CK_c_441_n N_CK_c_442_n N_CK_c_443_n N_CK_c_444_n
+ N_CK_c_445_n CK PM_SKY130_OSU_SC_12T_HS__DFF_1%CK
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%A_32_115# N_A_32_115#_M1008_s
+ N_A_32_115#_M1022_s N_A_32_115#_M1013_g N_A_32_115#_M1004_g
+ N_A_32_115#_c_648_n N_A_32_115#_c_650_n N_A_32_115#_c_651_n
+ N_A_32_115#_c_652_n N_A_32_115#_M1015_g N_A_32_115#_M1006_g
+ N_A_32_115#_c_657_n N_A_32_115#_c_658_n N_A_32_115#_c_680_n
+ N_A_32_115#_c_661_n N_A_32_115#_c_662_n N_A_32_115#_c_685_n
+ N_A_32_115#_c_663_n N_A_32_115#_c_665_n N_A_32_115#_c_667_n
+ N_A_32_115#_c_668_n PM_SKY130_OSU_SC_12T_HS__DFF_1%A_32_115#
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%A_243_89# N_A_243_89#_M1001_d
+ N_A_243_89#_M1017_d N_A_243_89#_c_759_n N_A_243_89#_M1025_g
+ N_A_243_89#_c_762_n N_A_243_89#_c_763_n N_A_243_89#_c_764_n
+ N_A_243_89#_M1011_g N_A_243_89#_c_766_n N_A_243_89#_M1003_g
+ N_A_243_89#_c_768_n N_A_243_89#_M1005_g N_A_243_89#_c_772_n
+ N_A_243_89#_c_773_n N_A_243_89#_c_774_n N_A_243_89#_c_775_n
+ N_A_243_89#_c_776_n N_A_243_89#_c_777_n N_A_243_89#_c_792_n
+ N_A_243_89#_c_781_n N_A_243_89#_c_797_n N_A_243_89#_c_782_n
+ N_A_243_89#_c_783_n N_A_243_89#_c_784_n N_A_243_89#_c_785_n
+ PM_SKY130_OSU_SC_12T_HS__DFF_1%A_243_89#
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%A_785_89# N_A_785_89#_M1009_d
+ N_A_785_89#_M1023_d N_A_785_89#_M1000_g N_A_785_89#_M1016_g
+ N_A_785_89#_c_957_n N_A_785_89#_M1010_g N_A_785_89#_M1024_g
+ N_A_785_89#_c_962_n N_A_785_89#_c_964_n N_A_785_89#_c_965_n
+ N_A_785_89#_c_966_n N_A_785_89#_c_967_n N_A_785_89#_c_968_n
+ N_A_785_89#_c_971_n N_A_785_89#_c_972_n N_A_785_89#_c_973_n
+ N_A_785_89#_c_974_n N_A_785_89#_c_975_n N_A_785_89#_c_976_n
+ N_A_785_89#_c_977_n N_A_785_89#_c_978_n N_A_785_89#_c_979_n
+ PM_SKY130_OSU_SC_12T_HS__DFF_1%A_785_89#
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%A_623_115# N_A_623_115#_M1012_d
+ N_A_623_115#_M1003_d N_A_623_115#_c_1117_n N_A_623_115#_M1009_g
+ N_A_623_115#_M1023_g N_A_623_115#_c_1122_n N_A_623_115#_c_1124_n
+ N_A_623_115#_c_1154_n N_A_623_115#_c_1184_n N_A_623_115#_c_1143_n
+ N_A_623_115#_c_1125_n N_A_623_115#_c_1126_n N_A_623_115#_c_1129_n
+ N_A_623_115#_c_1131_n N_A_623_115#_c_1132_n N_A_623_115#_c_1133_n
+ N_A_623_115#_c_1135_n N_A_623_115#_c_1136_n
+ PM_SKY130_OSU_SC_12T_HS__DFF_1%A_623_115#
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%ON N_ON_M1010_s N_ON_M1024_s N_ON_M1002_g
+ N_ON_M1018_g N_ON_c_1244_n N_ON_c_1245_n N_ON_c_1248_n N_ON_c_1249_n
+ N_ON_c_1250_n N_ON_c_1252_n N_ON_c_1253_n N_ON_c_1254_n N_ON_c_1255_n
+ N_ON_c_1256_n ON PM_SKY130_OSU_SC_12T_HS__DFF_1%ON
x_PM_SKY130_OSU_SC_12T_HS__DFF_1%Q N_Q_M1002_d N_Q_M1018_d N_Q_c_1320_n
+ N_Q_c_1326_n N_Q_c_1322_n N_Q_c_1323_n N_Q_c_1330_n N_Q_c_1324_n Q
+ PM_SKY130_OSU_SC_12T_HS__DFF_1%Q
cc_1 N_GND_M1008_b N_A_75_248#_c_284_n 0.0206783f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=1.24
cc_2 N_GND_c_2_p N_A_75_248#_c_284_n 0.00606474f $X=0.63 $Y=0.152 $X2=0.475
+ $Y2=1.24
cc_3 N_GND_c_3_p N_A_75_248#_c_284_n 0.00308284f $X=0.715 $Y=0.755 $X2=0.475
+ $Y2=1.24
cc_4 N_GND_c_4_p N_A_75_248#_c_284_n 0.00468827f $X=6.46 $Y=0.19 $X2=0.475
+ $Y2=1.24
cc_5 N_GND_M1008_b N_A_75_248#_c_288_n 0.0143449f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=1.39
cc_6 N_GND_M1008_b N_A_75_248#_c_289_n 0.0223136f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.285
cc_7 N_GND_M1008_b N_A_75_248#_c_290_n 0.0431517f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.12
cc_8 N_GND_M1008_b N_A_75_248#_c_291_n 0.018477f $X=-0.045 $Y=0 $X2=1.405
+ $Y2=1.285
cc_9 N_GND_c_3_p N_A_75_248#_c_291_n 0.00456782f $X=0.715 $Y=0.755 $X2=1.405
+ $Y2=1.285
cc_10 N_GND_M1008_b N_A_75_248#_c_293_n 0.00315644f $X=-0.045 $Y=0 $X2=0.71
+ $Y2=1.285
cc_11 N_GND_c_3_p N_A_75_248#_c_293_n 0.00460441f $X=0.715 $Y=0.755 $X2=0.71
+ $Y2=1.285
cc_12 N_GND_M1008_b N_A_75_248#_c_295_n 0.00140975f $X=-0.045 $Y=0 $X2=1.49
+ $Y2=1.2
cc_13 N_GND_M1008_b N_A_75_248#_c_296_n 0.00329831f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.285
cc_14 N_GND_M1008_b N_A_75_248#_c_297_n 0.012703f $X=-0.045 $Y=0 $X2=0.567
+ $Y2=2.12
cc_15 N_GND_M1008_b N_A_75_248#_c_298_n 0.00311983f $X=-0.045 $Y=0 $X2=1.49
+ $Y2=0.755
cc_16 N_GND_c_16_p N_A_75_248#_c_298_n 0.0145844f $X=2.38 $Y=0.152 $X2=1.49
+ $Y2=0.755
cc_17 N_GND_c_4_p N_A_75_248#_c_298_n 0.0098977f $X=6.46 $Y=0.19 $X2=1.49
+ $Y2=0.755
cc_18 N_GND_M1008_b N_D_M1007_g 0.0319343f $X=-0.045 $Y=0 $X2=0.93 $Y2=0.85
cc_19 N_GND_c_3_p N_D_M1007_g 0.00308284f $X=0.715 $Y=0.755 $X2=0.93 $Y2=0.85
cc_20 N_GND_c_16_p N_D_M1007_g 0.00606474f $X=2.38 $Y=0.152 $X2=0.93 $Y2=0.85
cc_21 N_GND_c_4_p N_D_M1007_g 0.00468827f $X=6.46 $Y=0.19 $X2=0.93 $Y2=0.85
cc_22 N_GND_M1008_b N_D_M1021_g 0.0297434f $X=-0.045 $Y=0 $X2=0.93 $Y2=3.235
cc_23 N_GND_M1008_b N_D_c_378_n 0.0271295f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.74
cc_24 N_GND_M1008_b N_D_c_379_n 0.00311208f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.74
cc_25 N_GND_M1008_b D 0.00874486f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.74
cc_26 N_GND_M1008_b N_CK_c_416_n 0.0307739f $X=-0.045 $Y=0 $X2=4.43 $Y2=2.45
cc_27 N_GND_M1008_b N_CK_c_417_n 0.0449017f $X=-0.045 $Y=0 $X2=4.485 $Y2=2.12
cc_28 N_GND_M1008_b N_CK_c_418_n 0.0247685f $X=-0.045 $Y=0 $X2=1.38 $Y2=2.285
cc_29 N_GND_M1008_b N_CK_c_419_n 0.0254952f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.4
cc_30 N_GND_M1008_b N_CK_c_420_n 0.017381f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.235
cc_31 N_GND_c_16_p N_CK_c_420_n 0.00606474f $X=2.38 $Y=0.152 $X2=1.83 $Y2=1.235
cc_32 N_GND_c_4_p N_CK_c_420_n 0.00468827f $X=6.46 $Y=0.19 $X2=1.83 $Y2=1.235
cc_33 N_GND_M1008_b N_CK_c_423_n 0.0268494f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.4
cc_34 N_GND_M1008_b N_CK_c_424_n 0.0174883f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.235
cc_35 N_GND_c_35_p N_CK_c_424_n 0.00606474f $X=4.13 $Y=0.152 $X2=3.1 $Y2=1.235
cc_36 N_GND_c_4_p N_CK_c_424_n 0.00468827f $X=6.46 $Y=0.19 $X2=3.1 $Y2=1.235
cc_37 N_GND_M1008_b N_CK_c_427_n 0.0223817f $X=-0.045 $Y=0 $X2=3.55 $Y2=2.285
cc_38 N_GND_M1008_b N_CK_c_428_n 0.0166942f $X=-0.045 $Y=0 $X2=4.457 $Y2=1.205
cc_39 N_GND_c_39_p N_CK_c_428_n 0.00308284f $X=4.215 $Y=0.755 $X2=4.457
+ $Y2=1.205
cc_40 N_GND_c_40_p N_CK_c_428_n 0.00606474f $X=5.08 $Y=0.152 $X2=4.457 $Y2=1.205
cc_41 N_GND_c_41_p N_CK_c_428_n 0.00365683f $X=5.165 $Y=0.755 $X2=4.457
+ $Y2=1.205
cc_42 N_GND_c_4_p N_CK_c_428_n 0.00468827f $X=6.46 $Y=0.19 $X2=4.457 $Y2=1.205
cc_43 N_GND_M1008_b N_CK_c_433_n 0.0140293f $X=-0.045 $Y=0 $X2=4.457 $Y2=1.355
cc_44 N_GND_M1008_b N_CK_c_434_n 0.00530209f $X=-0.045 $Y=0 $X2=1.745 $Y2=2.11
cc_45 N_GND_M1008_b N_CK_c_435_n 0.00995082f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.4
cc_46 N_GND_M1008_b N_CK_c_436_n 0.00850752f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.4
cc_47 N_GND_M1008_b N_CK_c_437_n 0.00428249f $X=-0.045 $Y=0 $X2=3.465 $Y2=2.11
cc_48 N_GND_M1008_b N_CK_c_438_n 5.00459e-19 $X=-0.045 $Y=0 $X2=3.185 $Y2=2.11
cc_49 N_GND_M1008_b N_CK_c_439_n 7.09602e-19 $X=-0.045 $Y=0 $X2=4.575 $Y2=2.11
cc_50 N_GND_M1008_b N_CK_c_440_n 0.00290411f $X=-0.045 $Y=0 $X2=1.35 $Y2=2.11
cc_51 N_GND_M1008_b N_CK_c_441_n 0.00150017f $X=-0.045 $Y=0 $X2=3.58 $Y2=2.11
cc_52 N_GND_M1008_b N_CK_c_442_n 0.0328858f $X=-0.045 $Y=0 $X2=3.435 $Y2=2.11
cc_53 N_GND_M1008_b N_CK_c_443_n 0.00558706f $X=-0.045 $Y=0 $X2=1.495 $Y2=2.11
cc_54 N_GND_M1008_b N_CK_c_444_n 0.0134637f $X=-0.045 $Y=0 $X2=4.43 $Y2=2.11
cc_55 N_GND_M1008_b N_CK_c_445_n 0.0021042f $X=-0.045 $Y=0 $X2=3.725 $Y2=2.11
cc_56 N_GND_M1008_b CK 0.00144846f $X=-0.045 $Y=0 $X2=4.575 $Y2=2.11
cc_57 N_GND_M1008_b N_A_32_115#_M1013_g 0.0171592f $X=-0.045 $Y=0 $X2=2.25
+ $Y2=0.85
cc_58 N_GND_c_16_p N_A_32_115#_M1013_g 0.00606474f $X=2.38 $Y=0.152 $X2=2.25
+ $Y2=0.85
cc_59 N_GND_c_59_p N_A_32_115#_M1013_g 0.00308284f $X=2.465 $Y=0.74 $X2=2.25
+ $Y2=0.85
cc_60 N_GND_c_4_p N_A_32_115#_M1013_g 0.00468827f $X=6.46 $Y=0.19 $X2=2.25
+ $Y2=0.85
cc_61 N_GND_M1008_b N_A_32_115#_c_648_n 0.0240502f $X=-0.045 $Y=0 $X2=2.605
+ $Y2=1.4
cc_62 N_GND_c_59_p N_A_32_115#_c_648_n 9.75298e-19 $X=2.465 $Y=0.74 $X2=2.605
+ $Y2=1.4
cc_63 N_GND_M1008_b N_A_32_115#_c_650_n 0.0105855f $X=-0.045 $Y=0 $X2=2.325
+ $Y2=1.4
cc_64 N_GND_M1008_b N_A_32_115#_c_651_n 0.022671f $X=-0.045 $Y=0 $X2=2.605
+ $Y2=2.285
cc_65 N_GND_M1008_b N_A_32_115#_c_652_n 0.0103324f $X=-0.045 $Y=0 $X2=2.325
+ $Y2=2.285
cc_66 N_GND_M1008_b N_A_32_115#_M1015_g 0.0171447f $X=-0.045 $Y=0 $X2=2.68
+ $Y2=0.85
cc_67 N_GND_c_59_p N_A_32_115#_M1015_g 0.00308284f $X=2.465 $Y=0.74 $X2=2.68
+ $Y2=0.85
cc_68 N_GND_c_35_p N_A_32_115#_M1015_g 0.00606474f $X=4.13 $Y=0.152 $X2=2.68
+ $Y2=0.85
cc_69 N_GND_c_4_p N_A_32_115#_M1015_g 0.00468827f $X=6.46 $Y=0.19 $X2=2.68
+ $Y2=0.85
cc_70 N_GND_M1008_b N_A_32_115#_c_657_n 0.0456538f $X=-0.045 $Y=0 $X2=0.17
+ $Y2=2.695
cc_71 N_GND_M1008_b N_A_32_115#_c_658_n 0.0046518f $X=-0.045 $Y=0 $X2=0.285
+ $Y2=0.755
cc_72 N_GND_c_2_p N_A_32_115#_c_658_n 0.00729833f $X=0.63 $Y=0.152 $X2=0.285
+ $Y2=0.755
cc_73 N_GND_c_4_p N_A_32_115#_c_658_n 0.00474439f $X=6.46 $Y=0.19 $X2=0.285
+ $Y2=0.755
cc_74 N_GND_M1008_b N_A_32_115#_c_661_n 0.00822335f $X=-0.045 $Y=0 $X2=2.42
+ $Y2=2.285
cc_75 N_GND_M1008_b N_A_32_115#_c_662_n 0.0203007f $X=-0.045 $Y=0 $X2=0.285
+ $Y2=1.37
cc_76 N_GND_M1008_b N_A_32_115#_c_663_n 0.00385085f $X=-0.045 $Y=0 $X2=2.42
+ $Y2=1.4
cc_77 N_GND_c_59_p N_A_32_115#_c_663_n 0.00620301f $X=2.465 $Y=0.74 $X2=2.42
+ $Y2=1.4
cc_78 N_GND_M1008_b N_A_32_115#_c_665_n 0.0225524f $X=-0.045 $Y=0 $X2=2.185
+ $Y2=1.37
cc_79 N_GND_c_3_p N_A_32_115#_c_665_n 0.00118122f $X=0.715 $Y=0.755 $X2=2.185
+ $Y2=1.37
cc_80 N_GND_M1008_b N_A_32_115#_c_667_n 0.00468924f $X=-0.045 $Y=0 $X2=0.43
+ $Y2=1.37
cc_81 N_GND_M1008_b N_A_32_115#_c_668_n 3.72162e-19 $X=-0.045 $Y=0 $X2=2.33
+ $Y2=1.37
cc_82 N_GND_c_59_p N_A_32_115#_c_668_n 7.4089e-19 $X=2.465 $Y=0.74 $X2=2.33
+ $Y2=1.37
cc_83 N_GND_M1008_b N_A_243_89#_c_759_n 0.0156145f $X=-0.045 $Y=0 $X2=1.29
+ $Y2=1.205
cc_84 N_GND_c_16_p N_A_243_89#_c_759_n 0.00606474f $X=2.38 $Y=0.152 $X2=1.29
+ $Y2=1.205
cc_85 N_GND_c_4_p N_A_243_89#_c_759_n 0.00468827f $X=6.46 $Y=0.19 $X2=1.29
+ $Y2=1.205
cc_86 N_GND_M1008_b N_A_243_89#_c_762_n 0.0217401f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.775
cc_87 N_GND_M1008_b N_A_243_89#_c_763_n 0.0182441f $X=-0.045 $Y=0 $X2=1.815
+ $Y2=1.85
cc_88 N_GND_M1008_b N_A_243_89#_c_764_n 0.00766736f $X=-0.045 $Y=0 $X2=1.485
+ $Y2=1.85
cc_89 N_GND_M1008_b N_A_243_89#_M1011_g 0.0302127f $X=-0.045 $Y=0 $X2=1.89
+ $Y2=3.235
cc_90 N_GND_M1008_b N_A_243_89#_c_766_n 0.0552247f $X=-0.045 $Y=0 $X2=2.965
+ $Y2=1.85
cc_91 N_GND_M1008_b N_A_243_89#_M1003_g 0.0297952f $X=-0.045 $Y=0 $X2=3.04
+ $Y2=3.235
cc_92 N_GND_M1008_b N_A_243_89#_c_768_n 0.0182441f $X=-0.045 $Y=0 $X2=3.445
+ $Y2=1.85
cc_93 N_GND_M1008_b N_A_243_89#_M1005_g 0.0335991f $X=-0.045 $Y=0 $X2=3.64
+ $Y2=0.85
cc_94 N_GND_c_35_p N_A_243_89#_M1005_g 0.00606474f $X=4.13 $Y=0.152 $X2=3.64
+ $Y2=0.85
cc_95 N_GND_c_4_p N_A_243_89#_M1005_g 0.00468827f $X=6.46 $Y=0.19 $X2=3.64
+ $Y2=0.85
cc_96 N_GND_M1008_b N_A_243_89#_c_772_n 0.0143258f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.28
cc_97 N_GND_M1008_b N_A_243_89#_c_773_n 0.00426513f $X=-0.045 $Y=0 $X2=1.89
+ $Y2=1.85
cc_98 N_GND_M1008_b N_A_243_89#_c_774_n 0.00426513f $X=-0.045 $Y=0 $X2=3.04
+ $Y2=1.85
cc_99 N_GND_M1008_b N_A_243_89#_c_775_n 0.0281466f $X=-0.045 $Y=0 $X2=3.58
+ $Y2=1.74
cc_100 N_GND_M1008_b N_A_243_89#_c_776_n 0.00218483f $X=-0.045 $Y=0 $X2=3.58
+ $Y2=1.74
cc_101 N_GND_M1008_b N_A_243_89#_c_777_n 0.0151508f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=0.755
cc_102 N_GND_c_40_p N_A_243_89#_c_777_n 0.00749582f $X=5.08 $Y=0.152 $X2=4.645
+ $Y2=0.755
cc_103 N_GND_c_41_p N_A_243_89#_c_777_n 0.0153786f $X=5.165 $Y=0.755 $X2=4.645
+ $Y2=0.755
cc_104 N_GND_c_4_p N_A_243_89#_c_777_n 0.00476261f $X=6.46 $Y=0.19 $X2=4.645
+ $Y2=0.755
cc_105 N_GND_M1008_b N_A_243_89#_c_781_n 0.0115392f $X=-0.045 $Y=0 $X2=4.915
+ $Y2=2.62
cc_106 N_GND_M1008_b N_A_243_89#_c_782_n 0.0110805f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=1.74
cc_107 N_GND_M1008_b N_A_243_89#_c_783_n 0.00199631f $X=-0.045 $Y=0 $X2=3.725
+ $Y2=1.725
cc_108 N_GND_M1008_b N_A_243_89#_c_784_n 0.00257437f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=1.74
cc_109 N_GND_M1008_b N_A_243_89#_c_785_n 0.00682657f $X=-0.045 $Y=0 $X2=4.5
+ $Y2=1.74
cc_110 N_GND_M1008_b N_A_785_89#_M1000_g 0.032189f $X=-0.045 $Y=0 $X2=4 $Y2=0.85
cc_111 N_GND_c_35_p N_A_785_89#_M1000_g 0.00606474f $X=4.13 $Y=0.152 $X2=4
+ $Y2=0.85
cc_112 N_GND_c_39_p N_A_785_89#_M1000_g 0.00308284f $X=4.215 $Y=0.755 $X2=4
+ $Y2=0.85
cc_113 N_GND_c_4_p N_A_785_89#_M1000_g 0.00468827f $X=6.46 $Y=0.19 $X2=4
+ $Y2=0.85
cc_114 N_GND_M1008_b N_A_785_89#_M1016_g 0.0287643f $X=-0.045 $Y=0 $X2=4
+ $Y2=3.235
cc_115 N_GND_M1008_b N_A_785_89#_c_957_n 0.0524798f $X=-0.045 $Y=0 $X2=6.28
+ $Y2=1.905
cc_116 N_GND_M1008_b N_A_785_89#_M1010_g 0.0225944f $X=-0.045 $Y=0 $X2=6.33
+ $Y2=0.85
cc_117 N_GND_c_117_p N_A_785_89#_M1010_g 0.00606474f $X=6.46 $Y=0.152 $X2=6.33
+ $Y2=0.85
cc_118 N_GND_c_118_p N_A_785_89#_M1010_g 0.00308284f $X=6.545 $Y=0.74 $X2=6.33
+ $Y2=0.85
cc_119 N_GND_c_4_p N_A_785_89#_M1010_g 0.00468827f $X=6.46 $Y=0.19 $X2=6.33
+ $Y2=0.85
cc_120 N_GND_M1008_b N_A_785_89#_c_962_n 0.0263051f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=1.74
cc_121 N_GND_c_39_p N_A_785_89#_c_962_n 0.00144867f $X=4.215 $Y=0.755 $X2=4.06
+ $Y2=1.74
cc_122 N_GND_M1008_b N_A_785_89#_c_964_n 0.026659f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=2.36
cc_123 N_GND_M1008_b N_A_785_89#_c_965_n 0.00533488f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=2.49
cc_124 N_GND_M1008_b N_A_785_89#_c_966_n 8.68018e-19 $X=-0.045 $Y=0 $X2=4.062
+ $Y2=1.812
cc_125 N_GND_M1008_b N_A_785_89#_c_967_n 0.00374026f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=2.48
cc_126 N_GND_M1008_b N_A_785_89#_c_968_n 0.0137272f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=0.755
cc_127 N_GND_c_117_p N_A_785_89#_c_968_n 0.0074445f $X=6.46 $Y=0.152 $X2=5.595
+ $Y2=0.755
cc_128 N_GND_c_4_p N_A_785_89#_c_968_n 0.00476261f $X=6.46 $Y=0.19 $X2=5.595
+ $Y2=0.755
cc_129 N_GND_M1008_b N_A_785_89#_c_971_n 0.0135339f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=2.955
cc_130 N_GND_M1008_b N_A_785_89#_c_972_n 0.012202f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=1.74
cc_131 N_GND_M1008_b N_A_785_89#_c_973_n 0.00243106f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=1.74
cc_132 N_GND_M1008_b N_A_785_89#_c_974_n 0.00259135f $X=-0.045 $Y=0 $X2=4.935
+ $Y2=2.48
cc_133 N_GND_M1008_b N_A_785_89#_c_975_n 0.00122267f $X=-0.045 $Y=0 $X2=4.205
+ $Y2=2.48
cc_134 N_GND_M1008_b N_A_785_89#_c_976_n 0.0053881f $X=-0.045 $Y=0 $X2=5.007
+ $Y2=2.395
cc_135 N_GND_M1008_b N_A_785_89#_c_977_n 0.0342039f $X=-0.045 $Y=0 $X2=6.08
+ $Y2=1.74
cc_136 N_GND_M1008_b N_A_785_89#_c_978_n 8.85102e-19 $X=-0.045 $Y=0 $X2=5.08
+ $Y2=1.74
cc_137 N_GND_M1008_b N_A_785_89#_c_979_n 0.00114171f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=1.74
cc_138 N_GND_M1008_b N_A_623_115#_c_1117_n 0.0221119f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=1.235
cc_139 N_GND_c_41_p N_A_623_115#_c_1117_n 0.00502587f $X=5.165 $Y=0.755 $X2=5.38
+ $Y2=1.235
cc_140 N_GND_c_117_p N_A_623_115#_c_1117_n 0.00606474f $X=6.46 $Y=0.152 $X2=5.38
+ $Y2=1.235
cc_141 N_GND_c_4_p N_A_623_115#_c_1117_n 0.00468827f $X=6.46 $Y=0.19 $X2=5.38
+ $Y2=1.235
cc_142 N_GND_M1008_b N_A_623_115#_M1023_g 0.0576696f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=3.235
cc_143 N_GND_M1008_b N_A_623_115#_c_1122_n 0.0484026f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=1.4
cc_144 N_GND_c_41_p N_A_623_115#_c_1122_n 0.00372615f $X=5.165 $Y=0.755 $X2=5.38
+ $Y2=1.4
cc_145 N_GND_M1008_b N_A_623_115#_c_1124_n 0.010671f $X=-0.045 $Y=0 $X2=2.76
+ $Y2=1.37
cc_146 N_GND_M1008_b N_A_623_115#_c_1125_n 0.00862295f $X=-0.045 $Y=0 $X2=3.44
+ $Y2=1.34
cc_147 N_GND_M1008_b N_A_623_115#_c_1126_n 0.00312748f $X=-0.045 $Y=0 $X2=3.34
+ $Y2=0.755
cc_148 N_GND_c_35_p N_A_623_115#_c_1126_n 0.0152394f $X=4.13 $Y=0.152 $X2=3.34
+ $Y2=0.755
cc_149 N_GND_c_4_p N_A_623_115#_c_1126_n 0.00994746f $X=6.46 $Y=0.19 $X2=3.34
+ $Y2=0.755
cc_150 N_GND_M1008_b N_A_623_115#_c_1129_n 0.00170347f $X=-0.045 $Y=0 $X2=5.175
+ $Y2=1.37
cc_151 N_GND_c_41_p N_A_623_115#_c_1129_n 0.00509045f $X=5.165 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_152 N_GND_M1008_b N_A_623_115#_c_1131_n 0.00412066f $X=-0.045 $Y=0 $X2=3.295
+ $Y2=1.37
cc_153 N_GND_M1008_b N_A_623_115#_c_1132_n 0.00645439f $X=-0.045 $Y=0 $X2=2.905
+ $Y2=1.37
cc_154 N_GND_M1008_b N_A_623_115#_c_1133_n 0.0298833f $X=-0.045 $Y=0 $X2=5.03
+ $Y2=1.37
cc_155 N_GND_c_39_p N_A_623_115#_c_1133_n 0.00727398f $X=4.215 $Y=0.755 $X2=5.03
+ $Y2=1.37
cc_156 N_GND_M1008_b N_A_623_115#_c_1135_n 0.00473166f $X=-0.045 $Y=0 $X2=3.585
+ $Y2=1.37
cc_157 N_GND_M1008_b N_A_623_115#_c_1136_n 7.10158e-19 $X=-0.045 $Y=0 $X2=5.175
+ $Y2=1.37
cc_158 N_GND_c_41_p N_A_623_115#_c_1136_n 0.00387467f $X=5.165 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_159 N_GND_M1008_b N_ON_M1002_g 0.0597145f $X=-0.045 $Y=0 $X2=6.76 $Y2=0.85
cc_160 N_GND_c_118_p N_ON_M1002_g 0.00308284f $X=6.545 $Y=0.74 $X2=6.76 $Y2=0.85
cc_161 N_GND_c_4_p N_ON_M1002_g 0.00468827f $X=6.46 $Y=0.19 $X2=6.76 $Y2=0.85
cc_162 N_GND_M1008_b N_ON_M1018_g 0.0148936f $X=-0.045 $Y=0 $X2=6.76 $Y2=3.235
cc_163 N_GND_M1008_b N_ON_c_1244_n 0.0285256f $X=-0.045 $Y=0 $X2=6.7 $Y2=2.015
cc_164 N_GND_M1008_b N_ON_c_1245_n 0.00515004f $X=-0.045 $Y=0 $X2=6.115 $Y2=0.74
cc_165 N_GND_c_117_p N_ON_c_1245_n 0.00757793f $X=6.46 $Y=0.152 $X2=6.115
+ $Y2=0.74
cc_166 N_GND_c_4_p N_ON_c_1245_n 0.00476261f $X=6.46 $Y=0.19 $X2=6.115 $Y2=0.74
cc_167 N_GND_M1008_b N_ON_c_1248_n 0.00173247f $X=-0.045 $Y=0 $X2=6.115
+ $Y2=2.195
cc_168 N_GND_M1008_b N_ON_c_1249_n 0.00445021f $X=-0.045 $Y=0 $X2=6.115
+ $Y2=3.615
cc_169 N_GND_M1008_b N_ON_c_1250_n 0.00951514f $X=-0.045 $Y=0 $X2=6.615 $Y2=1.4
cc_170 N_GND_c_118_p N_ON_c_1250_n 0.00738334f $X=6.545 $Y=0.74 $X2=6.615
+ $Y2=1.4
cc_171 N_GND_M1008_b N_ON_c_1252_n 0.0026304f $X=-0.045 $Y=0 $X2=6.2 $Y2=1.4
cc_172 N_GND_M1008_b N_ON_c_1253_n 0.0130744f $X=-0.045 $Y=0 $X2=6.615 $Y2=2.11
cc_173 N_GND_M1008_b N_ON_c_1254_n 0.00154829f $X=-0.045 $Y=0 $X2=6.702
+ $Y2=1.658
cc_174 N_GND_M1008_b N_ON_c_1255_n 5.47532e-19 $X=-0.045 $Y=0 $X2=6.7 $Y2=2.015
cc_175 N_GND_M1008_b N_ON_c_1256_n 5.06249e-19 $X=-0.045 $Y=0 $X2=6.702
+ $Y2=1.745
cc_176 N_GND_M1008_b ON 0.00962953f $X=-0.045 $Y=0 $X2=6.115 $Y2=2.11
cc_177 N_GND_M1008_b N_Q_c_1320_n 0.00885446f $X=-0.045 $Y=0 $X2=6.975 $Y2=0.74
cc_178 N_GND_c_4_p N_Q_c_1320_n 0.00468662f $X=6.46 $Y=0.19 $X2=6.975 $Y2=0.74
cc_179 N_GND_M1008_b N_Q_c_1322_n 0.060171f $X=-0.045 $Y=0 $X2=7.09 $Y2=2.395
cc_180 N_GND_M1008_b N_Q_c_1323_n 0.00345218f $X=-0.045 $Y=0 $X2=7.09 $Y2=2.48
cc_181 N_GND_M1008_b N_Q_c_1324_n 0.0141022f $X=-0.045 $Y=0 $X2=7.09 $Y2=1.07
cc_182 N_GND_M1008_b Q 0.00636397f $X=-0.045 $Y=0 $X2=6.97 $Y2=2.48
cc_183 N_VDD_M1022_b N_A_75_248#_M1022_g 0.0224266f $X=-0.045 $Y=2.425 $X2=0.5
+ $Y2=3.235
cc_184 N_VDD_c_184_p N_A_75_248#_M1022_g 0.00606474f $X=0.63 $Y=4.287 $X2=0.5
+ $Y2=3.235
cc_185 N_VDD_c_185_p N_A_75_248#_M1022_g 0.00337744f $X=0.715 $Y=3.295 $X2=0.5
+ $Y2=3.235
cc_186 N_VDD_c_186_p N_A_75_248#_M1022_g 0.00468827f $X=6.46 $Y=4.25 $X2=0.5
+ $Y2=3.235
cc_187 N_VDD_M1022_b N_A_75_248#_c_289_n 0.00631278f $X=-0.045 $Y=2.425 $X2=0.51
+ $Y2=2.285
cc_188 N_VDD_M1022_b N_A_75_248#_c_306_n 0.00145465f $X=-0.045 $Y=2.425
+ $X2=0.625 $Y2=2.62
cc_189 N_VDD_M1022_d N_A_75_248#_c_307_n 0.00447048f $X=0.575 $Y=2.605 $X2=1.42
+ $Y2=2.705
cc_190 N_VDD_c_185_p N_A_75_248#_c_307_n 0.00499116f $X=0.715 $Y=3.295 $X2=1.42
+ $Y2=2.705
cc_191 N_VDD_M1022_d N_A_75_248#_c_309_n 0.00106276f $X=0.575 $Y=2.605 $X2=0.71
+ $Y2=2.705
cc_192 N_VDD_c_185_p N_A_75_248#_c_309_n 0.00488762f $X=0.715 $Y=3.295 $X2=0.71
+ $Y2=2.705
cc_193 N_VDD_M1022_b N_A_75_248#_c_311_n 0.00313975f $X=-0.045 $Y=2.425 $X2=1.59
+ $Y2=2.955
cc_194 N_VDD_c_194_p N_A_75_248#_c_311_n 0.0149076f $X=2.38 $Y=4.287 $X2=1.59
+ $Y2=2.955
cc_195 N_VDD_c_186_p N_A_75_248#_c_311_n 0.00958198f $X=6.46 $Y=4.25 $X2=1.59
+ $Y2=2.955
cc_196 N_VDD_M1022_b N_A_75_248#_c_296_n 2.34911e-19 $X=-0.045 $Y=2.425 $X2=0.51
+ $Y2=2.285
cc_197 N_VDD_M1022_b N_D_M1021_g 0.0196482f $X=-0.045 $Y=2.425 $X2=0.93
+ $Y2=3.235
cc_198 N_VDD_c_185_p N_D_M1021_g 0.00337744f $X=0.715 $Y=3.295 $X2=0.93
+ $Y2=3.235
cc_199 N_VDD_c_194_p N_D_M1021_g 0.00606474f $X=2.38 $Y=4.287 $X2=0.93 $Y2=3.235
cc_200 N_VDD_c_186_p N_D_M1021_g 0.00468827f $X=6.46 $Y=4.25 $X2=0.93 $Y2=3.235
cc_201 N_VDD_M1022_b N_CK_M1014_g 0.0201249f $X=-0.045 $Y=2.425 $X2=1.29
+ $Y2=3.235
cc_202 N_VDD_c_194_p N_CK_M1014_g 0.00606474f $X=2.38 $Y=4.287 $X2=1.29
+ $Y2=3.235
cc_203 N_VDD_c_186_p N_CK_M1014_g 0.00468827f $X=6.46 $Y=4.25 $X2=1.29 $Y2=3.235
cc_204 N_VDD_M1022_b N_CK_M1019_g 0.0201163f $X=-0.045 $Y=2.425 $X2=3.64
+ $Y2=3.235
cc_205 N_VDD_c_205_p N_CK_M1019_g 0.00606474f $X=4.13 $Y=4.287 $X2=3.64
+ $Y2=3.235
cc_206 N_VDD_c_186_p N_CK_M1019_g 0.00468827f $X=6.46 $Y=4.25 $X2=3.64 $Y2=3.235
cc_207 N_VDD_M1022_b N_CK_c_416_n 0.007968f $X=-0.045 $Y=2.425 $X2=4.43 $Y2=2.45
cc_208 N_VDD_M1022_b N_CK_M1017_g 0.0218804f $X=-0.045 $Y=2.425 $X2=4.43
+ $Y2=3.235
cc_209 N_VDD_c_209_p N_CK_M1017_g 0.0047242f $X=4.215 $Y=3.21 $X2=4.43 $Y2=3.235
cc_210 N_VDD_c_210_p N_CK_M1017_g 0.00606474f $X=5.08 $Y=4.287 $X2=4.43
+ $Y2=3.235
cc_211 N_VDD_c_211_p N_CK_M1017_g 0.00455736f $X=5.165 $Y=3.295 $X2=4.43
+ $Y2=3.235
cc_212 N_VDD_c_186_p N_CK_M1017_g 0.00468827f $X=6.46 $Y=4.25 $X2=4.43 $Y2=3.235
cc_213 N_VDD_M1022_b N_CK_c_418_n 0.0065467f $X=-0.045 $Y=2.425 $X2=1.38
+ $Y2=2.285
cc_214 N_VDD_M1022_b N_CK_c_427_n 0.00654388f $X=-0.045 $Y=2.425 $X2=3.55
+ $Y2=2.285
cc_215 N_VDD_M1022_b N_CK_c_439_n 0.0010436f $X=-0.045 $Y=2.425 $X2=4.575
+ $Y2=2.11
cc_216 N_VDD_M1022_b N_CK_c_440_n 9.30704e-19 $X=-0.045 $Y=2.425 $X2=1.35
+ $Y2=2.11
cc_217 N_VDD_M1022_b N_CK_c_441_n 0.00253381f $X=-0.045 $Y=2.425 $X2=3.58
+ $Y2=2.11
cc_218 N_VDD_M1022_b N_A_32_115#_M1004_g 0.0192219f $X=-0.045 $Y=2.425 $X2=2.25
+ $Y2=3.235
cc_219 N_VDD_c_194_p N_A_32_115#_M1004_g 0.00606474f $X=2.38 $Y=4.287 $X2=2.25
+ $Y2=3.235
cc_220 N_VDD_c_220_p N_A_32_115#_M1004_g 0.00337744f $X=2.465 $Y=3.295 $X2=2.25
+ $Y2=3.235
cc_221 N_VDD_c_186_p N_A_32_115#_M1004_g 0.00468827f $X=6.46 $Y=4.25 $X2=2.25
+ $Y2=3.235
cc_222 N_VDD_c_220_p N_A_32_115#_c_651_n 8.24975e-19 $X=2.465 $Y=3.295 $X2=2.605
+ $Y2=2.285
cc_223 N_VDD_M1022_b N_A_32_115#_M1006_g 0.0181098f $X=-0.045 $Y=2.425 $X2=2.68
+ $Y2=3.235
cc_224 N_VDD_c_220_p N_A_32_115#_M1006_g 0.00337744f $X=2.465 $Y=3.295 $X2=2.68
+ $Y2=3.235
cc_225 N_VDD_c_205_p N_A_32_115#_M1006_g 0.00606474f $X=4.13 $Y=4.287 $X2=2.68
+ $Y2=3.235
cc_226 N_VDD_c_186_p N_A_32_115#_M1006_g 0.00468827f $X=6.46 $Y=4.25 $X2=2.68
+ $Y2=3.235
cc_227 N_VDD_M1022_b N_A_32_115#_c_657_n 0.0120505f $X=-0.045 $Y=2.425 $X2=0.17
+ $Y2=2.695
cc_228 N_VDD_M1022_b N_A_32_115#_c_680_n 0.00156053f $X=-0.045 $Y=2.425
+ $X2=0.285 $Y2=2.955
cc_229 N_VDD_c_184_p N_A_32_115#_c_680_n 0.00736239f $X=0.63 $Y=4.287 $X2=0.285
+ $Y2=2.955
cc_230 N_VDD_c_186_p N_A_32_115#_c_680_n 0.00476261f $X=6.46 $Y=4.25 $X2=0.285
+ $Y2=2.955
cc_231 N_VDD_M1022_b N_A_32_115#_c_661_n 0.00424346f $X=-0.045 $Y=2.425 $X2=2.42
+ $Y2=2.285
cc_232 N_VDD_c_220_p N_A_32_115#_c_661_n 0.004428f $X=2.465 $Y=3.295 $X2=2.42
+ $Y2=2.285
cc_233 N_VDD_M1022_b N_A_32_115#_c_685_n 0.0093744f $X=-0.045 $Y=2.425 $X2=0.285
+ $Y2=2.78
cc_234 N_VDD_M1022_b N_A_243_89#_M1011_g 0.0214581f $X=-0.045 $Y=2.425 $X2=1.89
+ $Y2=3.235
cc_235 N_VDD_c_194_p N_A_243_89#_M1011_g 0.00606474f $X=2.38 $Y=4.287 $X2=1.89
+ $Y2=3.235
cc_236 N_VDD_c_186_p N_A_243_89#_M1011_g 0.00468827f $X=6.46 $Y=4.25 $X2=1.89
+ $Y2=3.235
cc_237 N_VDD_M1022_b N_A_243_89#_M1003_g 0.0214271f $X=-0.045 $Y=2.425 $X2=3.04
+ $Y2=3.235
cc_238 N_VDD_c_205_p N_A_243_89#_M1003_g 0.00606474f $X=4.13 $Y=4.287 $X2=3.04
+ $Y2=3.235
cc_239 N_VDD_c_186_p N_A_243_89#_M1003_g 0.00468827f $X=6.46 $Y=4.25 $X2=3.04
+ $Y2=3.235
cc_240 N_VDD_M1022_b N_A_243_89#_c_792_n 0.00156053f $X=-0.045 $Y=2.425
+ $X2=4.645 $Y2=2.955
cc_241 N_VDD_c_210_p N_A_243_89#_c_792_n 0.00749582f $X=5.08 $Y=4.287 $X2=4.645
+ $Y2=2.955
cc_242 N_VDD_c_211_p N_A_243_89#_c_792_n 0.0341747f $X=5.165 $Y=3.295 $X2=4.645
+ $Y2=2.955
cc_243 N_VDD_c_186_p N_A_243_89#_c_792_n 0.00476261f $X=6.46 $Y=4.25 $X2=4.645
+ $Y2=2.955
cc_244 N_VDD_M1022_b N_A_243_89#_c_781_n 0.00543969f $X=-0.045 $Y=2.425
+ $X2=4.915 $Y2=2.62
cc_245 N_VDD_M1022_b N_A_243_89#_c_797_n 0.0119291f $X=-0.045 $Y=2.425 $X2=4.915
+ $Y2=2.705
cc_246 N_VDD_M1022_b N_A_785_89#_M1016_g 0.0178558f $X=-0.045 $Y=2.425 $X2=4
+ $Y2=3.235
cc_247 N_VDD_c_205_p N_A_785_89#_M1016_g 0.00606474f $X=4.13 $Y=4.287 $X2=4
+ $Y2=3.235
cc_248 N_VDD_c_209_p N_A_785_89#_M1016_g 0.0047242f $X=4.215 $Y=3.21 $X2=4
+ $Y2=3.235
cc_249 N_VDD_c_186_p N_A_785_89#_M1016_g 0.00468827f $X=6.46 $Y=4.25 $X2=4
+ $Y2=3.235
cc_250 N_VDD_M1022_b N_A_785_89#_c_965_n 0.0277135f $X=-0.045 $Y=2.425 $X2=6.305
+ $Y2=2.49
cc_251 N_VDD_c_251_p N_A_785_89#_c_965_n 0.00606474f $X=6.46 $Y=4.287 $X2=6.305
+ $Y2=2.49
cc_252 N_VDD_c_252_p N_A_785_89#_c_965_n 0.00354579f $X=6.545 $Y=3.615 $X2=6.305
+ $Y2=2.49
cc_253 N_VDD_c_186_p N_A_785_89#_c_965_n 0.00468827f $X=6.46 $Y=4.25 $X2=6.305
+ $Y2=2.49
cc_254 N_VDD_M1022_b N_A_785_89#_c_967_n 0.00241422f $X=-0.045 $Y=2.425 $X2=4.06
+ $Y2=2.48
cc_255 N_VDD_c_209_p N_A_785_89#_c_967_n 0.00121222f $X=4.215 $Y=3.21 $X2=4.06
+ $Y2=2.48
cc_256 N_VDD_M1022_b N_A_785_89#_c_971_n 0.00576734f $X=-0.045 $Y=2.425
+ $X2=5.595 $Y2=2.955
cc_257 N_VDD_c_251_p N_A_785_89#_c_971_n 0.0074445f $X=6.46 $Y=4.287 $X2=5.595
+ $Y2=2.955
cc_258 N_VDD_c_186_p N_A_785_89#_c_971_n 0.00476261f $X=6.46 $Y=4.25 $X2=5.595
+ $Y2=2.955
cc_259 N_VDD_M1022_b N_A_785_89#_c_974_n 0.011211f $X=-0.045 $Y=2.425 $X2=4.935
+ $Y2=2.48
cc_260 N_VDD_c_209_p N_A_785_89#_c_974_n 0.00492996f $X=4.215 $Y=3.21 $X2=4.935
+ $Y2=2.48
cc_261 N_VDD_M1022_b N_A_785_89#_c_975_n 0.00594814f $X=-0.045 $Y=2.425
+ $X2=4.205 $Y2=2.48
cc_262 N_VDD_c_209_p N_A_785_89#_c_975_n 0.00366258f $X=4.215 $Y=3.21 $X2=4.205
+ $Y2=2.48
cc_263 N_VDD_M1022_b N_A_623_115#_M1023_g 0.0260072f $X=-0.045 $Y=2.425 $X2=5.38
+ $Y2=3.235
cc_264 N_VDD_c_211_p N_A_623_115#_M1023_g 0.00636672f $X=5.165 $Y=3.295 $X2=5.38
+ $Y2=3.235
cc_265 N_VDD_c_251_p N_A_623_115#_M1023_g 0.00606474f $X=6.46 $Y=4.287 $X2=5.38
+ $Y2=3.235
cc_266 N_VDD_c_186_p N_A_623_115#_M1023_g 0.00468827f $X=6.46 $Y=4.25 $X2=5.38
+ $Y2=3.235
cc_267 N_VDD_M1022_b N_A_623_115#_c_1124_n 0.00167876f $X=-0.045 $Y=2.425
+ $X2=2.76 $Y2=1.37
cc_268 N_VDD_M1022_b N_A_623_115#_c_1143_n 0.00313975f $X=-0.045 $Y=2.425
+ $X2=3.34 $Y2=3.295
cc_269 N_VDD_c_205_p N_A_623_115#_c_1143_n 0.0151257f $X=4.13 $Y=4.287 $X2=3.34
+ $Y2=3.295
cc_270 N_VDD_c_186_p N_A_623_115#_c_1143_n 0.00958198f $X=6.46 $Y=4.25 $X2=3.34
+ $Y2=3.295
cc_271 N_VDD_M1022_b N_ON_M1018_g 0.0267313f $X=-0.045 $Y=2.425 $X2=6.76
+ $Y2=3.235
cc_272 N_VDD_c_252_p N_ON_M1018_g 0.00354579f $X=6.545 $Y=3.615 $X2=6.76
+ $Y2=3.235
cc_273 N_VDD_c_273_p N_ON_M1018_g 0.00606474f $X=6.46 $Y=4.25 $X2=6.76 $Y2=3.235
cc_274 N_VDD_c_186_p N_ON_M1018_g 0.00468827f $X=6.46 $Y=4.25 $X2=6.76 $Y2=3.235
cc_275 N_VDD_M1022_b N_ON_c_1249_n 0.00535667f $X=-0.045 $Y=2.425 $X2=6.115
+ $Y2=3.615
cc_276 N_VDD_c_251_p N_ON_c_1249_n 0.00757793f $X=6.46 $Y=4.287 $X2=6.115
+ $Y2=3.615
cc_277 N_VDD_c_186_p N_ON_c_1249_n 0.00476261f $X=6.46 $Y=4.25 $X2=6.115
+ $Y2=3.615
cc_278 N_VDD_M1022_b N_Q_c_1326_n 0.00156053f $X=-0.045 $Y=2.425 $X2=6.975
+ $Y2=3.615
cc_279 N_VDD_c_273_p N_Q_c_1326_n 0.00757793f $X=6.46 $Y=4.25 $X2=6.975
+ $Y2=3.615
cc_280 N_VDD_c_186_p N_Q_c_1326_n 0.00476261f $X=6.46 $Y=4.25 $X2=6.975
+ $Y2=3.615
cc_281 N_VDD_M1022_b N_Q_c_1323_n 0.0111162f $X=-0.045 $Y=2.425 $X2=7.09
+ $Y2=2.48
cc_282 N_VDD_M1022_b N_Q_c_1330_n 0.00144175f $X=-0.045 $Y=2.425 $X2=6.972
+ $Y2=2.88
cc_283 N_VDD_M1022_b Q 0.00549803f $X=-0.045 $Y=2.425 $X2=6.97 $Y2=2.48
cc_284 N_A_75_248#_c_284_n N_D_M1007_g 0.0247367f $X=0.475 $Y=1.24 $X2=0.93
+ $Y2=0.85
cc_285 N_A_75_248#_c_290_n N_D_M1007_g 0.022942f $X=0.51 $Y=2.12 $X2=0.93
+ $Y2=0.85
cc_286 N_A_75_248#_c_291_n N_D_M1007_g 0.0146593f $X=1.405 $Y=1.285 $X2=0.93
+ $Y2=0.85
cc_287 N_A_75_248#_c_297_n N_D_M1007_g 0.00559668f $X=0.567 $Y=2.12 $X2=0.93
+ $Y2=0.85
cc_288 N_A_75_248#_M1022_g N_D_M1021_g 0.0342437f $X=0.5 $Y=3.235 $X2=0.93
+ $Y2=3.235
cc_289 N_A_75_248#_c_289_n N_D_M1021_g 0.0194268f $X=0.51 $Y=2.285 $X2=0.93
+ $Y2=3.235
cc_290 N_A_75_248#_c_306_n N_D_M1021_g 0.00559668f $X=0.625 $Y=2.62 $X2=0.93
+ $Y2=3.235
cc_291 N_A_75_248#_c_307_n N_D_M1021_g 0.019095f $X=1.42 $Y=2.705 $X2=0.93
+ $Y2=3.235
cc_292 N_A_75_248#_c_291_n N_D_c_378_n 0.00207628f $X=1.405 $Y=1.285 $X2=0.99
+ $Y2=1.74
cc_293 N_A_75_248#_c_296_n N_D_c_378_n 0.00559668f $X=0.51 $Y=2.285 $X2=0.99
+ $Y2=1.74
cc_294 N_A_75_248#_c_291_n N_D_c_379_n 0.0086486f $X=1.405 $Y=1.285 $X2=0.99
+ $Y2=1.74
cc_295 N_A_75_248#_c_297_n N_D_c_379_n 0.0187793f $X=0.567 $Y=2.12 $X2=0.99
+ $Y2=1.74
cc_296 N_A_75_248#_c_291_n D 0.00200799f $X=1.405 $Y=1.285 $X2=0.99 $Y2=1.74
cc_297 N_A_75_248#_c_297_n D 0.007232f $X=0.567 $Y=2.12 $X2=0.99 $Y2=1.74
cc_298 N_A_75_248#_c_307_n N_CK_M1014_g 0.0156056f $X=1.42 $Y=2.705 $X2=1.29
+ $Y2=3.235
cc_299 N_A_75_248#_c_307_n N_CK_c_418_n 0.00248712f $X=1.42 $Y=2.705 $X2=1.38
+ $Y2=2.285
cc_300 N_A_75_248#_c_291_n N_CK_c_419_n 7.46335e-19 $X=1.405 $Y=1.285 $X2=1.83
+ $Y2=1.4
cc_301 N_A_75_248#_c_298_n N_CK_c_419_n 0.00190388f $X=1.49 $Y=0.755 $X2=1.83
+ $Y2=1.4
cc_302 N_A_75_248#_c_291_n N_CK_c_420_n 9.05754e-19 $X=1.405 $Y=1.285 $X2=1.83
+ $Y2=1.235
cc_303 N_A_75_248#_c_295_n N_CK_c_420_n 0.00540119f $X=1.49 $Y=1.2 $X2=1.83
+ $Y2=1.235
cc_304 N_A_75_248#_c_291_n N_CK_c_434_n 0.00160862f $X=1.405 $Y=1.285 $X2=1.745
+ $Y2=2.11
cc_305 N_A_75_248#_c_307_n N_CK_c_434_n 0.0081057f $X=1.42 $Y=2.705 $X2=1.745
+ $Y2=2.11
cc_306 N_A_75_248#_c_291_n N_CK_c_435_n 0.00989572f $X=1.405 $Y=1.285 $X2=1.83
+ $Y2=1.4
cc_307 N_A_75_248#_c_298_n N_CK_c_435_n 6.02618e-19 $X=1.49 $Y=0.755 $X2=1.83
+ $Y2=1.4
cc_308 N_A_75_248#_c_291_n N_CK_c_440_n 0.00263105f $X=1.405 $Y=1.285 $X2=1.35
+ $Y2=2.11
cc_309 N_A_75_248#_c_307_n N_CK_c_440_n 0.0111655f $X=1.42 $Y=2.705 $X2=1.35
+ $Y2=2.11
cc_310 N_A_75_248#_c_296_n N_CK_c_440_n 0.00703951f $X=0.51 $Y=2.285 $X2=1.35
+ $Y2=2.11
cc_311 N_A_75_248#_c_297_n N_CK_c_440_n 0.00315097f $X=0.567 $Y=2.12 $X2=1.35
+ $Y2=2.11
cc_312 N_A_75_248#_c_307_n N_CK_c_442_n 0.00596172f $X=1.42 $Y=2.705 $X2=3.435
+ $Y2=2.11
cc_313 N_A_75_248#_c_307_n N_CK_c_443_n 0.00395573f $X=1.42 $Y=2.705 $X2=1.495
+ $Y2=2.11
cc_314 N_A_75_248#_c_297_n N_CK_c_443_n 0.00642669f $X=0.567 $Y=2.12 $X2=1.495
+ $Y2=2.11
cc_315 N_A_75_248#_M1022_g N_A_32_115#_c_657_n 0.00498045f $X=0.5 $Y=3.235
+ $X2=0.17 $Y2=2.695
cc_316 N_A_75_248#_c_290_n N_A_32_115#_c_657_n 0.0218335f $X=0.51 $Y=2.12
+ $X2=0.17 $Y2=2.695
cc_317 N_A_75_248#_c_306_n N_A_32_115#_c_657_n 0.00821014f $X=0.625 $Y=2.62
+ $X2=0.17 $Y2=2.695
cc_318 N_A_75_248#_c_309_n N_A_32_115#_c_657_n 0.00395316f $X=0.71 $Y=2.705
+ $X2=0.17 $Y2=2.695
cc_319 N_A_75_248#_c_296_n N_A_32_115#_c_657_n 0.0245251f $X=0.51 $Y=2.285
+ $X2=0.17 $Y2=2.695
cc_320 N_A_75_248#_c_297_n N_A_32_115#_c_657_n 0.0334082f $X=0.567 $Y=2.12
+ $X2=0.17 $Y2=2.695
cc_321 N_A_75_248#_c_284_n N_A_32_115#_c_658_n 0.00546712f $X=0.475 $Y=1.24
+ $X2=0.285 $Y2=0.755
cc_322 N_A_75_248#_c_284_n N_A_32_115#_c_662_n 0.00165831f $X=0.475 $Y=1.24
+ $X2=0.285 $Y2=1.37
cc_323 N_A_75_248#_c_288_n N_A_32_115#_c_662_n 0.00460749f $X=0.475 $Y=1.39
+ $X2=0.285 $Y2=1.37
cc_324 N_A_75_248#_c_293_n N_A_32_115#_c_662_n 0.0125535f $X=0.71 $Y=1.285
+ $X2=0.285 $Y2=1.37
cc_325 N_A_75_248#_c_297_n N_A_32_115#_c_662_n 0.00592135f $X=0.567 $Y=2.12
+ $X2=0.285 $Y2=1.37
cc_326 N_A_75_248#_c_288_n N_A_32_115#_c_665_n 0.0047054f $X=0.475 $Y=1.39
+ $X2=2.185 $Y2=1.37
cc_327 N_A_75_248#_c_290_n N_A_32_115#_c_665_n 0.0043937f $X=0.51 $Y=2.12
+ $X2=2.185 $Y2=1.37
cc_328 N_A_75_248#_c_291_n N_A_32_115#_c_665_n 0.0597786f $X=1.405 $Y=1.285
+ $X2=2.185 $Y2=1.37
cc_329 N_A_75_248#_c_293_n N_A_32_115#_c_665_n 0.00750079f $X=0.71 $Y=1.285
+ $X2=2.185 $Y2=1.37
cc_330 N_A_75_248#_c_297_n N_A_32_115#_c_665_n 0.0143756f $X=0.567 $Y=2.12
+ $X2=2.185 $Y2=1.37
cc_331 N_A_75_248#_c_298_n N_A_32_115#_c_665_n 0.0070752f $X=1.49 $Y=0.755
+ $X2=2.185 $Y2=1.37
cc_332 N_A_75_248#_c_288_n N_A_32_115#_c_667_n 0.00387046f $X=0.475 $Y=1.39
+ $X2=0.43 $Y2=1.37
cc_333 N_A_75_248#_c_290_n N_A_32_115#_c_667_n 0.00369116f $X=0.51 $Y=2.12
+ $X2=0.43 $Y2=1.37
cc_334 N_A_75_248#_c_293_n N_A_32_115#_c_667_n 8.15236e-19 $X=0.71 $Y=1.285
+ $X2=0.43 $Y2=1.37
cc_335 N_A_75_248#_c_297_n N_A_32_115#_c_667_n 8.59347e-19 $X=0.567 $Y=2.12
+ $X2=0.43 $Y2=1.37
cc_336 N_A_75_248#_c_291_n N_A_243_89#_c_759_n 0.0066768f $X=1.405 $Y=1.285
+ $X2=1.29 $Y2=1.205
cc_337 N_A_75_248#_c_295_n N_A_243_89#_c_759_n 0.00317892f $X=1.49 $Y=1.2
+ $X2=1.29 $Y2=1.205
cc_338 N_A_75_248#_c_291_n N_A_243_89#_c_762_n 0.00333286f $X=1.405 $Y=1.285
+ $X2=1.41 $Y2=1.775
cc_339 N_A_75_248#_c_307_n N_A_243_89#_c_763_n 6.56088e-19 $X=1.42 $Y=2.705
+ $X2=1.815 $Y2=1.85
cc_340 N_A_75_248#_c_291_n N_A_243_89#_c_772_n 0.00993421f $X=1.405 $Y=1.285
+ $X2=1.41 $Y2=1.28
cc_341 N_A_75_248#_c_307_n A_201_521# 0.00732587f $X=1.42 $Y=2.705 $X2=1.005
+ $Y2=2.605
cc_342 N_D_M1021_g N_CK_c_418_n 0.111906f $X=0.93 $Y=3.235 $X2=1.38 $Y2=2.285
cc_343 N_D_c_379_n N_CK_c_435_n 0.00479659f $X=0.99 $Y=1.74 $X2=1.83 $Y2=1.4
cc_344 D N_CK_c_435_n 0.00555005f $X=0.99 $Y=1.74 $X2=1.83 $Y2=1.4
cc_345 N_D_M1021_g N_CK_c_440_n 0.00358312f $X=0.93 $Y=3.235 $X2=1.35 $Y2=2.11
cc_346 N_D_M1021_g N_CK_c_443_n 0.00542304f $X=0.93 $Y=3.235 $X2=1.495 $Y2=2.11
cc_347 D N_CK_c_443_n 0.00375733f $X=0.99 $Y=1.74 $X2=1.495 $Y2=2.11
cc_348 N_D_M1007_g N_A_32_115#_c_665_n 0.00223521f $X=0.93 $Y=0.85 $X2=2.185
+ $Y2=1.37
cc_349 N_D_c_378_n N_A_32_115#_c_665_n 7.9412e-19 $X=0.99 $Y=1.74 $X2=2.185
+ $Y2=1.37
cc_350 N_D_c_379_n N_A_32_115#_c_665_n 0.00111625f $X=0.99 $Y=1.74 $X2=2.185
+ $Y2=1.37
cc_351 D N_A_32_115#_c_665_n 0.0353362f $X=0.99 $Y=1.74 $X2=2.185 $Y2=1.37
cc_352 N_D_M1007_g N_A_243_89#_c_759_n 0.0553906f $X=0.93 $Y=0.85 $X2=1.29
+ $Y2=1.205
cc_353 N_D_M1007_g N_A_243_89#_c_762_n 0.00886317f $X=0.93 $Y=0.85 $X2=1.41
+ $Y2=1.775
cc_354 N_D_c_378_n N_A_243_89#_c_762_n 0.0214858f $X=0.99 $Y=1.74 $X2=1.41
+ $Y2=1.775
cc_355 N_D_c_379_n N_A_243_89#_c_762_n 0.00166174f $X=0.99 $Y=1.74 $X2=1.41
+ $Y2=1.775
cc_356 D N_A_243_89#_c_762_n 0.00338565f $X=0.99 $Y=1.74 $X2=1.41 $Y2=1.775
cc_357 N_D_M1021_g N_A_243_89#_c_764_n 8.72885e-19 $X=0.93 $Y=3.235 $X2=1.485
+ $Y2=1.85
cc_358 D N_A_243_89#_c_764_n 4.62757e-19 $X=0.99 $Y=1.74 $X2=1.485 $Y2=1.85
cc_359 N_CK_c_420_n N_A_32_115#_M1013_g 0.0342837f $X=1.83 $Y=1.235 $X2=2.25
+ $Y2=0.85
cc_360 N_CK_c_435_n N_A_32_115#_M1013_g 0.00109085f $X=1.83 $Y=1.4 $X2=2.25
+ $Y2=0.85
cc_361 N_CK_c_423_n N_A_32_115#_c_648_n 0.033846f $X=3.1 $Y=1.4 $X2=2.605
+ $Y2=1.4
cc_362 N_CK_c_436_n N_A_32_115#_c_648_n 3.18936e-19 $X=3.1 $Y=1.4 $X2=2.605
+ $Y2=1.4
cc_363 N_CK_c_419_n N_A_32_115#_c_650_n 0.0342837f $X=1.83 $Y=1.4 $X2=2.325
+ $Y2=1.4
cc_364 N_CK_c_442_n N_A_32_115#_c_651_n 0.00765556f $X=3.435 $Y=2.11 $X2=2.605
+ $Y2=2.285
cc_365 N_CK_c_442_n N_A_32_115#_c_652_n 0.00673865f $X=3.435 $Y=2.11 $X2=2.325
+ $Y2=2.285
cc_366 N_CK_c_424_n N_A_32_115#_M1015_g 0.033846f $X=3.1 $Y=1.235 $X2=2.68
+ $Y2=0.85
cc_367 N_CK_c_419_n N_A_32_115#_c_661_n 8.1208e-19 $X=1.83 $Y=1.4 $X2=2.42
+ $Y2=2.285
cc_368 N_CK_c_434_n N_A_32_115#_c_661_n 0.00402252f $X=1.745 $Y=2.11 $X2=2.42
+ $Y2=2.285
cc_369 N_CK_c_435_n N_A_32_115#_c_661_n 0.0202707f $X=1.83 $Y=1.4 $X2=2.42
+ $Y2=2.285
cc_370 N_CK_c_442_n N_A_32_115#_c_661_n 0.0206843f $X=3.435 $Y=2.11 $X2=2.42
+ $Y2=2.285
cc_371 N_CK_c_419_n N_A_32_115#_c_663_n 6.279e-19 $X=1.83 $Y=1.4 $X2=2.42
+ $Y2=1.4
cc_372 N_CK_c_435_n N_A_32_115#_c_663_n 0.00643639f $X=1.83 $Y=1.4 $X2=2.42
+ $Y2=1.4
cc_373 N_CK_c_436_n N_A_32_115#_c_663_n 9.81026e-19 $X=3.1 $Y=1.4 $X2=2.42
+ $Y2=1.4
cc_374 N_CK_c_442_n N_A_32_115#_c_663_n 0.00102309f $X=3.435 $Y=2.11 $X2=2.42
+ $Y2=1.4
cc_375 N_CK_c_419_n N_A_32_115#_c_665_n 0.00577781f $X=1.83 $Y=1.4 $X2=2.185
+ $Y2=1.37
cc_376 N_CK_c_434_n N_A_32_115#_c_665_n 0.0043165f $X=1.745 $Y=2.11 $X2=2.185
+ $Y2=1.37
cc_377 N_CK_c_435_n N_A_32_115#_c_665_n 0.0204213f $X=1.83 $Y=1.4 $X2=2.185
+ $Y2=1.37
cc_378 N_CK_c_440_n N_A_32_115#_c_665_n 8.37938e-19 $X=1.35 $Y=2.11 $X2=2.185
+ $Y2=1.37
cc_379 N_CK_c_443_n N_A_32_115#_c_665_n 0.0126162f $X=1.495 $Y=2.11 $X2=2.185
+ $Y2=1.37
cc_380 N_CK_c_419_n N_A_32_115#_c_668_n 3.26623e-19 $X=1.83 $Y=1.4 $X2=2.33
+ $Y2=1.37
cc_381 N_CK_c_435_n N_A_32_115#_c_668_n 0.00141649f $X=1.83 $Y=1.4 $X2=2.33
+ $Y2=1.37
cc_382 N_CK_c_442_n N_A_32_115#_c_668_n 0.0129652f $X=3.435 $Y=2.11 $X2=2.33
+ $Y2=1.37
cc_383 N_CK_c_420_n N_A_243_89#_c_759_n 0.0152188f $X=1.83 $Y=1.235 $X2=1.29
+ $Y2=1.205
cc_384 N_CK_c_435_n N_A_243_89#_c_762_n 0.00602582f $X=1.83 $Y=1.4 $X2=1.41
+ $Y2=1.775
cc_385 N_CK_c_419_n N_A_243_89#_c_763_n 0.0183472f $X=1.83 $Y=1.4 $X2=1.815
+ $Y2=1.85
cc_386 N_CK_c_435_n N_A_243_89#_c_763_n 0.00665821f $X=1.83 $Y=1.4 $X2=1.815
+ $Y2=1.85
cc_387 N_CK_c_442_n N_A_243_89#_c_763_n 0.00549601f $X=3.435 $Y=2.11 $X2=1.815
+ $Y2=1.85
cc_388 N_CK_c_418_n N_A_243_89#_c_764_n 0.012591f $X=1.38 $Y=2.285 $X2=1.485
+ $Y2=1.85
cc_389 N_CK_c_434_n N_A_243_89#_c_764_n 0.00756374f $X=1.745 $Y=2.11 $X2=1.485
+ $Y2=1.85
cc_390 N_CK_c_440_n N_A_243_89#_c_764_n 0.00154604f $X=1.35 $Y=2.11 $X2=1.485
+ $Y2=1.85
cc_391 N_CK_c_443_n N_A_243_89#_c_764_n 0.00130179f $X=1.495 $Y=2.11 $X2=1.485
+ $Y2=1.85
cc_392 N_CK_M1014_g N_A_243_89#_M1011_g 0.0315947f $X=1.29 $Y=3.235 $X2=1.89
+ $Y2=3.235
cc_393 N_CK_c_418_n N_A_243_89#_M1011_g 0.014942f $X=1.38 $Y=2.285 $X2=1.89
+ $Y2=3.235
cc_394 N_CK_c_434_n N_A_243_89#_M1011_g 0.00849934f $X=1.745 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_395 N_CK_c_435_n N_A_243_89#_M1011_g 0.00368559f $X=1.83 $Y=1.4 $X2=1.89
+ $Y2=3.235
cc_396 N_CK_c_440_n N_A_243_89#_M1011_g 0.00148098f $X=1.35 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_397 N_CK_c_442_n N_A_243_89#_M1011_g 0.00937774f $X=3.435 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_398 N_CK_c_442_n N_A_243_89#_c_766_n 0.00615595f $X=3.435 $Y=2.11 $X2=2.965
+ $Y2=1.85
cc_399 N_CK_M1019_g N_A_243_89#_M1003_g 0.0316011f $X=3.64 $Y=3.235 $X2=3.04
+ $Y2=3.235
cc_400 N_CK_c_427_n N_A_243_89#_M1003_g 0.0138379f $X=3.55 $Y=2.285 $X2=3.04
+ $Y2=3.235
cc_401 N_CK_c_436_n N_A_243_89#_M1003_g 0.00305863f $X=3.1 $Y=1.4 $X2=3.04
+ $Y2=3.235
cc_402 N_CK_c_438_n N_A_243_89#_M1003_g 0.00692515f $X=3.185 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_403 N_CK_c_441_n N_A_243_89#_M1003_g 8.92314e-19 $X=3.58 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_404 N_CK_c_442_n N_A_243_89#_M1003_g 0.00496221f $X=3.435 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_405 N_CK_c_427_n N_A_243_89#_c_768_n 0.0199686f $X=3.55 $Y=2.285 $X2=3.445
+ $Y2=1.85
cc_406 N_CK_c_436_n N_A_243_89#_c_768_n 0.00708423f $X=3.1 $Y=1.4 $X2=3.445
+ $Y2=1.85
cc_407 N_CK_c_437_n N_A_243_89#_c_768_n 0.00731605f $X=3.465 $Y=2.11 $X2=3.445
+ $Y2=1.85
cc_408 N_CK_c_442_n N_A_243_89#_c_768_n 0.00530993f $X=3.435 $Y=2.11 $X2=3.445
+ $Y2=1.85
cc_409 N_CK_c_445_n N_A_243_89#_c_768_n 0.00125555f $X=3.725 $Y=2.11 $X2=3.445
+ $Y2=1.85
cc_410 N_CK_c_423_n N_A_243_89#_M1005_g 0.0132483f $X=3.1 $Y=1.4 $X2=3.64
+ $Y2=0.85
cc_411 N_CK_c_424_n N_A_243_89#_M1005_g 0.015655f $X=3.1 $Y=1.235 $X2=3.64
+ $Y2=0.85
cc_412 N_CK_c_436_n N_A_243_89#_M1005_g 9.94573e-19 $X=3.1 $Y=1.4 $X2=3.64
+ $Y2=0.85
cc_413 N_CK_c_419_n N_A_243_89#_c_772_n 0.0216996f $X=1.83 $Y=1.4 $X2=1.41
+ $Y2=1.28
cc_414 N_CK_c_420_n N_A_243_89#_c_772_n 9.76811e-19 $X=1.83 $Y=1.235 $X2=1.41
+ $Y2=1.28
cc_415 N_CK_c_440_n N_A_243_89#_c_772_n 2.43077e-19 $X=1.35 $Y=2.11 $X2=1.41
+ $Y2=1.28
cc_416 N_CK_c_435_n N_A_243_89#_c_773_n 0.00568091f $X=1.83 $Y=1.4 $X2=1.89
+ $Y2=1.85
cc_417 N_CK_c_423_n N_A_243_89#_c_774_n 0.0183472f $X=3.1 $Y=1.4 $X2=3.04
+ $Y2=1.85
cc_418 N_CK_c_436_n N_A_243_89#_c_774_n 0.00436024f $X=3.1 $Y=1.4 $X2=3.04
+ $Y2=1.85
cc_419 N_CK_c_436_n N_A_243_89#_c_775_n 0.00327058f $X=3.1 $Y=1.4 $X2=3.58
+ $Y2=1.74
cc_420 N_CK_c_441_n N_A_243_89#_c_775_n 0.00136839f $X=3.58 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_421 N_CK_c_427_n N_A_243_89#_c_776_n 7.64371e-19 $X=3.55 $Y=2.285 $X2=3.58
+ $Y2=1.74
cc_422 N_CK_c_436_n N_A_243_89#_c_776_n 0.00799667f $X=3.1 $Y=1.4 $X2=3.58
+ $Y2=1.74
cc_423 N_CK_c_437_n N_A_243_89#_c_776_n 0.00282541f $X=3.465 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_424 N_CK_c_441_n N_A_243_89#_c_776_n 0.0116376f $X=3.58 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_425 N_CK_c_444_n N_A_243_89#_c_776_n 5.17303e-19 $X=4.43 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_426 N_CK_c_445_n N_A_243_89#_c_776_n 0.00180359f $X=3.725 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_427 N_CK_c_428_n N_A_243_89#_c_777_n 0.00641826f $X=4.457 $Y=1.205 $X2=4.645
+ $Y2=0.755
cc_428 N_CK_c_433_n N_A_243_89#_c_777_n 0.0125898f $X=4.457 $Y=1.355 $X2=4.645
+ $Y2=0.755
cc_429 N_CK_c_416_n N_A_243_89#_c_781_n 0.00318866f $X=4.43 $Y=2.45 $X2=4.915
+ $Y2=2.62
cc_430 N_CK_M1017_g N_A_243_89#_c_781_n 0.00395773f $X=4.43 $Y=3.235 $X2=4.915
+ $Y2=2.62
cc_431 N_CK_c_417_n N_A_243_89#_c_781_n 0.00561766f $X=4.485 $Y=2.12 $X2=4.915
+ $Y2=2.62
cc_432 N_CK_c_439_n N_A_243_89#_c_781_n 0.0277441f $X=4.575 $Y=2.11 $X2=4.915
+ $Y2=2.62
cc_433 CK N_A_243_89#_c_781_n 0.00256489f $X=4.575 $Y=2.11 $X2=4.915 $Y2=2.62
cc_434 N_CK_c_416_n N_A_243_89#_c_797_n 0.00233394f $X=4.43 $Y=2.45 $X2=4.915
+ $Y2=2.705
cc_435 N_CK_c_439_n N_A_243_89#_c_797_n 0.00601935f $X=4.575 $Y=2.11 $X2=4.915
+ $Y2=2.705
cc_436 N_CK_c_416_n N_A_243_89#_c_782_n 0.00178821f $X=4.43 $Y=2.45 $X2=4.645
+ $Y2=1.74
cc_437 N_CK_c_417_n N_A_243_89#_c_782_n 0.00516589f $X=4.485 $Y=2.12 $X2=4.645
+ $Y2=1.74
cc_438 N_CK_c_439_n N_A_243_89#_c_782_n 0.00622889f $X=4.575 $Y=2.11 $X2=4.645
+ $Y2=1.74
cc_439 CK N_A_243_89#_c_782_n 7.47532e-19 $X=4.575 $Y=2.11 $X2=4.645 $Y2=1.74
cc_440 N_CK_c_436_n N_A_243_89#_c_783_n 0.00363658f $X=3.1 $Y=1.4 $X2=3.725
+ $Y2=1.725
cc_441 N_CK_c_441_n N_A_243_89#_c_783_n 5.68393e-19 $X=3.58 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_442 N_CK_c_442_n N_A_243_89#_c_783_n 0.00163817f $X=3.435 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_443 N_CK_c_445_n N_A_243_89#_c_783_n 0.0296304f $X=3.725 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_444 N_CK_c_416_n N_A_243_89#_c_784_n 2.36275e-19 $X=4.43 $Y=2.45 $X2=4.645
+ $Y2=1.74
cc_445 N_CK_c_417_n N_A_243_89#_c_784_n 0.00251055f $X=4.485 $Y=2.12 $X2=4.645
+ $Y2=1.74
cc_446 N_CK_c_439_n N_A_243_89#_c_784_n 0.00129883f $X=4.575 $Y=2.11 $X2=4.645
+ $Y2=1.74
cc_447 CK N_A_243_89#_c_784_n 0.0226502f $X=4.575 $Y=2.11 $X2=4.645 $Y2=1.74
cc_448 N_CK_c_417_n N_A_243_89#_c_785_n 0.00278025f $X=4.485 $Y=2.12 $X2=4.5
+ $Y2=1.74
cc_449 N_CK_c_433_n N_A_243_89#_c_785_n 2.64649e-19 $X=4.457 $Y=1.355 $X2=4.5
+ $Y2=1.74
cc_450 N_CK_c_444_n N_A_243_89#_c_785_n 0.0538111f $X=4.43 $Y=2.11 $X2=4.5
+ $Y2=1.74
cc_451 CK N_A_243_89#_c_785_n 0.00582134f $X=4.575 $Y=2.11 $X2=4.5 $Y2=1.74
cc_452 N_CK_c_417_n N_A_785_89#_M1000_g 0.00866378f $X=4.485 $Y=2.12 $X2=4
+ $Y2=0.85
cc_453 N_CK_c_428_n N_A_785_89#_M1000_g 0.0236863f $X=4.457 $Y=1.205 $X2=4
+ $Y2=0.85
cc_454 N_CK_c_416_n N_A_785_89#_M1016_g 0.0389285f $X=4.43 $Y=2.45 $X2=4
+ $Y2=3.235
cc_455 N_CK_c_417_n N_A_785_89#_M1016_g 0.0139901f $X=4.485 $Y=2.12 $X2=4
+ $Y2=3.235
cc_456 N_CK_c_427_n N_A_785_89#_M1016_g 0.11066f $X=3.55 $Y=2.285 $X2=4
+ $Y2=3.235
cc_457 N_CK_c_439_n N_A_785_89#_M1016_g 5.87562e-19 $X=4.575 $Y=2.11 $X2=4
+ $Y2=3.235
cc_458 N_CK_c_441_n N_A_785_89#_M1016_g 0.0026293f $X=3.58 $Y=2.11 $X2=4
+ $Y2=3.235
cc_459 N_CK_c_444_n N_A_785_89#_M1016_g 0.00326152f $X=4.43 $Y=2.11 $X2=4
+ $Y2=3.235
cc_460 N_CK_c_445_n N_A_785_89#_M1016_g 0.00113587f $X=3.725 $Y=2.11 $X2=4
+ $Y2=3.235
cc_461 N_CK_c_417_n N_A_785_89#_c_962_n 0.0205509f $X=4.485 $Y=2.12 $X2=4.06
+ $Y2=1.74
cc_462 N_CK_c_444_n N_A_785_89#_c_962_n 7.38456e-19 $X=4.43 $Y=2.11 $X2=4.06
+ $Y2=1.74
cc_463 N_CK_c_417_n N_A_785_89#_c_966_n 8.16378e-19 $X=4.485 $Y=2.12 $X2=4.062
+ $Y2=1.812
cc_464 N_CK_c_416_n N_A_785_89#_c_967_n 0.00276728f $X=4.43 $Y=2.45 $X2=4.06
+ $Y2=2.48
cc_465 N_CK_c_417_n N_A_785_89#_c_967_n 0.00438365f $X=4.485 $Y=2.12 $X2=4.06
+ $Y2=2.48
cc_466 N_CK_c_427_n N_A_785_89#_c_967_n 0.00220762f $X=3.55 $Y=2.285 $X2=4.06
+ $Y2=2.48
cc_467 N_CK_c_439_n N_A_785_89#_c_967_n 0.0149594f $X=4.575 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_468 N_CK_c_441_n N_A_785_89#_c_967_n 0.0145646f $X=3.58 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_469 N_CK_c_444_n N_A_785_89#_c_967_n 0.0141886f $X=4.43 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_470 N_CK_c_445_n N_A_785_89#_c_967_n 0.00207435f $X=3.725 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_471 CK N_A_785_89#_c_967_n 0.00191287f $X=4.575 $Y=2.11 $X2=4.06 $Y2=2.48
cc_472 N_CK_c_416_n N_A_785_89#_c_974_n 0.00433036f $X=4.43 $Y=2.45 $X2=4.935
+ $Y2=2.48
cc_473 N_CK_M1017_g N_A_785_89#_c_974_n 0.00888384f $X=4.43 $Y=3.235 $X2=4.935
+ $Y2=2.48
cc_474 N_CK_c_439_n N_A_785_89#_c_974_n 0.00642476f $X=4.575 $Y=2.11 $X2=4.935
+ $Y2=2.48
cc_475 N_CK_c_444_n N_A_785_89#_c_974_n 0.0190758f $X=4.43 $Y=2.11 $X2=4.935
+ $Y2=2.48
cc_476 CK N_A_785_89#_c_974_n 0.025144f $X=4.575 $Y=2.11 $X2=4.935 $Y2=2.48
cc_477 N_CK_c_416_n N_A_785_89#_c_975_n 4.83733e-19 $X=4.43 $Y=2.45 $X2=4.205
+ $Y2=2.48
cc_478 N_CK_M1017_g N_A_785_89#_c_975_n 4.63789e-19 $X=4.43 $Y=3.235 $X2=4.205
+ $Y2=2.48
cc_479 N_CK_c_427_n N_A_785_89#_c_975_n 0.00406973f $X=3.55 $Y=2.285 $X2=4.205
+ $Y2=2.48
cc_480 N_CK_c_439_n N_A_785_89#_c_975_n 7.97287e-19 $X=4.575 $Y=2.11 $X2=4.205
+ $Y2=2.48
cc_481 N_CK_c_441_n N_A_785_89#_c_975_n 0.00250268f $X=3.58 $Y=2.11 $X2=4.205
+ $Y2=2.48
cc_482 N_CK_c_444_n N_A_785_89#_c_975_n 0.0252575f $X=4.43 $Y=2.11 $X2=4.205
+ $Y2=2.48
cc_483 N_CK_c_439_n N_A_785_89#_c_976_n 0.00120049f $X=4.575 $Y=2.11 $X2=5.007
+ $Y2=2.395
cc_484 CK N_A_785_89#_c_976_n 0.0189169f $X=4.575 $Y=2.11 $X2=5.007 $Y2=2.395
cc_485 N_CK_c_416_n N_A_623_115#_M1023_g 0.00468822f $X=4.43 $Y=2.45 $X2=5.38
+ $Y2=3.235
cc_486 N_CK_c_433_n N_A_623_115#_c_1122_n 0.00711103f $X=4.457 $Y=1.355 $X2=5.38
+ $Y2=1.4
cc_487 N_CK_c_423_n N_A_623_115#_c_1124_n 0.0018894f $X=3.1 $Y=1.4 $X2=2.76
+ $Y2=1.37
cc_488 N_CK_c_436_n N_A_623_115#_c_1124_n 0.0516585f $X=3.1 $Y=1.4 $X2=2.76
+ $Y2=1.37
cc_489 N_CK_c_438_n N_A_623_115#_c_1124_n 0.0116464f $X=3.185 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_490 N_CK_c_441_n N_A_623_115#_c_1124_n 0.00640739f $X=3.58 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_491 N_CK_c_442_n N_A_623_115#_c_1124_n 0.020359f $X=3.435 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_492 N_CK_c_445_n N_A_623_115#_c_1124_n 5.47744e-19 $X=3.725 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_493 N_CK_c_427_n N_A_623_115#_c_1154_n 0.00248712f $X=3.55 $Y=2.285 $X2=3.17
+ $Y2=2.705
cc_494 N_CK_c_437_n N_A_623_115#_c_1154_n 0.007489f $X=3.465 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_495 N_CK_c_438_n N_A_623_115#_c_1154_n 0.00323798f $X=3.185 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_496 N_CK_c_441_n N_A_623_115#_c_1154_n 0.00351845f $X=3.58 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_497 N_CK_c_442_n N_A_623_115#_c_1154_n 0.0125804f $X=3.435 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_498 N_CK_c_445_n N_A_623_115#_c_1154_n 8.86004e-19 $X=3.725 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_499 N_CK_c_423_n N_A_623_115#_c_1125_n 0.00131946f $X=3.1 $Y=1.4 $X2=3.44
+ $Y2=1.34
cc_500 N_CK_c_424_n N_A_623_115#_c_1125_n 0.00403992f $X=3.1 $Y=1.235 $X2=3.44
+ $Y2=1.34
cc_501 N_CK_c_436_n N_A_623_115#_c_1125_n 0.014622f $X=3.1 $Y=1.4 $X2=3.44
+ $Y2=1.34
cc_502 N_CK_c_437_n N_A_623_115#_c_1125_n 0.00112312f $X=3.465 $Y=2.11 $X2=3.44
+ $Y2=1.34
cc_503 N_CK_c_442_n N_A_623_115#_c_1125_n 9.66728e-19 $X=3.435 $Y=2.11 $X2=3.44
+ $Y2=1.34
cc_504 N_CK_c_423_n N_A_623_115#_c_1126_n 0.00217193f $X=3.1 $Y=1.4 $X2=3.34
+ $Y2=0.755
cc_505 N_CK_c_436_n N_A_623_115#_c_1126_n 8.41917e-19 $X=3.1 $Y=1.4 $X2=3.34
+ $Y2=0.755
cc_506 N_CK_c_423_n N_A_623_115#_c_1131_n 0.00611127f $X=3.1 $Y=1.4 $X2=3.295
+ $Y2=1.37
cc_507 N_CK_c_436_n N_A_623_115#_c_1131_n 0.0178129f $X=3.1 $Y=1.4 $X2=3.295
+ $Y2=1.37
cc_508 N_CK_c_437_n N_A_623_115#_c_1131_n 0.00291459f $X=3.465 $Y=2.11 $X2=3.295
+ $Y2=1.37
cc_509 N_CK_c_423_n N_A_623_115#_c_1132_n 6.81488e-19 $X=3.1 $Y=1.4 $X2=2.905
+ $Y2=1.37
cc_510 N_CK_c_436_n N_A_623_115#_c_1132_n 0.00134743f $X=3.1 $Y=1.4 $X2=2.905
+ $Y2=1.37
cc_511 N_CK_c_442_n N_A_623_115#_c_1132_n 0.0128239f $X=3.435 $Y=2.11 $X2=2.905
+ $Y2=1.37
cc_512 N_CK_c_417_n N_A_623_115#_c_1133_n 0.00322503f $X=4.485 $Y=2.12 $X2=5.03
+ $Y2=1.37
cc_513 N_CK_c_433_n N_A_623_115#_c_1133_n 0.0102398f $X=4.457 $Y=1.355 $X2=5.03
+ $Y2=1.37
cc_514 N_CK_c_423_n N_A_623_115#_c_1135_n 5.48392e-19 $X=3.1 $Y=1.4 $X2=3.585
+ $Y2=1.37
cc_515 N_CK_c_436_n N_A_623_115#_c_1135_n 8.69968e-19 $X=3.1 $Y=1.4 $X2=3.585
+ $Y2=1.37
cc_516 N_A_32_115#_c_665_n N_A_243_89#_c_762_n 0.00256272f $X=2.185 $Y=1.37
+ $X2=1.41 $Y2=1.775
cc_517 N_A_32_115#_c_665_n N_A_243_89#_c_763_n 0.00290011f $X=2.185 $Y=1.37
+ $X2=1.815 $Y2=1.85
cc_518 N_A_32_115#_c_652_n N_A_243_89#_M1011_g 0.113994f $X=2.325 $Y=2.285
+ $X2=1.89 $Y2=3.235
cc_519 N_A_32_115#_c_661_n N_A_243_89#_M1011_g 0.00435172f $X=2.42 $Y=2.285
+ $X2=1.89 $Y2=3.235
cc_520 N_A_32_115#_c_650_n N_A_243_89#_c_766_n 0.0342442f $X=2.325 $Y=1.4
+ $X2=2.965 $Y2=1.85
cc_521 N_A_32_115#_c_652_n N_A_243_89#_c_766_n 0.0355605f $X=2.325 $Y=2.285
+ $X2=2.965 $Y2=1.85
cc_522 N_A_32_115#_c_661_n N_A_243_89#_c_766_n 0.0111197f $X=2.42 $Y=2.285
+ $X2=2.965 $Y2=1.85
cc_523 N_A_32_115#_c_663_n N_A_243_89#_c_766_n 8.22237e-19 $X=2.42 $Y=1.4
+ $X2=2.965 $Y2=1.85
cc_524 N_A_32_115#_c_665_n N_A_243_89#_c_766_n 0.00477469f $X=2.185 $Y=1.37
+ $X2=2.965 $Y2=1.85
cc_525 N_A_32_115#_c_668_n N_A_243_89#_c_766_n 3.93645e-19 $X=2.33 $Y=1.37
+ $X2=2.965 $Y2=1.85
cc_526 N_A_32_115#_c_651_n N_A_243_89#_M1003_g 0.110621f $X=2.605 $Y=2.285
+ $X2=3.04 $Y2=3.235
cc_527 N_A_32_115#_M1004_g N_A_623_115#_c_1124_n 9.36754e-19 $X=2.25 $Y=3.235
+ $X2=2.76 $Y2=1.37
cc_528 N_A_32_115#_c_648_n N_A_623_115#_c_1124_n 0.0077615f $X=2.605 $Y=1.4
+ $X2=2.76 $Y2=1.37
cc_529 N_A_32_115#_c_651_n N_A_623_115#_c_1124_n 0.00729195f $X=2.605 $Y=2.285
+ $X2=2.76 $Y2=1.37
cc_530 N_A_32_115#_M1006_g N_A_623_115#_c_1124_n 0.00479454f $X=2.68 $Y=3.235
+ $X2=2.76 $Y2=1.37
cc_531 N_A_32_115#_c_661_n N_A_623_115#_c_1124_n 0.0700092f $X=2.42 $Y=2.285
+ $X2=2.76 $Y2=1.37
cc_532 N_A_32_115#_c_663_n N_A_623_115#_c_1124_n 0.0104545f $X=2.42 $Y=1.4
+ $X2=2.76 $Y2=1.37
cc_533 N_A_32_115#_c_668_n N_A_623_115#_c_1124_n 3.63286e-19 $X=2.33 $Y=1.37
+ $X2=2.76 $Y2=1.37
cc_534 N_A_32_115#_M1004_g N_A_623_115#_c_1184_n 9.13132e-19 $X=2.25 $Y=3.235
+ $X2=2.845 $Y2=2.705
cc_535 N_A_32_115#_M1006_g N_A_623_115#_c_1184_n 0.0096885f $X=2.68 $Y=3.235
+ $X2=2.845 $Y2=2.705
cc_536 N_A_32_115#_c_648_n N_A_623_115#_c_1132_n 0.00169405f $X=2.605 $Y=1.4
+ $X2=2.905 $Y2=1.37
cc_537 N_A_32_115#_M1015_g N_A_623_115#_c_1132_n 0.00605065f $X=2.68 $Y=0.85
+ $X2=2.905 $Y2=1.37
cc_538 N_A_32_115#_c_663_n N_A_623_115#_c_1132_n 0.00135424f $X=2.42 $Y=1.4
+ $X2=2.905 $Y2=1.37
cc_539 N_A_32_115#_c_668_n N_A_623_115#_c_1132_n 0.0241344f $X=2.33 $Y=1.37
+ $X2=2.905 $Y2=1.37
cc_540 N_A_243_89#_M1005_g N_A_785_89#_M1000_g 0.0470074f $X=3.64 $Y=0.85 $X2=4
+ $Y2=0.85
cc_541 N_A_243_89#_c_775_n N_A_785_89#_c_962_n 0.0470074f $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_542 N_A_243_89#_c_776_n N_A_785_89#_c_962_n 8.11121e-19 $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_543 N_A_243_89#_c_782_n N_A_785_89#_c_962_n 5.33708e-19 $X=4.645 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_544 N_A_243_89#_c_783_n N_A_785_89#_c_962_n 9.00828e-19 $X=3.725 $Y=1.725
+ $X2=4.06 $Y2=1.74
cc_545 N_A_243_89#_c_784_n N_A_785_89#_c_962_n 4.49351e-19 $X=4.645 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_546 N_A_243_89#_c_785_n N_A_785_89#_c_962_n 0.00295157f $X=4.5 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_547 N_A_243_89#_c_775_n N_A_785_89#_c_966_n 7.48149e-19 $X=3.58 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_548 N_A_243_89#_c_776_n N_A_785_89#_c_966_n 0.0079274f $X=3.58 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_549 N_A_243_89#_c_777_n N_A_785_89#_c_966_n 0.00254242f $X=4.645 $Y=0.755
+ $X2=4.062 $Y2=1.812
cc_550 N_A_243_89#_c_782_n N_A_785_89#_c_966_n 0.00340323f $X=4.645 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_551 N_A_243_89#_c_783_n N_A_785_89#_c_966_n 0.00135239f $X=3.725 $Y=1.725
+ $X2=4.062 $Y2=1.812
cc_552 N_A_243_89#_c_784_n N_A_785_89#_c_966_n 0.00101182f $X=4.645 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_553 N_A_243_89#_c_785_n N_A_785_89#_c_966_n 0.0115044f $X=4.5 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_554 N_A_243_89#_c_775_n N_A_785_89#_c_967_n 6.69855e-19 $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_555 N_A_243_89#_c_776_n N_A_785_89#_c_967_n 6.26362e-19 $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_556 N_A_243_89#_c_782_n N_A_785_89#_c_967_n 7.11909e-19 $X=4.645 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_557 N_A_243_89#_c_783_n N_A_785_89#_c_967_n 0.00136024f $X=3.725 $Y=1.725
+ $X2=4.06 $Y2=2.48
cc_558 N_A_243_89#_c_784_n N_A_785_89#_c_967_n 9.62563e-19 $X=4.645 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_559 N_A_243_89#_c_781_n N_A_785_89#_c_971_n 0.0162069f $X=4.915 $Y=2.62
+ $X2=5.595 $Y2=2.955
cc_560 N_A_243_89#_c_782_n N_A_785_89#_c_971_n 6.20209e-19 $X=4.645 $Y=1.74
+ $X2=5.595 $Y2=2.955
cc_561 N_A_243_89#_c_782_n N_A_785_89#_c_973_n 0.0038586f $X=4.645 $Y=1.74
+ $X2=5.595 $Y2=1.74
cc_562 N_A_243_89#_c_781_n N_A_785_89#_c_974_n 0.0170279f $X=4.915 $Y=2.62
+ $X2=4.935 $Y2=2.48
cc_563 N_A_243_89#_c_797_n N_A_785_89#_c_974_n 0.0134665f $X=4.915 $Y=2.705
+ $X2=4.935 $Y2=2.48
cc_564 N_A_243_89#_c_782_n N_A_785_89#_c_974_n 0.00186509f $X=4.645 $Y=1.74
+ $X2=4.935 $Y2=2.48
cc_565 N_A_243_89#_c_784_n N_A_785_89#_c_974_n 0.0032354f $X=4.645 $Y=1.74
+ $X2=4.935 $Y2=2.48
cc_566 N_A_243_89#_c_781_n N_A_785_89#_c_976_n 0.0176818f $X=4.915 $Y=2.62
+ $X2=5.007 $Y2=2.395
cc_567 N_A_243_89#_c_782_n N_A_785_89#_c_976_n 9.38674e-19 $X=4.645 $Y=1.74
+ $X2=5.007 $Y2=2.395
cc_568 N_A_243_89#_c_782_n N_A_785_89#_c_978_n 0.00750891f $X=4.645 $Y=1.74
+ $X2=5.08 $Y2=1.74
cc_569 N_A_243_89#_c_784_n N_A_785_89#_c_978_n 0.0197438f $X=4.645 $Y=1.74
+ $X2=5.08 $Y2=1.74
cc_570 N_A_243_89#_c_777_n N_A_623_115#_c_1117_n 0.00729796f $X=4.645 $Y=0.755
+ $X2=5.38 $Y2=1.235
cc_571 N_A_243_89#_c_777_n N_A_623_115#_M1023_g 0.00186304f $X=4.645 $Y=0.755
+ $X2=5.38 $Y2=3.235
cc_572 N_A_243_89#_c_792_n N_A_623_115#_M1023_g 0.00781432f $X=4.645 $Y=2.955
+ $X2=5.38 $Y2=3.235
cc_573 N_A_243_89#_c_781_n N_A_623_115#_M1023_g 0.0105293f $X=4.915 $Y=2.62
+ $X2=5.38 $Y2=3.235
cc_574 N_A_243_89#_c_797_n N_A_623_115#_M1023_g 0.00340068f $X=4.915 $Y=2.705
+ $X2=5.38 $Y2=3.235
cc_575 N_A_243_89#_c_782_n N_A_623_115#_M1023_g 0.00296549f $X=4.645 $Y=1.74
+ $X2=5.38 $Y2=3.235
cc_576 N_A_243_89#_c_784_n N_A_623_115#_M1023_g 5.83966e-19 $X=4.645 $Y=1.74
+ $X2=5.38 $Y2=3.235
cc_577 N_A_243_89#_c_777_n N_A_623_115#_c_1122_n 0.00323378f $X=4.645 $Y=0.755
+ $X2=5.38 $Y2=1.4
cc_578 N_A_243_89#_c_766_n N_A_623_115#_c_1124_n 0.0121637f $X=2.965 $Y=1.85
+ $X2=2.76 $Y2=1.37
cc_579 N_A_243_89#_M1003_g N_A_623_115#_c_1124_n 0.0104621f $X=3.04 $Y=3.235
+ $X2=2.76 $Y2=1.37
cc_580 N_A_243_89#_c_766_n N_A_623_115#_c_1154_n 5.88705e-19 $X=2.965 $Y=1.85
+ $X2=3.17 $Y2=2.705
cc_581 N_A_243_89#_M1003_g N_A_623_115#_c_1154_n 0.0162544f $X=3.04 $Y=3.235
+ $X2=3.17 $Y2=2.705
cc_582 N_A_243_89#_c_768_n N_A_623_115#_c_1154_n 6.306e-19 $X=3.445 $Y=1.85
+ $X2=3.17 $Y2=2.705
cc_583 N_A_243_89#_M1005_g N_A_623_115#_c_1125_n 0.0111789f $X=3.64 $Y=0.85
+ $X2=3.44 $Y2=1.34
cc_584 N_A_243_89#_c_775_n N_A_623_115#_c_1125_n 0.0019278f $X=3.58 $Y=1.74
+ $X2=3.44 $Y2=1.34
cc_585 N_A_243_89#_c_776_n N_A_623_115#_c_1125_n 0.00649516f $X=3.58 $Y=1.74
+ $X2=3.44 $Y2=1.34
cc_586 N_A_243_89#_c_783_n N_A_623_115#_c_1125_n 3.68943e-19 $X=3.725 $Y=1.725
+ $X2=3.44 $Y2=1.34
cc_587 N_A_243_89#_c_777_n N_A_623_115#_c_1129_n 0.00848647f $X=4.645 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_588 N_A_243_89#_c_766_n N_A_623_115#_c_1131_n 0.0015396f $X=2.965 $Y=1.85
+ $X2=3.295 $Y2=1.37
cc_589 N_A_243_89#_c_768_n N_A_623_115#_c_1131_n 0.00243388f $X=3.445 $Y=1.85
+ $X2=3.295 $Y2=1.37
cc_590 N_A_243_89#_c_774_n N_A_623_115#_c_1131_n 5.01668e-19 $X=3.04 $Y=1.85
+ $X2=3.295 $Y2=1.37
cc_591 N_A_243_89#_c_766_n N_A_623_115#_c_1132_n 0.00117411f $X=2.965 $Y=1.85
+ $X2=2.905 $Y2=1.37
cc_592 N_A_243_89#_M1005_g N_A_623_115#_c_1133_n 0.0076805f $X=3.64 $Y=0.85
+ $X2=5.03 $Y2=1.37
cc_593 N_A_243_89#_c_777_n N_A_623_115#_c_1133_n 0.0231229f $X=4.645 $Y=0.755
+ $X2=5.03 $Y2=1.37
cc_594 N_A_243_89#_c_782_n N_A_623_115#_c_1133_n 0.0081736f $X=4.645 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_595 N_A_243_89#_c_784_n N_A_623_115#_c_1133_n 0.0251744f $X=4.645 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_596 N_A_243_89#_c_785_n N_A_623_115#_c_1133_n 0.0641247f $X=4.5 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_597 N_A_243_89#_M1005_g N_A_623_115#_c_1135_n 0.00332547f $X=3.64 $Y=0.85
+ $X2=3.585 $Y2=1.37
cc_598 N_A_243_89#_c_775_n N_A_623_115#_c_1135_n 6.54323e-19 $X=3.58 $Y=1.74
+ $X2=3.585 $Y2=1.37
cc_599 N_A_243_89#_c_776_n N_A_623_115#_c_1135_n 0.00311003f $X=3.58 $Y=1.74
+ $X2=3.585 $Y2=1.37
cc_600 N_A_243_89#_c_783_n N_A_623_115#_c_1135_n 0.0279665f $X=3.725 $Y=1.725
+ $X2=3.585 $Y2=1.37
cc_601 N_A_243_89#_c_777_n N_A_623_115#_c_1136_n 0.00149153f $X=4.645 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_602 N_A_785_89#_c_968_n N_A_623_115#_c_1117_n 0.0212717f $X=5.595 $Y=0.755
+ $X2=5.38 $Y2=1.235
cc_603 N_A_785_89#_c_957_n N_A_623_115#_M1023_g 0.00462538f $X=6.28 $Y=1.905
+ $X2=5.38 $Y2=3.235
cc_604 N_A_785_89#_c_971_n N_A_623_115#_M1023_g 0.0232766f $X=5.595 $Y=2.955
+ $X2=5.38 $Y2=3.235
cc_605 N_A_785_89#_c_973_n N_A_623_115#_M1023_g 0.0024326f $X=5.595 $Y=1.74
+ $X2=5.38 $Y2=3.235
cc_606 N_A_785_89#_c_976_n N_A_623_115#_M1023_g 0.0141612f $X=5.007 $Y=2.395
+ $X2=5.38 $Y2=3.235
cc_607 N_A_785_89#_c_977_n N_A_623_115#_M1023_g 0.0162618f $X=6.08 $Y=1.74
+ $X2=5.38 $Y2=3.235
cc_608 N_A_785_89#_c_978_n N_A_623_115#_c_1122_n 0.00424614f $X=5.08 $Y=1.74
+ $X2=5.38 $Y2=1.4
cc_609 N_A_785_89#_c_968_n N_A_623_115#_c_1129_n 0.012913f $X=5.595 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_610 N_A_785_89#_c_977_n N_A_623_115#_c_1129_n 7.77735e-19 $X=6.08 $Y=1.74
+ $X2=5.175 $Y2=1.37
cc_611 N_A_785_89#_c_978_n N_A_623_115#_c_1129_n 0.004937f $X=5.08 $Y=1.74
+ $X2=5.175 $Y2=1.37
cc_612 N_A_785_89#_M1000_g N_A_623_115#_c_1133_n 0.0105151f $X=4 $Y=0.85
+ $X2=5.03 $Y2=1.37
cc_613 N_A_785_89#_c_962_n N_A_623_115#_c_1133_n 7.90759e-19 $X=4.06 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_614 N_A_785_89#_c_966_n N_A_623_115#_c_1133_n 0.00516488f $X=4.062 $Y=1.812
+ $X2=5.03 $Y2=1.37
cc_615 N_A_785_89#_c_978_n N_A_623_115#_c_1133_n 0.0082117f $X=5.08 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_616 N_A_785_89#_c_968_n N_A_623_115#_c_1136_n 0.0033865f $X=5.595 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_617 N_A_785_89#_c_978_n N_A_623_115#_c_1136_n 0.0258498f $X=5.08 $Y=1.74
+ $X2=5.175 $Y2=1.37
cc_618 N_A_785_89#_c_957_n N_ON_M1002_g 0.0154305f $X=6.28 $Y=1.905 $X2=6.76
+ $Y2=0.85
cc_619 N_A_785_89#_M1010_g N_ON_M1002_g 0.0253877f $X=6.33 $Y=0.85 $X2=6.76
+ $Y2=0.85
cc_620 N_A_785_89#_c_972_n N_ON_M1002_g 6.55283e-19 $X=6.215 $Y=1.74 $X2=6.76
+ $Y2=0.85
cc_621 N_A_785_89#_c_964_n N_ON_M1018_g 0.00630133f $X=6.305 $Y=2.36 $X2=6.76
+ $Y2=3.235
cc_622 N_A_785_89#_c_965_n N_ON_M1018_g 0.0506162f $X=6.305 $Y=2.49 $X2=6.76
+ $Y2=3.235
cc_623 N_A_785_89#_c_957_n N_ON_c_1244_n 0.0212297f $X=6.28 $Y=1.905 $X2=6.7
+ $Y2=2.015
cc_624 N_A_785_89#_c_957_n N_ON_c_1245_n 0.00188672f $X=6.28 $Y=1.905 $X2=6.115
+ $Y2=0.74
cc_625 N_A_785_89#_M1010_g N_ON_c_1245_n 0.00922835f $X=6.33 $Y=0.85 $X2=6.115
+ $Y2=0.74
cc_626 N_A_785_89#_c_968_n N_ON_c_1245_n 0.0321547f $X=5.595 $Y=0.755 $X2=6.115
+ $Y2=0.74
cc_627 N_A_785_89#_c_957_n N_ON_c_1248_n 0.00289364f $X=6.28 $Y=1.905 $X2=6.115
+ $Y2=2.195
cc_628 N_A_785_89#_c_971_n N_ON_c_1248_n 0.00525727f $X=5.595 $Y=2.955 $X2=6.115
+ $Y2=2.195
cc_629 N_A_785_89#_c_972_n N_ON_c_1248_n 0.0101349f $X=6.215 $Y=1.74 $X2=6.115
+ $Y2=2.195
cc_630 N_A_785_89#_c_979_n N_ON_c_1248_n 3.37612e-19 $X=6.215 $Y=1.74 $X2=6.115
+ $Y2=2.195
cc_631 N_A_785_89#_c_964_n N_ON_c_1249_n 0.0120965f $X=6.305 $Y=2.36 $X2=6.115
+ $Y2=3.615
cc_632 N_A_785_89#_c_965_n N_ON_c_1249_n 0.0210894f $X=6.305 $Y=2.49 $X2=6.115
+ $Y2=3.615
cc_633 N_A_785_89#_c_971_n N_ON_c_1249_n 0.0721092f $X=5.595 $Y=2.955 $X2=6.115
+ $Y2=3.615
cc_634 N_A_785_89#_c_957_n N_ON_c_1250_n 0.0192889f $X=6.28 $Y=1.905 $X2=6.615
+ $Y2=1.4
cc_635 N_A_785_89#_c_972_n N_ON_c_1250_n 0.0110497f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=1.4
cc_636 N_A_785_89#_c_979_n N_ON_c_1250_n 0.00387586f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=1.4
cc_637 N_A_785_89#_c_957_n N_ON_c_1252_n 0.00308111f $X=6.28 $Y=1.905 $X2=6.2
+ $Y2=1.4
cc_638 N_A_785_89#_c_968_n N_ON_c_1252_n 0.00869401f $X=5.595 $Y=0.755 $X2=6.2
+ $Y2=1.4
cc_639 N_A_785_89#_c_972_n N_ON_c_1252_n 0.0120752f $X=6.215 $Y=1.74 $X2=6.2
+ $Y2=1.4
cc_640 N_A_785_89#_c_977_n N_ON_c_1252_n 0.00132729f $X=6.08 $Y=1.74 $X2=6.2
+ $Y2=1.4
cc_641 N_A_785_89#_c_979_n N_ON_c_1252_n 0.00306734f $X=6.215 $Y=1.74 $X2=6.2
+ $Y2=1.4
cc_642 N_A_785_89#_c_957_n N_ON_c_1253_n 2.65797e-19 $X=6.28 $Y=1.905 $X2=6.615
+ $Y2=2.11
cc_643 N_A_785_89#_c_964_n N_ON_c_1253_n 0.0141863f $X=6.305 $Y=2.36 $X2=6.615
+ $Y2=2.11
cc_644 N_A_785_89#_c_965_n N_ON_c_1253_n 0.00208656f $X=6.305 $Y=2.49 $X2=6.615
+ $Y2=2.11
cc_645 N_A_785_89#_c_972_n N_ON_c_1253_n 0.00957264f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=2.11
cc_646 N_A_785_89#_c_979_n N_ON_c_1253_n 0.00261089f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=2.11
cc_647 N_A_785_89#_c_957_n N_ON_c_1254_n 0.00380215f $X=6.28 $Y=1.905 $X2=6.702
+ $Y2=1.658
cc_648 N_A_785_89#_c_972_n N_ON_c_1254_n 0.00996181f $X=6.215 $Y=1.74 $X2=6.702
+ $Y2=1.658
cc_649 N_A_785_89#_c_979_n N_ON_c_1254_n 0.00251327f $X=6.215 $Y=1.74 $X2=6.702
+ $Y2=1.658
cc_650 N_A_785_89#_c_957_n N_ON_c_1255_n 0.00152939f $X=6.28 $Y=1.905 $X2=6.7
+ $Y2=2.015
cc_651 N_A_785_89#_c_979_n N_ON_c_1255_n 0.00137139f $X=6.215 $Y=1.74 $X2=6.7
+ $Y2=2.015
cc_652 N_A_785_89#_c_957_n ON 0.00197254f $X=6.28 $Y=1.905 $X2=6.115 $Y2=2.11
cc_653 N_A_785_89#_c_964_n ON 0.0039793f $X=6.305 $Y=2.36 $X2=6.115 $Y2=2.11
cc_654 N_A_785_89#_c_971_n ON 0.00761812f $X=5.595 $Y=2.955 $X2=6.115 $Y2=2.11
cc_655 N_A_785_89#_c_972_n ON 0.00222181f $X=6.215 $Y=1.74 $X2=6.115 $Y2=2.11
cc_656 N_A_785_89#_c_977_n ON 0.0192933f $X=6.08 $Y=1.74 $X2=6.115 $Y2=2.11
cc_657 N_A_785_89#_c_979_n ON 0.0183431f $X=6.215 $Y=1.74 $X2=6.115 $Y2=2.11
cc_658 N_A_785_89#_c_965_n Q 0.0010185f $X=6.305 $Y=2.49 $X2=6.97 $Y2=2.48
cc_659 N_A_623_115#_c_1154_n A_551_521# 0.0031646f $X=3.17 $Y=2.705 $X2=2.755
+ $Y2=2.605
cc_660 N_A_623_115#_c_1184_n A_551_521# 0.00144354f $X=2.845 $Y=2.705 $X2=2.755
+ $Y2=2.605
cc_661 N_ON_M1002_g N_Q_c_1322_n 0.0301628f $X=6.76 $Y=0.85 $X2=7.09 $Y2=2.395
cc_662 N_ON_c_1250_n N_Q_c_1322_n 0.0113726f $X=6.615 $Y=1.4 $X2=7.09 $Y2=2.395
cc_663 N_ON_c_1253_n N_Q_c_1322_n 0.0111434f $X=6.615 $Y=2.11 $X2=7.09 $Y2=2.395
cc_664 N_ON_c_1254_n N_Q_c_1322_n 0.0155777f $X=6.702 $Y=1.658 $X2=7.09
+ $Y2=2.395
cc_665 N_ON_c_1255_n N_Q_c_1322_n 0.0164341f $X=6.7 $Y=2.015 $X2=7.09 $Y2=2.395
cc_666 N_ON_M1018_g N_Q_c_1323_n 0.00583168f $X=6.76 $Y=3.235 $X2=7.09 $Y2=2.48
cc_667 N_ON_M1018_g N_Q_c_1330_n 0.0123536f $X=6.76 $Y=3.235 $X2=6.972 $Y2=2.88
cc_668 N_ON_M1002_g N_Q_c_1324_n 0.00384319f $X=6.76 $Y=0.85 $X2=7.09 $Y2=1.07
cc_669 N_ON_M1018_g Q 0.0140528f $X=6.76 $Y=3.235 $X2=6.97 $Y2=2.48
cc_670 N_ON_c_1249_n Q 0.00550321f $X=6.115 $Y=3.615 $X2=6.97 $Y2=2.48
cc_671 N_ON_c_1253_n Q 0.00287022f $X=6.615 $Y=2.11 $X2=6.97 $Y2=2.48
