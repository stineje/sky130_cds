* File: sky130_osu_sc_18T_ls__inv_3.spice
* Created: Fri Nov 12 14:17:29 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_ls__inv_3.pex.spice"
.subckt sky130_osu_sc_18T_ls__inv_3  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1000 N_GND_M1000_d N_A_M1000_g N_Y_M1000_s N_GND_M1000_b NSHORT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1000_s N_GND_M1000_b NSHORT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_GND_M1001_d N_A_M1003_g N_Y_M1003_s N_GND_M1000_b NSHORT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VDD_M1002_s N_VDD_M1002_b PHIGHVT L=0.15 W=3
+ AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2 SB=75001
+ A=0.45 P=6.3 MULT=1
MM1004 N_Y_M1002_d N_A_M1004_g N_VDD_M1004_s N_VDD_M1002_b PHIGHVT L=0.15 W=3
+ AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75000.6
+ A=0.45 P=6.3 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VDD_M1004_s N_VDD_M1002_b PHIGHVT L=0.15 W=3
+ AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX6_noxref N_GND_M1000_b N_VDD_M1002_b NWDIODE A=7.296 P=11.44
pX7_noxref noxref_5 A A PROBETYPE=1
pX8_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__inv_3.pxi.spice"
*
.ends
*
*
