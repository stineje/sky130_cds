* File: sky130_osu_sc_15T_ls__nand2_1.pxi.spice
* Created: Fri Nov 12 14:58:21 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__NAND2_1%GND N_GND_M1001_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_9_p GND N_GND_c_3_p PM_SKY130_OSU_SC_15T_LS__NAND2_1%GND
x_PM_SKY130_OSU_SC_15T_LS__NAND2_1%VDD N_VDD_M1000_s N_VDD_M1003_d N_VDD_M1000_b
+ N_VDD_c_27_p N_VDD_c_28_p N_VDD_c_37_p VDD N_VDD_c_29_p
+ PM_SKY130_OSU_SC_15T_LS__NAND2_1%VDD
x_PM_SKY130_OSU_SC_15T_LS__NAND2_1%A N_A_M1002_g N_A_M1000_g N_A_c_50_n
+ N_A_c_51_n A PM_SKY130_OSU_SC_15T_LS__NAND2_1%A
x_PM_SKY130_OSU_SC_15T_LS__NAND2_1%B N_B_M1001_g N_B_M1003_g N_B_c_82_n
+ N_B_c_84_n N_B_c_85_n B PM_SKY130_OSU_SC_15T_LS__NAND2_1%B
x_PM_SKY130_OSU_SC_15T_LS__NAND2_1%Y N_Y_M1002_s N_Y_M1000_d N_Y_c_115_n
+ N_Y_c_118_n N_Y_c_119_n N_Y_c_120_n Y N_Y_c_123_n
+ PM_SKY130_OSU_SC_15T_LS__NAND2_1%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.0889283f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1002_b N_A_M1000_g 0.00342256f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_5 N_GND_M1002_b N_A_c_50_n 0.0490341f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.425
cc_6 N_GND_M1002_b N_A_c_51_n 0.00856875f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.425
cc_7 N_GND_M1002_b N_B_M1001_g 0.0461967f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_8 N_GND_c_2_p N_B_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.945
cc_9 N_GND_c_9_p N_B_M1001_g 0.00866533f $X=1.05 $Y=0.865 $X2=0.835 $Y2=0.945
cc_10 N_GND_c_3_p N_B_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.945
cc_11 N_GND_M1002_b N_B_M1003_g 0.0316271f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_12 N_GND_M1002_b N_B_c_82_n 0.0353546f $X=-0.045 $Y=0 $X2=0.915 $Y2=1.96
cc_13 N_GND_c_9_p N_B_c_82_n 0.00231535f $X=1.05 $Y=0.865 $X2=0.915 $Y2=1.96
cc_14 N_GND_M1002_b N_B_c_84_n 0.0195876f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.7
cc_15 N_GND_M1002_b N_B_c_85_n 0.0122574f $X=-0.045 $Y=0 $X2=1.06 $Y2=1.96
cc_16 N_GND_M1002_b B 0.00492682f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.7
cc_17 N_GND_M1002_b N_Y_c_115_n 0.00156053f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.865
cc_18 N_GND_c_2_p N_Y_c_115_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26 $Y2=0.865
cc_19 N_GND_c_3_p N_Y_c_115_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26 $Y2=0.865
cc_20 N_GND_M1002_b N_Y_c_118_n 0.00851145f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.33
cc_21 N_GND_c_9_p N_Y_c_119_n 6.82281e-19 $X=1.05 $Y=0.865 $X2=0.605 $Y2=1.22
cc_22 N_GND_M1002_b N_Y_c_120_n 0.0206417f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.22
cc_23 N_GND_c_9_p N_Y_c_120_n 5.67165e-19 $X=1.05 $Y=0.865 $X2=0.405 $Y2=1.22
cc_24 N_GND_M1002_b Y 0.013296f $X=-0.045 $Y=0 $X2=0.68 $Y2=2.09
cc_25 N_GND_M1002_b N_Y_c_123_n 0.00518799f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.33
cc_26 N_VDD_M1000_b N_A_M1000_g 0.0229548f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_27 N_VDD_c_27_p N_A_M1000_g 0.00751602f $X=0.26 $Y=3.885 $X2=0.475 $Y2=3.825
cc_28 N_VDD_c_28_p N_A_M1000_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475 $Y2=3.825
cc_29 N_VDD_c_29_p N_A_M1000_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=3.825
cc_30 N_VDD_M1000_s N_A_c_51_n 0.00953431f $X=0.135 $Y=2.825 $X2=0.32 $Y2=2.425
cc_31 N_VDD_M1000_b N_A_c_51_n 0.00618364f $X=-0.045 $Y=2.645 $X2=0.32 $Y2=2.425
cc_32 N_VDD_c_27_p N_A_c_51_n 0.00252874f $X=0.26 $Y=3.885 $X2=0.32 $Y2=2.425
cc_33 N_VDD_M1000_s A 0.0150401f $X=0.135 $Y=2.825 $X2=0.32 $Y2=3.07
cc_34 N_VDD_c_27_p A 0.00522047f $X=0.26 $Y=3.885 $X2=0.32 $Y2=3.07
cc_35 N_VDD_M1000_b N_B_M1003_g 0.0226242f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_36 N_VDD_c_28_p N_B_M1003_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905 $Y2=3.825
cc_37 N_VDD_c_37_p N_B_M1003_g 0.00751602f $X=1.12 $Y=3.545 $X2=0.905 $Y2=3.825
cc_38 N_VDD_c_29_p N_B_M1003_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.905 $Y2=3.825
cc_39 N_VDD_M1000_b N_B_c_84_n 0.00337476f $X=-0.045 $Y=2.645 $X2=1.06 $Y2=2.7
cc_40 N_VDD_c_37_p N_B_c_84_n 0.00252359f $X=1.12 $Y=3.545 $X2=1.06 $Y2=2.7
cc_41 N_VDD_M1000_b B 0.012337f $X=-0.045 $Y=2.645 $X2=1.06 $Y2=2.7
cc_42 N_VDD_c_37_p B 0.00509939f $X=1.12 $Y=3.545 $X2=1.06 $Y2=2.7
cc_43 N_VDD_M1000_b N_Y_c_118_n 0.00501659f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.33
cc_44 N_VDD_c_28_p N_Y_c_118_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69 $Y2=2.33
cc_45 N_VDD_c_29_p N_Y_c_118_n 0.00434939f $X=1.02 $Y=5.36 $X2=0.69 $Y2=2.33
cc_46 N_A_M1002_g N_B_M1001_g 0.105421f $X=0.475 $Y=0.945 $X2=0.835 $Y2=0.945
cc_47 N_A_M1002_g N_B_M1003_g 0.044872f $X=0.475 $Y=0.945 $X2=0.905 $Y2=3.825
cc_48 N_A_M1002_g N_B_c_84_n 0.00112963f $X=0.475 $Y=0.945 $X2=1.06 $Y2=2.7
cc_49 N_A_M1002_g N_B_c_85_n 0.00282768f $X=0.475 $Y=0.945 $X2=1.06 $Y2=1.96
cc_50 A N_Y_M1000_d 0.00263091f $X=0.32 $Y=3.07 $X2=0.55 $Y2=2.825
cc_51 N_A_M1002_g N_Y_c_115_n 0.00740756f $X=0.475 $Y=0.945 $X2=0.26 $Y2=0.865
cc_52 N_A_M1002_g N_Y_c_118_n 0.00554573f $X=0.475 $Y=0.945 $X2=0.69 $Y2=2.33
cc_53 N_A_c_51_n N_Y_c_118_n 0.0420549f $X=0.32 $Y=2.425 $X2=0.69 $Y2=2.33
cc_54 A N_Y_c_118_n 0.00831114f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.33
cc_55 N_A_M1002_g N_Y_c_119_n 0.0136921f $X=0.475 $Y=0.945 $X2=0.605 $Y2=1.22
cc_56 N_A_M1002_g N_Y_c_120_n 0.00380596f $X=0.475 $Y=0.945 $X2=0.405 $Y2=1.22
cc_57 N_A_M1002_g Y 0.0123501f $X=0.475 $Y=0.945 $X2=0.68 $Y2=2.09
cc_58 N_A_M1002_g N_Y_c_123_n 0.00216533f $X=0.475 $Y=0.945 $X2=0.69 $Y2=2.33
cc_59 N_A_c_50_n N_Y_c_123_n 0.00278592f $X=0.32 $Y=2.425 $X2=0.69 $Y2=2.33
cc_60 N_A_c_51_n N_Y_c_123_n 0.00474021f $X=0.32 $Y=2.425 $X2=0.69 $Y2=2.33
cc_61 A N_Y_c_123_n 0.00150969f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.33
cc_62 N_B_M1003_g N_Y_c_118_n 0.00568509f $X=0.905 $Y=3.825 $X2=0.69 $Y2=2.33
cc_63 N_B_c_82_n N_Y_c_118_n 2.88224e-19 $X=0.915 $Y=1.96 $X2=0.69 $Y2=2.33
cc_64 N_B_c_84_n N_Y_c_118_n 0.0295869f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_65 N_B_c_85_n N_Y_c_118_n 0.00144012f $X=1.06 $Y=1.96 $X2=0.69 $Y2=2.33
cc_66 B N_Y_c_118_n 0.00831114f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_67 N_B_M1001_g N_Y_c_119_n 0.00790819f $X=0.835 $Y=0.945 $X2=0.605 $Y2=1.22
cc_68 N_B_M1001_g Y 0.0185298f $X=0.835 $Y=0.945 $X2=0.68 $Y2=2.09
cc_69 N_B_M1003_g Y 0.00128442f $X=0.905 $Y=3.825 $X2=0.68 $Y2=2.09
cc_70 N_B_c_82_n Y 0.00398874f $X=0.915 $Y=1.96 $X2=0.68 $Y2=2.09
cc_71 N_B_c_84_n Y 0.0066619f $X=1.06 $Y=2.7 $X2=0.68 $Y2=2.09
cc_72 N_B_c_85_n Y 0.0139756f $X=1.06 $Y=1.96 $X2=0.68 $Y2=2.09
cc_73 N_B_M1003_g N_Y_c_123_n 0.00339349f $X=0.905 $Y=3.825 $X2=0.69 $Y2=2.33
cc_74 N_B_c_82_n N_Y_c_123_n 0.00170653f $X=0.915 $Y=1.96 $X2=0.69 $Y2=2.33
cc_75 N_B_c_84_n N_Y_c_123_n 0.00640429f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_76 N_B_c_85_n N_Y_c_123_n 0.00261701f $X=1.06 $Y=1.96 $X2=0.69 $Y2=2.33
cc_77 B N_Y_c_123_n 0.0028041f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_78 N_Y_c_119_n A_110_115# 0.0109071f $X=0.605 $Y=1.22 $X2=0.55 $Y2=0.575
