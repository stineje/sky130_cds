magic
tech sky130A
magscale 1 2
timestamp 1600380937
<< checkpaint >>
rect -1260 -1260 1261 1261
<< nwell >>
rect -9 581 814 1341
<< nmos >>
rect 80 115 110 315
rect 152 115 182 315
rect 252 115 282 315
rect 338 115 368 315
rect 424 115 454 315
rect 510 115 540 315
rect 596 115 626 315
rect 682 115 712 315
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
rect 338 617 368 1217
rect 424 617 454 1217
rect 510 617 540 1217
rect 596 617 626 1217
rect 682 617 712 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 115 152 315
rect 182 267 252 315
rect 182 131 193 267
rect 227 131 252 267
rect 182 115 252 131
rect 282 267 338 315
rect 282 131 293 267
rect 327 131 338 267
rect 282 115 338 131
rect 368 267 424 315
rect 368 131 379 267
rect 413 131 424 267
rect 368 115 424 131
rect 454 267 510 315
rect 454 131 465 267
rect 499 131 510 267
rect 454 115 510 131
rect 540 267 596 315
rect 540 131 551 267
rect 585 131 596 267
rect 540 115 596 131
rect 626 267 682 315
rect 626 131 637 267
rect 671 131 682 267
rect 626 115 682 131
rect 712 267 765 315
rect 712 131 723 267
rect 757 131 765 267
rect 712 115 765 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 166 1217
rect 110 725 121 1201
rect 155 725 166 1201
rect 110 617 166 725
rect 196 1201 252 1217
rect 196 725 207 1201
rect 241 725 252 1201
rect 196 617 252 725
rect 282 1201 338 1217
rect 282 657 293 1201
rect 327 657 338 1201
rect 282 617 338 657
rect 368 1201 424 1217
rect 368 657 379 1201
rect 413 657 424 1201
rect 368 617 424 657
rect 454 1201 510 1217
rect 454 657 465 1201
rect 499 657 510 1201
rect 454 617 510 657
rect 540 1201 596 1217
rect 540 657 551 1201
rect 585 657 596 1201
rect 540 617 596 657
rect 626 1201 682 1217
rect 626 657 637 1201
rect 671 657 682 1201
rect 626 617 682 657
rect 712 1201 765 1217
rect 712 657 723 1201
rect 757 657 765 1201
rect 712 617 765 657
<< ndiffc >>
rect 35 131 69 267
rect 193 131 227 267
rect 293 131 327 267
rect 379 131 413 267
rect 465 131 499 267
rect 551 131 585 267
rect 637 131 671 267
rect 723 131 757 267
<< pdiffc >>
rect 35 793 69 1201
rect 121 725 155 1201
rect 207 725 241 1201
rect 293 657 327 1201
rect 379 657 413 1201
rect 465 657 499 1201
rect 551 657 585 1201
rect 637 657 671 1201
rect 723 657 757 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 338 1217 368 1244
rect 424 1217 454 1243
rect 510 1217 540 1243
rect 596 1217 626 1243
rect 682 1217 712 1243
rect 80 586 110 617
rect 20 570 110 586
rect 20 536 30 570
rect 64 536 110 570
rect 20 520 110 536
rect 80 315 110 520
rect 166 519 196 617
rect 252 592 282 617
rect 338 592 368 617
rect 424 592 454 617
rect 510 592 540 617
rect 596 592 626 617
rect 682 592 712 617
rect 252 562 712 592
rect 152 502 210 519
rect 152 468 166 502
rect 200 468 210 502
rect 152 452 210 468
rect 152 315 182 452
rect 252 420 282 562
rect 252 404 306 420
rect 252 370 262 404
rect 296 384 306 404
rect 596 384 626 562
rect 296 370 712 384
rect 252 354 712 370
rect 252 315 282 354
rect 338 315 368 354
rect 424 315 454 354
rect 510 315 540 354
rect 596 315 626 354
rect 682 315 712 354
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
rect 338 89 368 115
rect 424 89 454 115
rect 510 89 540 115
rect 596 89 626 115
rect 682 89 712 115
<< polycont >>
rect 30 536 64 570
rect 166 468 200 502
rect 262 370 296 404
<< locali >>
rect 0 1305 814 1332
rect 0 1271 51 1305
rect 85 1271 187 1305
rect 221 1271 323 1305
rect 357 1271 459 1305
rect 493 1271 595 1305
rect 629 1271 814 1305
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 98 725 121 743
rect 98 709 155 725
rect 207 1201 241 1271
rect 207 709 241 725
rect 293 1201 327 1217
rect 30 570 64 649
rect 30 520 64 536
rect 98 404 132 709
rect 166 502 200 575
rect 293 535 327 657
rect 379 1201 413 1271
rect 379 641 413 657
rect 465 1201 499 1217
rect 465 535 499 657
rect 551 1201 585 1271
rect 551 641 585 657
rect 637 1201 671 1217
rect 637 535 671 657
rect 723 1201 757 1271
rect 723 641 757 657
rect 166 452 200 468
rect 35 370 262 404
rect 296 370 312 404
rect 35 267 69 370
rect 35 115 69 131
rect 193 267 227 283
rect 193 61 227 131
rect 293 267 327 279
rect 293 115 327 131
rect 379 267 413 283
rect 379 61 413 131
rect 465 267 499 279
rect 465 115 499 131
rect 551 267 585 283
rect 551 61 585 131
rect 637 267 671 279
rect 637 115 671 131
rect 723 267 757 283
rect 723 61 757 131
rect 0 27 51 61
rect 85 27 187 61
rect 221 27 323 61
rect 357 27 459 61
rect 493 27 595 61
rect 629 27 814 61
rect 0 0 814 27
<< viali >>
rect 30 649 64 683
rect 166 575 200 609
rect 293 501 327 535
rect 465 501 499 535
rect 637 501 671 535
rect 293 279 327 313
rect 465 279 499 313
rect 637 279 671 313
<< metal1 >>
rect 0 1271 814 1332
rect 18 683 76 689
rect 18 649 30 683
rect 64 649 98 683
rect 18 643 76 649
rect 154 609 212 615
rect 132 575 166 609
rect 200 575 212 609
rect 154 569 212 575
rect 281 535 339 541
rect 453 535 511 541
rect 625 535 683 541
rect 281 501 293 535
rect 327 501 465 535
rect 499 501 637 535
rect 671 501 683 535
rect 281 495 339 501
rect 453 495 511 501
rect 625 495 683 501
rect 293 319 327 495
rect 465 319 499 495
rect 637 319 671 495
rect 281 313 339 319
rect 453 313 511 319
rect 625 313 683 319
rect 281 279 293 313
rect 327 279 465 313
rect 499 279 637 313
rect 671 279 683 313
rect 281 273 339 279
rect 453 273 511 279
rect 625 273 683 279
rect 0 0 814 61
<< labels >>
rlabel metal1 68 44 68 44 1 gnd
rlabel metal1 68 1288 68 1288 1 vdd
rlabel metal1 184 592 184 592 1 B
port 1 n
rlabel metal1 48 666 48 666 1 A
port 2 n
rlabel metal1 311 444 311 444 1 Y
port 3 n
<< end >>
