* File: sky130_osu_sc_18T_hs__ant.pex.spice
* Created: Thu Oct 29 17:06:22 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__ANT%GND 5 11
r13 5 11 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=0.17 $X2=0.34
+ $Y2=0.17
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ANT%VDD 1 7 11 15 17
r7 17 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=6.49 $X2=0.34
+ $Y2=6.49
r8 15 23 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r9 11 14 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r10 9 15 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.605 $Y2=6.507
r11 9 14 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r12 7 23 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r13 1 14 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r14 1 11 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ANT%A 1 3 12 16 20 23 26 30 34 36 38 41 46
r20 46 48 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=2.59
+ $X2=0.362 $Y2=2.755
r21 46 47 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=2.59
+ $X2=0.362 $Y2=2.425
r22 41 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.59 $X2=0.32 $Y2=2.59
r23 38 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.59
+ $X2=0.32 $Y2=2.59
r24 32 34 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.69 $Y=1.915
+ $X2=0.69 $Y2=0.825
r25 31 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.26
+ $Y2=2
r26 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=2
+ $X2=0.69 $Y2=1.915
r27 30 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=2 $X2=0.345
+ $Y2=2
r28 26 28 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r29 24 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=2.59
r30 24 26 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=3.455
r31 23 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.505
+ $X2=0.26 $Y2=2.59
r32 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2
r33 22 23 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2.505
r34 18 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.915
+ $X2=0.26 $Y2=2
r35 18 20 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.26 $Y=1.915
+ $X2=0.26 $Y2=0.825
r36 16 48 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.755
r37 12 47 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.425
r38 3 28 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r39 3 26 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r40 1 34 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
r41 1 20 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

