magic
tech sky130A
magscale 1 2
timestamp 1606864597
<< checkpaint >>
rect -801 1315 1753 2575
rect -1209 -1243 1753 1315
<< nwell >>
rect -9 581 553 1341
<< nmos >>
rect 80 115 110 315
rect 270 115 300 315
rect 356 115 386 315
<< pmoshvt >>
rect 80 617 110 1217
rect 270 617 300 1217
rect 356 617 386 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 163 315
rect 110 131 121 267
rect 155 131 163 267
rect 110 115 163 131
rect 217 267 270 315
rect 217 131 225 267
rect 259 131 270 267
rect 217 115 270 131
rect 300 267 356 315
rect 300 131 311 267
rect 345 131 356 267
rect 300 115 356 131
rect 386 267 439 315
rect 386 131 397 267
rect 431 131 439 267
rect 386 115 439 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 163 1217
rect 110 657 121 1201
rect 155 657 163 1201
rect 110 617 163 657
rect 217 1201 270 1217
rect 217 657 225 1201
rect 259 657 270 1201
rect 217 617 270 657
rect 300 1201 356 1217
rect 300 657 311 1201
rect 345 657 356 1201
rect 300 617 356 657
rect 386 1201 439 1217
rect 386 657 397 1201
rect 431 657 439 1201
rect 386 617 439 657
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 225 131 259 267
rect 311 131 345 267
rect 397 131 431 267
<< pdiffc >>
rect 35 793 69 1201
rect 121 657 155 1201
rect 225 657 259 1201
rect 311 657 345 1201
rect 397 657 431 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 435 1271 459 1305
rect 493 1271 517 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 459 1271 493 1305
<< poly >>
rect 80 1232 300 1262
rect 80 1217 110 1232
rect 270 1217 300 1232
rect 356 1217 386 1243
rect 80 494 110 617
rect 270 591 300 617
rect 152 555 218 565
rect 152 521 168 555
rect 202 541 218 555
rect 356 541 386 617
rect 202 521 386 541
rect 152 511 386 521
rect 27 478 110 494
rect 27 444 37 478
rect 71 469 110 478
rect 71 444 386 469
rect 27 439 386 444
rect 27 428 110 439
rect 80 315 110 428
rect 152 387 218 397
rect 152 353 168 387
rect 202 373 218 387
rect 202 353 300 373
rect 152 343 300 353
rect 270 315 300 343
rect 356 315 386 439
rect 80 89 110 115
rect 270 89 300 115
rect 356 89 386 115
<< polycont >>
rect 168 521 202 555
rect 37 444 71 478
rect 168 353 202 387
<< locali >>
rect 0 1311 550 1332
rect 0 1271 459 1311
rect 493 1271 550 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 37 478 71 649
rect 37 428 71 444
rect 121 571 155 657
rect 225 1201 259 1217
rect 311 1201 345 1217
rect 225 623 270 657
rect 236 609 270 623
rect 121 555 202 571
rect 121 521 168 555
rect 121 505 202 521
rect 121 403 155 505
rect 121 387 202 403
rect 121 353 168 387
rect 121 337 202 353
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 337
rect 236 301 270 575
rect 311 461 345 657
rect 397 1201 431 1217
rect 397 535 431 657
rect 121 115 155 131
rect 225 267 270 301
rect 311 267 345 279
rect 225 115 259 131
rect 311 115 345 131
rect 397 267 431 501
rect 397 115 431 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 550 61
rect 0 0 550 21
<< viali >>
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 37 649 71 683
rect 236 575 270 609
rect 311 427 345 461
rect 397 501 431 535
rect 311 279 345 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1311 550 1332
rect 0 1277 459 1311
rect 493 1277 550 1311
rect 0 1271 550 1277
rect 25 683 83 689
rect 25 649 37 683
rect 71 649 117 683
rect 25 643 83 649
rect 224 609 282 615
rect 190 575 236 609
rect 270 575 282 609
rect 224 569 282 575
rect 385 535 443 541
rect 351 501 397 535
rect 431 501 443 535
rect 385 495 443 501
rect 299 461 357 467
rect 299 427 311 461
rect 345 427 357 461
rect 299 421 357 427
rect 311 319 345 421
rect 299 313 357 319
rect 299 279 311 313
rect 345 279 357 313
rect 299 273 357 279
rect 0 55 550 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 550 55
rect 0 0 550 21
<< labels >>
rlabel metal1 54 666 54 666 1 S0
port 1 n
rlabel metal1 328 444 328 444 1 Y
port 2 n
rlabel metal1 253 592 253 592 1 A0
port 3 n
rlabel metal1 414 518 414 518 1 A1
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 476 1284 476 1284 1 vdd
<< end >>
