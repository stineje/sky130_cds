* File: sky130_osu_sc_12T_ls__addf_1.pex.spice
* Created: Fri Nov 12 15:33:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%GND 1 2 3 4 5 81 83 91 93 103 105 111
+ 112 125 127 134 146 154 156
c175 103 0 1.20197e-19 $X=2.34 $Y=0.755
c176 81 0 1.04223e-19 $X=-0.045 $Y=0
r177 154 156 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r178 136 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=0.152
+ $X2=6.32 $Y2=0.152
r179 132 150 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.152
r180 132 134 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.74
r181 128 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.152
+ $X2=5.31 $Y2=0.152
r182 127 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.152
+ $X2=6.32 $Y2=0.152
r183 123 149 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.152
r184 123 125 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.755
r185 113 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0.152
+ $X2=3.2 $Y2=0.152
r186 112 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=0.152
+ $X2=5.31 $Y2=0.152
r187 111 146 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.615
+ $X2=3.2 $Y2=0.7
r188 110 148 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.152
r189 110 111 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.615
r190 105 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.152
+ $X2=3.2 $Y2=0.152
r191 101 103 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.34 $Y=0.305
+ $X2=2.34 $Y2=0.755
r192 94 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r193 89 141 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r194 89 91 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r195 83 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r196 81 156 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r197 81 154 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r198 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.34 $Y2=0.305
r199 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.255 $Y2=0.152
r200 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.425 $Y2=0.152
r201 81 136 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.46 $Y=0.152
+ $X2=6.405 $Y2=0.152
r202 81 127 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.235 $Y2=0.152
r203 81 128 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.395 $Y2=0.152
r204 81 112 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=0.152
+ $X2=5.225 $Y2=0.152
r205 81 113 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.285 $Y2=0.152
r206 81 105 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.115 $Y2=0.152
r207 81 106 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.425 $Y2=0.152
r208 81 93 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.255 $Y2=0.152
r209 81 94 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r210 81 83 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r211 5 134 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.195
+ $Y=0.575 $X2=6.32 $Y2=0.74
r212 4 125 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.17
+ $Y=0.575 $X2=5.31 $Y2=0.755
r213 3 146 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.575 $X2=3.2 $Y2=0.7
r214 2 103 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.575 $X2=2.34 $Y2=0.755
r215 1 91 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%VDD 1 2 3 4 5 61 63 70 72 80 82 88 90
+ 100 102 108 114 123 127
r124 123 127 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=6.46 $Y2=4.287
r125 114 127 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=4.25
+ $X2=6.46 $Y2=4.25
r126 112 121 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=4.287
+ $X2=6.32 $Y2=4.287
r127 112 114 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.405 $Y=4.287
+ $X2=6.46 $Y2=4.287
r128 108 111 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.32 $Y=2.955
+ $X2=6.32 $Y2=3.635
r129 106 121 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.32 $Y=4.135
+ $X2=6.32 $Y2=4.287
r130 106 111 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.32 $Y=4.135
+ $X2=6.32 $Y2=3.635
r131 103 120 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=4.287
+ $X2=5.31 $Y2=4.287
r132 103 105 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.395 $Y=4.287
+ $X2=5.78 $Y2=4.287
r133 102 121 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=4.287
+ $X2=6.32 $Y2=4.287
r134 102 105 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=6.235 $Y=4.287
+ $X2=5.78 $Y2=4.287
r135 98 120 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.31 $Y=4.135
+ $X2=5.31 $Y2=4.287
r136 98 100 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.31 $Y=4.135
+ $X2=5.31 $Y2=3.635
r137 95 97 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=4.42 $Y=4.287
+ $X2=5.1 $Y2=4.287
r138 93 95 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.74 $Y=4.287
+ $X2=4.42 $Y2=4.287
r139 91 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=4.287
+ $X2=3.2 $Y2=4.287
r140 91 93 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.285 $Y=4.287
+ $X2=3.74 $Y2=4.287
r141 90 120 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=4.287
+ $X2=5.31 $Y2=4.287
r142 90 97 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.225 $Y=4.287
+ $X2=5.1 $Y2=4.287
r143 86 119 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.2 $Y=4.135
+ $X2=3.2 $Y2=4.287
r144 86 88 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.2 $Y=4.135
+ $X2=3.2 $Y2=3.7
r145 83 118 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=4.287
+ $X2=2.34 $Y2=4.287
r146 83 85 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=2.425 $Y=4.287
+ $X2=3.06 $Y2=4.287
r147 82 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=4.287
+ $X2=3.2 $Y2=4.287
r148 82 85 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.115 $Y=4.287
+ $X2=3.06 $Y2=4.287
r149 78 118 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.34 $Y=4.135
+ $X2=2.34 $Y2=4.287
r150 78 80 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.34 $Y=4.135
+ $X2=2.34 $Y2=3.295
r151 75 77 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r152 73 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r153 73 75 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r154 72 118 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=4.287
+ $X2=2.34 $Y2=4.287
r155 72 77 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=2.255 $Y=4.287
+ $X2=1.7 $Y2=4.287
r156 68 116 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r157 68 70 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.635
r158 65 123 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r159 63 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r160 63 65 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r161 61 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=4.135 $X2=6.46 $Y2=4.22
r162 61 105 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=4.135 $X2=5.78 $Y2=4.22
r163 61 97 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=4.135 $X2=5.1 $Y2=4.22
r164 61 95 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=4.135 $X2=4.42 $Y2=4.22
r165 61 93 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r166 61 85 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r167 61 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r168 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r169 61 75 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r170 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r171 5 111 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=6.195
+ $Y=2.605 $X2=6.32 $Y2=3.635
r172 5 108 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=6.195
+ $Y=2.605 $X2=6.32 $Y2=2.955
r173 4 100 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=2.605 $X2=5.31 $Y2=3.635
r174 3 88 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=2.605 $X2=3.2 $Y2=3.7
r175 2 80 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=2.2
+ $Y=2.605 $X2=2.34 $Y2=3.295
r176 1 70 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%A 3 7 9 11 12 14 15 16 17 18 22 24 25 27
+ 28 30 33 36 41 44 45 47 50 51 53 54 56 60 62 65 70 71 72 73 75 82
c233 73 0 1.55125e-19 $X=2.64 $Y=1.74
c234 72 0 7.77159e-20 $X=5.01 $Y=1.74
c235 65 0 1.50611e-19 $X=2.495 $Y=1.65
c236 54 0 2.67871e-19 $X=5.13 $Y=2.445
c237 47 0 1.89896e-19 $X=2.555 $Y=2.405
c238 45 0 1.29217e-19 $X=2.495 $Y=1.815
c239 36 0 1.32911e-19 $X=5.095 $Y=3.235
c240 28 0 1.58366e-19 $X=2.555 $Y=2.48
c241 24 0 1.79385e-19 $X=2.435 $Y=2.33
c242 22 0 1.57982e-19 $X=2.495 $Y=1.65
c243 16 0 1.75108e-19 $X=2.2 $Y=1.28
r244 73 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.64 $Y=1.74
+ $X2=2.495 $Y2=1.74
r245 72 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.01 $Y=1.74
+ $X2=5.155 $Y2=1.74
r246 72 73 2.28203 $w=1.7e-07 $l=2.37e-06 $layer=MET1_cond $X=5.01 $Y=1.74
+ $X2=2.64 $Y2=1.74
r247 71 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=1.74
+ $X2=0.485 $Y2=1.74
r248 70 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.35 $Y=1.74
+ $X2=2.495 $Y2=1.74
r249 70 71 1.65616 $w=1.7e-07 $l=1.72e-06 $layer=MET1_cond $X=2.35 $Y=1.74
+ $X2=0.63 $Y2=1.74
r250 67 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.495 $Y=1.74
+ $X2=2.495 $Y2=1.74
r251 65 67 4.0073 $w=2.74e-07 $l=9e-08 $layer=LI1_cond $X=2.495 $Y=1.65
+ $X2=2.495 $Y2=1.74
r252 62 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.155 $Y=1.74
+ $X2=5.155 $Y2=1.74
r253 60 69 5.95303 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=1.455
+ $X2=5.155 $Y2=1.37
r254 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.155 $Y=1.455
+ $X2=5.155 $Y2=1.74
r255 56 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=1.74
+ $X2=0.485 $Y2=1.74
r256 53 54 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=5.13 $Y=2.295
+ $X2=5.13 $Y2=2.445
r257 52 53 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.165 $Y=1.535
+ $X2=5.165 $Y2=2.295
r258 50 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.37 $X2=5.155 $Y2=1.37
r259 50 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.37
+ $X2=5.155 $Y2=1.535
r260 50 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.37
+ $X2=5.155 $Y2=1.205
r261 46 47 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.435 $Y=2.405
+ $X2=2.555 $Y2=2.405
r262 41 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.74 $X2=0.485 $Y2=1.74
r263 41 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.74
+ $X2=0.485 $Y2=1.905
r264 41 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.74
+ $X2=0.485 $Y2=1.575
r265 36 54 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.095 $Y=3.235
+ $X2=5.095 $Y2=2.445
r266 33 51 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.095 $Y=0.835
+ $X2=5.095 $Y2=1.205
r267 28 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.555 $Y=2.48
+ $X2=2.555 $Y2=2.405
r268 28 30 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.555 $Y=2.48
+ $X2=2.555 $Y2=3.235
r269 25 44 15.2969 $w=2.1e-07 $l=1.00623e-07 $layer=POLY_cond $X=2.555 $Y=1.205
+ $X2=2.495 $Y2=1.28
r270 25 27 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.555 $Y=1.205
+ $X2=2.555 $Y2=0.835
r271 24 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=2.33
+ $X2=2.435 $Y2=2.405
r272 24 45 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.435 $Y=2.33
+ $X2=2.435 $Y2=1.815
r273 22 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.65 $X2=2.495 $Y2=1.65
r274 20 45 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.495 $Y=1.68
+ $X2=2.495 $Y2=1.815
r275 20 22 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.495 $Y=1.68
+ $X2=2.495 $Y2=1.65
r276 19 44 15.2969 $w=2.1e-07 $l=7.5e-08 $layer=POLY_cond $X=2.495 $Y=1.355
+ $X2=2.495 $Y2=1.28
r277 19 22 65.5412 $w=2.7e-07 $l=2.95e-07 $layer=POLY_cond $X=2.495 $Y=1.355
+ $X2=2.495 $Y2=1.65
r278 17 46 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=2.405
+ $X2=2.435 $Y2=2.405
r279 17 18 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=2.405
+ $X2=2.2 $Y2=2.405
r280 15 44 10.1846 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.36 $Y=1.28
+ $X2=2.495 $Y2=1.28
r281 15 16 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=1.28
+ $X2=2.2 $Y2=1.28
r282 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=2.48
+ $X2=2.2 $Y2=2.405
r283 12 14 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.125 $Y=2.48
+ $X2=2.125 $Y2=3.235
r284 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=1.205
+ $X2=2.2 $Y2=1.28
r285 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.125 $Y=1.205
+ $X2=2.125 $Y2=0.835
r286 7 43 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=1.905
r287 3 42 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%B 3 7 11 15 19 23 27 31 34 40 43 47 52
+ 56 58 60 63 70 72 78 80 81 83 85 86 87 88 97
c272 88 0 3.48262e-19 $X=3.12 $Y=2.48
c273 81 0 1.8823e-19 $X=0.63 $Y=2.48
c274 72 0 1.96262e-19 $X=0.485 $Y=2.28
c275 70 0 1.89283e-19 $X=4.265 $Y=2.48
c276 58 0 1.04223e-19 $X=2.1 $Y=2.48
c277 47 0 7.77159e-20 $X=4.265 $Y=2.135
c278 43 0 1.79385e-19 $X=2.975 $Y=1.655
c279 40 0 1.37671e-19 $X=2.015 $Y=1.95
c280 23 0 1.29405e-20 $X=2.985 $Y=3.235
r281 88 95 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.12 $Y=2.48
+ $X2=2.975 $Y2=2.48
r282 87 97 0.101907 $w=2.4e-07 $l=1.45e-07 $layer=MET1_cond $X=4.12 $Y=2.48
+ $X2=4.265 $Y2=2.48
r283 87 88 0.962882 $w=1.7e-07 $l=1e-06 $layer=MET1_cond $X=4.12 $Y=2.48
+ $X2=3.12 $Y2=2.48
r284 86 93 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.45 $Y=2.48
+ $X2=2.305 $Y2=2.48
r285 85 95 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.83 $Y=2.48
+ $X2=2.975 $Y2=2.48
r286 85 86 0.365895 $w=1.7e-07 $l=3.8e-07 $layer=MET1_cond $X=2.83 $Y=2.48
+ $X2=2.45 $Y2=2.48
r287 81 90 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=2.48
+ $X2=0.485 $Y2=2.48
r288 81 83 0.0144432 $w=1.7e-07 $l=1.5e-08 $layer=MET1_cond $X=0.63 $Y=2.48
+ $X2=0.645 $Y2=2.48
r289 80 93 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.16 $Y=2.48
+ $X2=2.305 $Y2=2.48
r290 80 83 1.45877 $w=1.7e-07 $l=1.515e-06 $layer=MET1_cond $X=2.16 $Y=2.48
+ $X2=0.645 $Y2=2.48
r291 75 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=2.48
+ $X2=0.485 $Y2=2.48
r292 72 75 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.485 $Y=2.28
+ $X2=0.485 $Y2=2.48
r293 70 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.265 $Y=2.48
+ $X2=4.265 $Y2=2.48
r294 68 78 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=2.22
+ $X2=4.265 $Y2=2.135
r295 68 70 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.265 $Y=2.22
+ $X2=4.265 $Y2=2.48
r296 66 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=2.48
+ $X2=2.975 $Y2=2.48
r297 63 66 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.975 $Y=1.655
+ $X2=2.975 $Y2=2.48
r298 60 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.305 $Y=2.48
+ $X2=2.305 $Y2=2.48
r299 58 60 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.1 $Y=2.48
+ $X2=2.305 $Y2=2.48
r300 54 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.015 $Y=2.395
+ $X2=2.1 $Y2=2.48
r301 54 56 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.015 $Y=2.395
+ $X2=2.015 $Y2=1.95
r302 50 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=2.28
+ $X2=0.485 $Y2=2.28
r303 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.57 $Y=2.28
+ $X2=0.895 $Y2=2.28
r304 47 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=2.135 $X2=4.265 $Y2=2.135
r305 47 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.135
+ $X2=4.265 $Y2=2.3
r306 47 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.135
+ $X2=4.265 $Y2=1.97
r307 43 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.655 $X2=2.975 $Y2=1.655
r308 43 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.655
+ $X2=2.975 $Y2=1.82
r309 43 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.655
+ $X2=2.975 $Y2=1.49
r310 40 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=1.95 $X2=2.015 $Y2=1.95
r311 37 40 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.765 $Y=1.95
+ $X2=2.015 $Y2=1.95
r312 34 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=2.28 $X2=0.895 $Y2=2.28
r313 34 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.28
+ $X2=0.895 $Y2=2.445
r314 34 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.28
+ $X2=0.895 $Y2=2.115
r315 31 49 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=4.275 $Y=3.235
+ $X2=4.275 $Y2=2.3
r316 27 48 581.989 $w=1.5e-07 $l=1.135e-06 $layer=POLY_cond $X=4.275 $Y=0.835
+ $X2=4.275 $Y2=1.97
r317 23 45 725.564 $w=1.5e-07 $l=1.415e-06 $layer=POLY_cond $X=2.985 $Y=3.235
+ $X2=2.985 $Y2=1.82
r318 19 44 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.985 $Y=0.835
+ $X2=2.985 $Y2=1.49
r319 13 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.115
+ $X2=1.765 $Y2=1.95
r320 13 15 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.765 $Y=2.115
+ $X2=1.765 $Y2=3.235
r321 9 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.785
+ $X2=1.765 $Y2=1.95
r322 9 11 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.765 $Y=1.785
+ $X2=1.765 $Y2=0.835
r323 7 36 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.445
r324 3 35 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=0.905 $Y=0.835
+ $X2=0.905 $Y2=2.115
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%CI 3 7 11 15 19 23 26 30 32 36 42 47 52
+ 53 54 55 57 64
c180 64 0 1.89283e-19 $X=4.745 $Y=2.11
c181 54 0 1.70419e-20 $X=4.6 $Y=2.11
c182 53 0 1.14581e-19 $X=1.48 $Y=2.11
c183 52 0 1.29217e-19 $X=3.25 $Y=2.11
c184 11 0 1.41673e-19 $X=3.415 $Y=0.835
c185 7 0 1.63624e-19 $X=1.335 $Y=3.235
r186 55 62 0.119415 $w=2.3e-07 $l=1.7e-07 $layer=MET1_cond $X=3.585 $Y=2.11
+ $X2=3.415 $Y2=2.11
r187 54 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.6 $Y=2.11
+ $X2=4.745 $Y2=2.11
r188 54 55 0.977326 $w=1.7e-07 $l=1.015e-06 $layer=MET1_cond $X=4.6 $Y=2.11
+ $X2=3.585 $Y2=2.11
r189 53 57 0.109791 $w=2.3e-07 $l=1.55e-07 $layer=MET1_cond $X=1.48 $Y=2.11
+ $X2=1.325 $Y2=2.11
r190 52 62 0.116207 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=3.25 $Y=2.11
+ $X2=3.415 $Y2=2.11
r191 52 53 1.7043 $w=1.7e-07 $l=1.77e-06 $layer=MET1_cond $X=3.25 $Y=2.11
+ $X2=1.48 $Y2=2.11
r192 50 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.745 $Y=2.11
+ $X2=4.745 $Y2=2.11
r193 47 50 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.745 $Y=1.92
+ $X2=4.745 $Y2=2.11
r194 42 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.415 $Y=2.11
+ $X2=3.415 $Y2=2.11
r195 39 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.325 $Y=2.11
+ $X2=1.325 $Y2=2.11
r196 36 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.325 $Y=1.74
+ $X2=1.325 $Y2=2.11
r197 32 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=1.92 $X2=4.745 $Y2=1.92
r198 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.92
+ $X2=4.745 $Y2=2.085
r199 32 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.92
+ $X2=4.745 $Y2=1.755
r200 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=2.11 $X2=3.415 $Y2=2.11
r201 26 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.74 $X2=1.325 $Y2=1.74
r202 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.74
+ $X2=1.325 $Y2=1.905
r203 26 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.74
+ $X2=1.325 $Y2=1.575
r204 23 34 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=4.685 $Y=3.235
+ $X2=4.685 $Y2=2.085
r205 19 33 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=4.685 $Y=0.835
+ $X2=4.685 $Y2=1.755
r206 13 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.275
+ $X2=3.415 $Y2=2.11
r207 13 15 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.415 $Y=2.275
+ $X2=3.415 $Y2=3.235
r208 9 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.945
+ $X2=3.415 $Y2=2.11
r209 9 11 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=3.415 $Y=1.945
+ $X2=3.415 $Y2=0.835
r210 7 28 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.335 $Y=3.235
+ $X2=1.335 $Y2=1.905
r211 3 27 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.335 $Y=0.835
+ $X2=1.335 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%CON 1 3 11 15 19 23 26 28 33 37 42 45 49
+ 53 56 62 64 65 66 67 74
c172 67 0 2.91173e-19 $X=4.1 $Y=1.37
c173 65 0 3.3309e-19 $X=1.81 $Y=1.37
c174 64 0 1.85295e-19 $X=3.855 $Y=1.37
c175 53 0 8.19432e-20 $X=1.665 $Y=2.637
c176 42 0 1.55125e-19 $X=1.665 $Y=1.37
c177 33 0 1.20197e-19 $X=1.55 $Y=0.755
c178 28 0 1.71092e-19 $X=6.41 $Y=2.26
c179 26 0 1.29042e-19 $X=3.845 $Y=1.455
c180 11 0 1.00659e-19 $X=3.845 $Y=0.835
r181 67 72 0.0937512 $w=2.3e-07 $l=1.3e-07 $layer=MET1_cond $X=4.1 $Y=1.37
+ $X2=3.97 $Y2=1.37
r182 66 74 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.995 $Y=1.37
+ $X2=6.14 $Y2=1.37
r183 66 67 1.82466 $w=1.7e-07 $l=1.895e-06 $layer=MET1_cond $X=5.995 $Y=1.37
+ $X2=4.1 $Y2=1.37
r184 65 69 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.81 $Y=1.37
+ $X2=1.665 $Y2=1.37
r185 64 72 0.0841272 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=3.855 $Y=1.37
+ $X2=3.97 $Y2=1.37
r186 64 65 1.96909 $w=1.7e-07 $l=2.045e-06 $layer=MET1_cond $X=3.855 $Y=1.37
+ $X2=1.81 $Y2=1.37
r187 60 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.14 $Y=1.37
+ $X2=6.14 $Y2=1.37
r188 60 62 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.14 $Y=1.37
+ $X2=6.41 $Y2=1.37
r189 58 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.97 $Y=1.37
+ $X2=3.97 $Y2=1.37
r190 56 58 7.36715 $w=2.07e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.412
+ $X2=3.97 $Y2=1.412
r191 51 53 6.89435 $w=1.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=2.637
+ $X2=1.665 $Y2=2.637
r192 47 49 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=1.2
+ $X2=1.665 $Y2=1.2
r193 43 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.455
+ $X2=6.41 $Y2=1.37
r194 43 45 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=6.41 $Y=1.455
+ $X2=6.41 $Y2=2.26
r195 42 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.665 $Y=1.37
+ $X2=1.665 $Y2=1.37
r196 40 53 1.22693 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=1.665 $Y=2.545
+ $X2=1.665 $Y2=2.637
r197 40 42 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.665 $Y=2.545
+ $X2=1.665 $Y2=1.37
r198 39 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.285
+ $X2=1.665 $Y2=1.2
r199 39 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.285
+ $X2=1.665 $Y2=1.37
r200 35 51 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.55 $Y=2.73
+ $X2=1.55 $Y2=2.637
r201 35 37 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.55 $Y=2.73
+ $X2=1.55 $Y2=3.295
r202 31 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.2
r203 31 33 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=0.755
r204 28 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=2.26 $X2=6.41 $Y2=2.26
r205 28 30 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.26
+ $X2=6.442 $Y2=2.425
r206 28 29 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.26
+ $X2=6.442 $Y2=2.095
r207 26 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.455 $X2=3.845 $Y2=1.455
r208 23 30 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.535 $Y=3.235
+ $X2=6.535 $Y2=2.425
r209 19 29 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=6.535 $Y=0.835
+ $X2=6.535 $Y2=2.095
r210 13 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.62
+ $X2=3.845 $Y2=1.455
r211 13 15 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=3.845 $Y=1.62
+ $X2=3.845 $Y2=3.235
r212 9 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.29
+ $X2=3.845 $Y2=1.455
r213 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.845 $Y=1.29
+ $X2=3.845 $Y2=0.835
r214 3 37 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.295
r215 1 33 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%A_784_115# 1 3 11 15 18 20 21 22 23 25
+ 27 30 32 35 37
c129 35 0 1.26797e-19 $X=4.06 $Y=0.74
c130 32 0 9.63581e-20 $X=5.415 $Y=2.77
c131 23 0 1.70419e-20 $X=4.06 $Y=2.94
c132 22 0 3.34795e-19 $X=3.93 $Y=1.795
c133 18 0 3.07391e-19 $X=5.585 $Y=2.275
c134 15 0 1.71513e-19 $X=5.585 $Y=3.235
c135 11 0 1.71092e-19 $X=5.585 $Y=0.835
r136 37 39 7.30282 $w=2.84e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=2.275
+ $X2=5.585 $Y2=2.275
r137 35 36 11.9608 $w=2.55e-07 $l=2.5e-07 $layer=LI1_cond $X=4.06 $Y=0.78
+ $X2=4.31 $Y2=0.78
r138 31 37 3.73949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=2.44
+ $X2=5.415 $Y2=2.275
r139 31 32 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.415 $Y=2.44
+ $X2=5.415 $Y2=2.77
r140 29 36 3.11056 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.31 $Y=0.95
+ $X2=4.31 $Y2=0.78
r141 29 30 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.31 $Y=0.95
+ $X2=4.31 $Y2=1.71
r142 28 33 3.40055 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=4.145 $Y=2.855
+ $X2=3.935 $Y2=2.855
r143 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.33 $Y=2.855
+ $X2=5.415 $Y2=2.77
r144 27 28 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=5.33 $Y=2.855
+ $X2=4.145 $Y2=2.855
r145 23 33 5.49396 $w=2.68e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.06 $Y=2.94
+ $X2=3.935 $Y2=2.855
r146 23 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.06 $Y=2.94
+ $X2=4.06 $Y2=3.295
r147 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.225 $Y=1.795
+ $X2=4.31 $Y2=1.71
r148 21 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.225 $Y=1.795
+ $X2=3.93 $Y2=1.795
r149 20 33 15.5089 $w=2.68e-07 $l=3.47095e-07 $layer=LI1_cond $X=3.845 $Y=2.55
+ $X2=3.935 $Y2=2.855
r150 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=1.88
+ $X2=3.93 $Y2=1.795
r151 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.845 $Y=1.88
+ $X2=3.845 $Y2=2.55
r152 18 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.585
+ $Y=2.275 $X2=5.585 $Y2=2.275
r153 13 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.44
+ $X2=5.585 $Y2=2.275
r154 13 15 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=5.585 $Y=2.44
+ $X2=5.585 $Y2=3.235
r155 9 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.11
+ $X2=5.585 $Y2=2.275
r156 9 11 653.777 $w=1.5e-07 $l=1.275e-06 $layer=POLY_cond $X=5.585 $Y=2.11
+ $X2=5.585 $Y2=0.835
r157 3 25 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=3.92
+ $Y=2.605 $X2=4.06 $Y2=3.295
r158 1 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.575 $X2=4.06 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%A_27_521# 1 2 11 13 17
c15 14 0 1.8823e-19 $X=0.345 $Y=2.98
r16 15 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.12 $Y=3.065
+ $X2=1.12 $Y2=3.295
r17 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=2.98
+ $X2=1.12 $Y2=3.065
r18 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=2.98
+ $X2=0.345 $Y2=2.98
r19 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.065
+ $X2=0.345 $Y2=2.98
r20 9 11 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.26 $Y=3.065
+ $X2=0.26 $Y2=3.295
r21 2 17 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.295
r22 1 11 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%A_526_521# 1 2 11 15 18
r15 13 15 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.63 $Y=3.315
+ $X2=3.63 $Y2=3.55
r16 12 18 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.855 $Y=3.23
+ $X2=2.77 $Y2=3.19
r17 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=3.23
+ $X2=3.63 $Y2=3.315
r18 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=3.23
+ $X2=2.855 $Y2=3.23
r19 2 15 600 $w=1.7e-07 $l=1.01258e-06 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=2.605 $X2=3.63 $Y2=3.55
r20 1 18 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=2.605 $X2=2.77 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%S 1 3 11 17 20 23 27 30
c51 30 0 1.32911e-19 $X=5.8 $Y=2.855
c52 27 0 1.41304e-19 $X=5.925 $Y=2.77
c53 23 0 1.66087e-19 $X=5.925 $Y=1.74
r54 25 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=2.77
+ $X2=5.925 $Y2=2.77
r55 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=1.74
+ $X2=5.925 $Y2=1.74
r56 20 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=2.685
+ $X2=5.925 $Y2=2.77
r57 19 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=1.825
+ $X2=5.925 $Y2=1.74
r58 19 20 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.925 $Y=1.825
+ $X2=5.925 $Y2=2.685
r59 15 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.8 $Y=2.855 $X2=5.8
+ $Y2=2.855
r60 15 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.855 $X2=5.8
+ $Y2=2.77
r61 15 17 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.8 $Y=2.855 $X2=5.8
+ $Y2=3.295
r62 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=1.655 $X2=5.8
+ $Y2=1.74
r63 9 11 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.8 $Y=1.655 $X2=5.8
+ $Y2=0.755
r64 3 17 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=5.66
+ $Y=2.605 $X2=5.8 $Y2=3.295
r65 1 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.66 $Y=0.575
+ $X2=5.8 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%CO 1 3 10 20
r16 15 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.75 $Y=2.955
+ $X2=6.75 $Y2=3.635
r17 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.75 $Y=2.48
+ $X2=6.75 $Y2=2.48
r18 13 15 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.75 $Y=2.48
+ $X2=6.75 $Y2=2.955
r19 10 13 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=6.75 $Y=0.755
+ $X2=6.75 $Y2=2.48
r20 3 17 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=2.605 $X2=6.75 $Y2=3.635
r21 3 15 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=2.605 $X2=6.75 $Y2=2.955
r22 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.61 $Y=0.575
+ $X2=6.75 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%A_27_115# 1 2 11 13 17 19
r27 19 20 13.626 $w=1.73e-07 $l=2.15e-07 $layer=LI1_cond $X=0.262 $Y=1.16
+ $X2=0.262 $Y2=0.945
r28 15 17 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.12 $Y=1.075
+ $X2=1.12 $Y2=0.755
r29 14 19 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.35 $Y=1.16
+ $X2=0.262 $Y2=1.16
r30 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=1.12 $Y2=1.075
r31 13 14 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.35 $Y2=1.16
r32 11 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.755
+ $X2=0.26 $Y2=0.945
r33 2 17 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
r34 1 11 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__ADDF_1%A_526_115# 1 2 11 13 14 17
c29 13 0 1.02903e-19 $X=3.545 $Y=1.115
r30 15 17 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.63 $Y=1.03
+ $X2=3.63 $Y2=0.755
r31 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=1.115
+ $X2=3.63 $Y2=1.03
r32 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=1.115
+ $X2=2.855 $Y2=1.115
r33 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.03
+ $X2=2.855 $Y2=1.115
r34 9 11 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.77 $Y=1.03
+ $X2=2.77 $Y2=0.755
r35 2 17 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.49 $Y=0.575
+ $X2=3.63 $Y2=0.755
r36 1 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.63 $Y=0.575
+ $X2=2.77 $Y2=0.755
.ends

