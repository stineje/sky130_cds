* File: sky130_osu_sc_15T_ms__tbufi_1.pxi.spice
* Created: Fri Nov 12 14:46:34 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__TBUFI_1%GND N_GND_M1003_d N_GND_M1003_b N_GND_c_3_p
+ N_GND_c_4_p GND N_GND_c_5_p PM_SKY130_OSU_SC_15T_MS__TBUFI_1%GND
x_PM_SKY130_OSU_SC_15T_MS__TBUFI_1%VDD N_VDD_M1004_d N_VDD_M1004_b N_VDD_c_40_p
+ N_VDD_c_41_p N_VDD_c_48_p VDD N_VDD_c_42_p
+ PM_SKY130_OSU_SC_15T_MS__TBUFI_1%VDD
x_PM_SKY130_OSU_SC_15T_MS__TBUFI_1%OE N_OE_c_60_n N_OE_c_61_n N_OE_M1003_g
+ N_OE_c_76_n N_OE_M1004_g N_OE_c_65_n N_OE_M1000_g N_OE_c_68_n N_OE_c_69_n
+ N_OE_c_71_n N_OE_c_73_n OE PM_SKY130_OSU_SC_15T_MS__TBUFI_1%OE
x_PM_SKY130_OSU_SC_15T_MS__TBUFI_1%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1004_s N_A_27_115#_M1002_g N_A_27_115#_c_126_n
+ N_A_27_115#_c_127_n N_A_27_115#_c_130_n N_A_27_115#_c_131_n
+ N_A_27_115#_c_132_n N_A_27_115#_c_133_n
+ PM_SKY130_OSU_SC_15T_MS__TBUFI_1%A_27_115#
x_PM_SKY130_OSU_SC_15T_MS__TBUFI_1%A N_A_M1005_g N_A_M1001_g N_A_c_178_n
+ N_A_c_179_n N_A_c_180_n A PM_SKY130_OSU_SC_15T_MS__TBUFI_1%A
x_PM_SKY130_OSU_SC_15T_MS__TBUFI_1%Y N_Y_M1005_d N_Y_M1001_d N_Y_c_224_n
+ N_Y_c_226_n Y N_Y_c_228_n N_Y_c_230_n PM_SKY130_OSU_SC_15T_MS__TBUFI_1%Y
cc_1 N_GND_M1003_b N_OE_c_60_n 0.0680245f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.6
cc_2 N_GND_M1003_b N_OE_c_61_n 0.0183291f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.39
cc_3 N_GND_c_3_p N_OE_c_61_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.39
cc_4 N_GND_c_4_p N_OE_c_61_n 0.00388248f $X=0.69 $Y=0.865 $X2=0.475 $Y2=1.39
cc_5 N_GND_c_5_p N_OE_c_61_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.39
cc_6 N_GND_M1003_b N_OE_c_65_n 0.0200336f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.39
cc_7 N_GND_c_4_p N_OE_c_65_n 0.00388248f $X=0.69 $Y=0.865 $X2=0.905 $Y2=1.39
cc_8 N_GND_c_5_p N_OE_c_65_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=1.39
cc_9 N_GND_M1003_b N_OE_c_68_n 0.00923524f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.675
cc_10 N_GND_M1003_b N_OE_c_69_n 0.0546824f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.59
cc_11 N_GND_c_4_p N_OE_c_69_n 0.00244833f $X=0.69 $Y=0.865 $X2=0.69 $Y2=1.59
cc_12 N_GND_M1003_b N_OE_c_71_n 0.00260472f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.59
cc_13 N_GND_c_4_p N_OE_c_71_n 0.00508043f $X=0.69 $Y=0.865 $X2=0.69 $Y2=1.59
cc_14 N_GND_M1003_b N_OE_c_73_n 7.18349e-19 $X=-0.045 $Y=0 $X2=0.69 $Y2=1.59
cc_15 N_GND_c_4_p N_OE_c_73_n 0.0046483f $X=0.69 $Y=0.865 $X2=0.69 $Y2=1.59
cc_16 N_GND_M1003_b OE 0.0107998f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.7
cc_17 N_GND_M1003_b N_A_27_115#_M1002_g 0.014739f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=3.825
cc_18 N_GND_M1003_b N_A_27_115#_c_126_n 0.0326306f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=2.22
cc_19 N_GND_M1003_b N_A_27_115#_c_127_n 0.0303682f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_20 N_GND_c_3_p N_A_27_115#_c_127_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_21 N_GND_c_5_p N_A_27_115#_c_127_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_22 N_GND_M1003_b N_A_27_115#_c_130_n 0.0116459f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.205
cc_23 N_GND_M1003_b N_A_27_115#_c_131_n 0.0101855f $X=-0.045 $Y=0 $X2=0.715
+ $Y2=2.22
cc_24 N_GND_M1003_b N_A_27_115#_c_132_n 0.00665288f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.22
cc_25 N_GND_M1003_b N_A_27_115#_c_133_n 0.00288071f $X=-0.045 $Y=0 $X2=0.8
+ $Y2=2.22
cc_26 N_GND_M1003_b N_A_M1005_g 0.0437489f $X=-0.045 $Y=0 $X2=1.265 $Y2=0.945
cc_27 N_GND_c_5_p N_A_M1005_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.265 $Y2=0.945
cc_28 N_GND_M1003_b N_A_M1001_g 0.0372976f $X=-0.045 $Y=0 $X2=1.265 $Y2=3.825
cc_29 N_GND_M1003_b N_A_c_178_n 0.0369358f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.83
cc_30 N_GND_M1003_b N_A_c_179_n 0.00459479f $X=-0.045 $Y=0 $X2=1.14 $Y2=3.07
cc_31 N_GND_M1003_b N_A_c_180_n 0.00983127f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.83
cc_32 N_GND_M1003_b N_Y_c_224_n 0.00913846f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.865
cc_33 N_GND_c_5_p N_Y_c_224_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.48 $Y2=0.865
cc_34 N_GND_M1003_b N_Y_c_226_n 0.0151339f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.33
cc_35 N_GND_M1003_b Y 0.0383474f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.56
cc_36 N_GND_M1003_b N_Y_c_228_n 0.0122638f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.22
cc_37 N_GND_c_4_p N_Y_c_228_n 9.45275e-19 $X=0.69 $Y=0.865 $X2=1.48 $Y2=1.22
cc_38 N_GND_M1003_b N_Y_c_230_n 0.0157299f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.33
cc_39 N_VDD_M1004_b N_OE_c_76_n 0.0187209f $X=-0.045 $Y=2.645 $X2=0.475 $Y2=2.75
cc_40 N_VDD_c_40_p N_OE_c_76_n 0.00496961f $X=0.605 $Y=5.397 $X2=0.475 $Y2=2.75
cc_41 N_VDD_c_41_p N_OE_c_76_n 0.00362996f $X=0.69 $Y=3.545 $X2=0.475 $Y2=2.75
cc_42 N_VDD_c_42_p N_OE_c_76_n 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=2.75
cc_43 N_VDD_M1004_b N_OE_c_68_n 0.0152497f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=2.675
cc_44 N_VDD_M1004_b OE 0.00599741f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.7
cc_45 N_VDD_c_41_p OE 0.00759884f $X=0.69 $Y=3.545 $X2=0.69 $Y2=2.7
cc_46 N_VDD_M1004_b N_A_27_115#_M1002_g 0.0192164f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_47 N_VDD_c_41_p N_A_27_115#_M1002_g 0.00362996f $X=0.69 $Y=3.545 $X2=0.905
+ $Y2=3.825
cc_48 N_VDD_c_48_p N_A_27_115#_M1002_g 0.00496961f $X=1.02 $Y=5.33 $X2=0.905
+ $Y2=3.825
cc_49 N_VDD_c_42_p N_A_27_115#_M1002_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.905
+ $Y2=3.825
cc_50 N_VDD_M1004_b N_A_27_115#_c_130_n 0.00845875f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.205
cc_51 N_VDD_c_40_p N_A_27_115#_c_130_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.205
cc_52 N_VDD_c_42_p N_A_27_115#_c_130_n 0.00435496f $X=1.02 $Y=5.36 $X2=0.26
+ $Y2=3.205
cc_53 N_VDD_M1004_b N_A_M1001_g 0.0230844f $X=-0.045 $Y=2.645 $X2=1.265
+ $Y2=3.825
cc_54 N_VDD_c_48_p N_A_M1001_g 0.00496961f $X=1.02 $Y=5.33 $X2=1.265 $Y2=3.825
cc_55 N_VDD_c_42_p N_A_M1001_g 0.00429146f $X=1.02 $Y=5.36 $X2=1.265 $Y2=3.825
cc_56 N_VDD_M1004_b N_A_c_179_n 5.73277e-19 $X=-0.045 $Y=2.645 $X2=1.14 $Y2=3.07
cc_57 N_VDD_M1004_b N_Y_c_226_n 0.0102055f $X=-0.045 $Y=2.645 $X2=1.48 $Y2=2.33
cc_58 N_VDD_c_48_p N_Y_c_226_n 0.00477009f $X=1.02 $Y=5.33 $X2=1.48 $Y2=2.33
cc_59 N_VDD_c_42_p N_Y_c_226_n 0.00435496f $X=1.02 $Y=5.36 $X2=1.48 $Y2=2.33
cc_60 N_OE_c_60_n N_A_27_115#_M1002_g 0.00266681f $X=0.27 $Y=2.6 $X2=0.905
+ $Y2=3.825
cc_61 N_OE_c_68_n N_A_27_115#_M1002_g 0.0402653f $X=0.475 $Y=2.675 $X2=0.905
+ $Y2=3.825
cc_62 OE N_A_27_115#_M1002_g 0.0135769f $X=0.69 $Y=2.7 $X2=0.905 $Y2=3.825
cc_63 N_OE_c_60_n N_A_27_115#_c_126_n 0.0126749f $X=0.27 $Y=2.6 $X2=0.905
+ $Y2=2.22
cc_64 N_OE_c_69_n N_A_27_115#_c_126_n 0.0119465f $X=0.69 $Y=1.59 $X2=0.905
+ $Y2=2.22
cc_65 N_OE_c_71_n N_A_27_115#_c_126_n 4.88301e-19 $X=0.69 $Y=1.59 $X2=0.905
+ $Y2=2.22
cc_66 OE N_A_27_115#_c_126_n 0.00242154f $X=0.69 $Y=2.7 $X2=0.905 $Y2=2.22
cc_67 N_OE_c_60_n N_A_27_115#_c_127_n 0.0232517f $X=0.27 $Y=2.6 $X2=0.26
+ $Y2=0.865
cc_68 N_OE_c_61_n N_A_27_115#_c_127_n 0.00957633f $X=0.475 $Y=1.39 $X2=0.26
+ $Y2=0.865
cc_69 N_OE_c_69_n N_A_27_115#_c_127_n 0.0135784f $X=0.69 $Y=1.59 $X2=0.26
+ $Y2=0.865
cc_70 N_OE_c_71_n N_A_27_115#_c_127_n 0.0116068f $X=0.69 $Y=1.59 $X2=0.26
+ $Y2=0.865
cc_71 N_OE_c_73_n N_A_27_115#_c_127_n 0.00367353f $X=0.69 $Y=1.59 $X2=0.26
+ $Y2=0.865
cc_72 OE N_A_27_115#_c_127_n 0.015341f $X=0.69 $Y=2.7 $X2=0.26 $Y2=0.865
cc_73 N_OE_c_60_n N_A_27_115#_c_130_n 0.0103172f $X=0.27 $Y=2.6 $X2=0.26
+ $Y2=3.205
cc_74 N_OE_c_76_n N_A_27_115#_c_130_n 0.00766083f $X=0.475 $Y=2.75 $X2=0.26
+ $Y2=3.205
cc_75 N_OE_c_68_n N_A_27_115#_c_130_n 0.00887831f $X=0.475 $Y=2.675 $X2=0.26
+ $Y2=3.205
cc_76 OE N_A_27_115#_c_130_n 0.0193905f $X=0.69 $Y=2.7 $X2=0.26 $Y2=3.205
cc_77 N_OE_c_68_n N_A_27_115#_c_131_n 0.00703932f $X=0.475 $Y=2.675 $X2=0.715
+ $Y2=2.22
cc_78 N_OE_c_69_n N_A_27_115#_c_131_n 0.00292172f $X=0.69 $Y=1.59 $X2=0.715
+ $Y2=2.22
cc_79 N_OE_c_71_n N_A_27_115#_c_131_n 0.00456286f $X=0.69 $Y=1.59 $X2=0.715
+ $Y2=2.22
cc_80 N_OE_c_73_n N_A_27_115#_c_131_n 0.00123496f $X=0.69 $Y=1.59 $X2=0.715
+ $Y2=2.22
cc_81 OE N_A_27_115#_c_131_n 0.0142208f $X=0.69 $Y=2.7 $X2=0.715 $Y2=2.22
cc_82 N_OE_c_60_n N_A_27_115#_c_132_n 0.00700951f $X=0.27 $Y=2.6 $X2=0.26
+ $Y2=2.22
cc_83 N_OE_c_60_n N_A_27_115#_c_133_n 7.28524e-19 $X=0.27 $Y=2.6 $X2=0.8
+ $Y2=2.22
cc_84 N_OE_c_69_n N_A_27_115#_c_133_n 7.06691e-19 $X=0.69 $Y=1.59 $X2=0.8
+ $Y2=2.22
cc_85 N_OE_c_71_n N_A_27_115#_c_133_n 0.00377605f $X=0.69 $Y=1.59 $X2=0.8
+ $Y2=2.22
cc_86 N_OE_c_73_n N_A_27_115#_c_133_n 0.00129814f $X=0.69 $Y=1.59 $X2=0.8
+ $Y2=2.22
cc_87 OE N_A_27_115#_c_133_n 0.0157069f $X=0.69 $Y=2.7 $X2=0.8 $Y2=2.22
cc_88 N_OE_c_65_n N_A_M1005_g 0.0674578f $X=0.905 $Y=1.39 $X2=1.265 $Y2=0.945
cc_89 N_OE_c_69_n N_A_M1005_g 0.00693622f $X=0.69 $Y=1.59 $X2=1.265 $Y2=0.945
cc_90 N_OE_c_71_n N_A_M1005_g 0.00287993f $X=0.69 $Y=1.59 $X2=1.265 $Y2=0.945
cc_91 OE N_A_c_178_n 2.30744e-19 $X=0.69 $Y=2.7 $X2=1.325 $Y2=1.83
cc_92 OE N_A_c_179_n 0.0257797f $X=0.69 $Y=2.7 $X2=1.14 $Y2=3.07
cc_93 N_OE_c_69_n N_A_c_180_n 2.20759e-19 $X=0.69 $Y=1.59 $X2=1.325 $Y2=1.83
cc_94 OE N_A_c_180_n 0.00765298f $X=0.69 $Y=2.7 $X2=1.325 $Y2=1.83
cc_95 N_OE_c_76_n A 8.46663e-19 $X=0.475 $Y=2.75 $X2=1.14 $Y2=3.07
cc_96 OE A 0.004991f $X=0.69 $Y=2.7 $X2=1.14 $Y2=3.07
cc_97 N_OE_c_69_n Y 2.15427e-19 $X=0.69 $Y=1.59 $X2=1.525 $Y2=1.56
cc_98 N_OE_c_71_n Y 0.00375884f $X=0.69 $Y=1.59 $X2=1.525 $Y2=1.56
cc_99 N_OE_c_73_n Y 0.0105247f $X=0.69 $Y=1.59 $X2=1.525 $Y2=1.56
cc_100 N_OE_c_65_n N_Y_c_228_n 0.00101819f $X=0.905 $Y=1.39 $X2=1.48 $Y2=1.22
cc_101 OE N_Y_c_230_n 0.0100845f $X=0.69 $Y=2.7 $X2=1.48 $Y2=2.33
cc_102 N_A_27_115#_c_126_n N_A_M1001_g 0.172375f $X=0.905 $Y=2.22 $X2=1.265
+ $Y2=3.825
cc_103 N_A_27_115#_c_133_n N_A_M1001_g 2.80054e-19 $X=0.8 $Y=2.22 $X2=1.265
+ $Y2=3.825
cc_104 N_A_27_115#_c_126_n N_A_c_179_n 0.0186036f $X=0.905 $Y=2.22 $X2=1.14
+ $Y2=3.07
cc_105 N_A_27_115#_c_133_n N_A_c_179_n 0.0209392f $X=0.8 $Y=2.22 $X2=1.14
+ $Y2=3.07
cc_106 N_A_27_115#_M1002_g A 0.01062f $X=0.905 $Y=3.825 $X2=1.14 $Y2=3.07
cc_107 N_A_27_115#_c_130_n A 0.00539687f $X=0.26 $Y=3.205 $X2=1.14 $Y2=3.07
cc_108 N_A_c_179_n A_196_565# 0.00616226f $X=1.14 $Y=3.07 $X2=0.98 $Y2=2.825
cc_109 A A_196_565# 0.0123769f $X=1.14 $Y=3.07 $X2=0.98 $Y2=2.825
cc_110 N_A_M1005_g N_Y_c_224_n 0.00740756f $X=1.265 $Y=0.945 $X2=1.48 $Y2=0.865
cc_111 N_A_c_178_n N_Y_c_224_n 8.70049e-19 $X=1.325 $Y=1.83 $X2=1.48 $Y2=0.865
cc_112 N_A_c_180_n N_Y_c_224_n 0.00216439f $X=1.325 $Y=1.83 $X2=1.48 $Y2=0.865
cc_113 N_A_M1001_g N_Y_c_226_n 0.0168888f $X=1.265 $Y=3.825 $X2=1.48 $Y2=2.33
cc_114 N_A_c_178_n N_Y_c_226_n 0.00102058f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
cc_115 N_A_c_179_n N_Y_c_226_n 0.049778f $X=1.14 $Y=3.07 $X2=1.48 $Y2=2.33
cc_116 N_A_c_180_n N_Y_c_226_n 0.00330615f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
cc_117 A N_Y_c_226_n 0.00706656f $X=1.14 $Y=3.07 $X2=1.48 $Y2=2.33
cc_118 N_A_M1005_g Y 0.00631192f $X=1.265 $Y=0.945 $X2=1.525 $Y2=1.56
cc_119 N_A_M1001_g Y 0.00511826f $X=1.265 $Y=3.825 $X2=1.525 $Y2=1.56
cc_120 N_A_c_178_n Y 0.0051471f $X=1.325 $Y=1.83 $X2=1.525 $Y2=1.56
cc_121 N_A_c_179_n Y 0.012418f $X=1.14 $Y=3.07 $X2=1.525 $Y2=1.56
cc_122 N_A_c_180_n Y 0.0167787f $X=1.325 $Y=1.83 $X2=1.525 $Y2=1.56
cc_123 N_A_M1005_g N_Y_c_228_n 0.00686905f $X=1.265 $Y=0.945 $X2=1.48 $Y2=1.22
cc_124 N_A_c_178_n N_Y_c_228_n 0.00129509f $X=1.325 $Y=1.83 $X2=1.48 $Y2=1.22
cc_125 N_A_c_180_n N_Y_c_228_n 0.00203451f $X=1.325 $Y=1.83 $X2=1.48 $Y2=1.22
cc_126 N_A_M1001_g N_Y_c_230_n 0.00445157f $X=1.265 $Y=3.825 $X2=1.48 $Y2=2.33
cc_127 N_A_c_178_n N_Y_c_230_n 0.00138163f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
cc_128 N_A_c_179_n N_Y_c_230_n 0.0031919f $X=1.14 $Y=3.07 $X2=1.48 $Y2=2.33
cc_129 N_A_c_180_n N_Y_c_230_n 0.00227834f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
