* File: sky130_osu_sc_15T_ls__oai22_l.pxi.spice
* Created: Fri Nov 12 14:59:03 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%GND N_GND_M1005_d N_GND_M1005_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_15T_LS__OAI22_L%GND
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%VDD N_VDD_M1001_s N_VDD_M1004_d N_VDD_M1001_b
+ N_VDD_c_48_p N_VDD_c_49_p N_VDD_c_67_p VDD N_VDD_c_50_p
+ PM_SKY130_OSU_SC_15T_LS__OAI22_L%VDD
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%A0 N_A0_c_73_n N_A0_M1005_g N_A0_M1001_g
+ N_A0_c_77_n N_A0_c_78_n N_A0_c_79_n N_A0_c_80_n A0
+ PM_SKY130_OSU_SC_15T_LS__OAI22_L%A0
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%A1 N_A1_M1007_g N_A1_M1000_g N_A1_c_113_n
+ N_A1_c_114_n N_A1_c_115_n A1 PM_SKY130_OSU_SC_15T_LS__OAI22_L%A1
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%B0 N_B0_M1002_g N_B0_M1003_g N_B0_c_164_n
+ N_B0_c_165_n N_B0_c_166_n B0 PM_SKY130_OSU_SC_15T_LS__OAI22_L%B0
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%B1 N_B1_M1004_g N_B1_M1006_g N_B1_c_212_n
+ N_B1_c_213_n N_B1_c_214_n N_B1_c_215_n B1 PM_SKY130_OSU_SC_15T_LS__OAI22_L%B1
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%Y N_Y_M1002_d N_Y_M1007_d N_Y_c_246_n
+ N_Y_c_258_n N_Y_c_250_n N_Y_c_285_p N_Y_c_242_n N_Y_c_277_n N_Y_c_243_n
+ N_Y_c_244_n Y PM_SKY130_OSU_SC_15T_LS__OAI22_L%Y
x_PM_SKY130_OSU_SC_15T_LS__OAI22_L%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1000_d N_A_27_115#_M1006_d N_A_27_115#_c_289_n
+ N_A_27_115#_c_292_n N_A_27_115#_c_302_n N_A_27_115#_c_294_n
+ N_A_27_115#_c_296_n N_A_27_115#_c_299_n
+ PM_SKY130_OSU_SC_15T_LS__OAI22_L%A_27_115#
cc_1 N_GND_M1005_b N_A0_c_73_n 0.0246907f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.44
cc_2 N_GND_c_2_p N_A0_c_73_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.44
cc_3 N_GND_c_3_p N_A0_c_73_n 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=1.44
cc_4 N_GND_c_4_p N_A0_c_73_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=1.44
cc_5 N_GND_M1005_b N_A0_c_77_n 0.0245194f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.515
cc_6 N_GND_M1005_b N_A0_c_78_n 0.0342831f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.5
cc_7 N_GND_M1005_b N_A0_c_79_n 0.0617326f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.335
cc_8 N_GND_M1005_b N_A0_c_80_n 0.0028102f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.5
cc_9 N_GND_M1005_b N_A1_M1007_g 0.0270201f $X=-0.045 $Y=0 $X2=0.835 $Y2=3.825
cc_10 N_GND_M1005_b N_A1_M1000_g 0.044324f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.945
cc_11 N_GND_c_3_p N_A1_M1000_g 0.00153861f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.945
cc_12 N_GND_c_4_p N_A1_M1000_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.905 $Y2=0.945
cc_13 N_GND_M1005_b N_A1_c_113_n 0.0318892f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.96
cc_14 N_GND_M1005_b N_A1_c_114_n 0.00628302f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.96
cc_15 N_GND_M1005_b N_A1_c_115_n 0.00134829f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.7
cc_16 N_GND_M1005_b A1 0.00271527f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.7
cc_17 N_GND_M1005_b N_B0_M1002_g 0.0223952f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.945
cc_18 N_GND_c_4_p N_B0_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335 $Y2=0.945
cc_19 N_GND_M1005_b N_B0_M1003_g 0.0427388f $X=-0.045 $Y=0 $X2=1.335 $Y2=3.825
cc_20 N_GND_M1005_b N_B0_c_164_n 0.0287877f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.64
cc_21 N_GND_M1005_b N_B0_c_165_n 0.00502228f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.33
cc_22 N_GND_M1005_b N_B0_c_166_n 0.00423567f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.64
cc_23 N_GND_M1005_b B0 0.0129888f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.33
cc_24 N_GND_M1005_b N_B1_M1006_g 0.0524354f $X=-0.045 $Y=0 $X2=1.765 $Y2=0.945
cc_25 N_GND_c_4_p N_B1_M1006_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765 $Y2=0.945
cc_26 N_GND_M1005_b N_B1_c_212_n 0.0319209f $X=-0.045 $Y=0 $X2=1.73 $Y2=2.55
cc_27 N_GND_M1005_b N_B1_c_213_n 0.00983533f $X=-0.045 $Y=0 $X2=1.73 $Y2=2.7
cc_28 N_GND_M1005_b N_B1_c_214_n 0.0576281f $X=-0.045 $Y=0 $X2=2.005 $Y2=1.965
cc_29 N_GND_M1005_b N_B1_c_215_n 0.0125315f $X=-0.045 $Y=0 $X2=2.005 $Y2=1.965
cc_30 N_GND_M1005_b B1 0.00895888f $X=-0.045 $Y=0 $X2=2.005 $Y2=1.965
cc_31 N_GND_M1005_b N_Y_c_242_n 0.00762457f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.59
cc_32 N_GND_M1005_b N_Y_c_243_n 0.00196399f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.475
cc_33 N_GND_M1005_b N_Y_c_244_n 5.70233e-19 $X=-0.045 $Y=0 $X2=1.665 $Y2=1.22
cc_34 N_GND_M1005_b Y 0.0039506f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.59
cc_35 N_GND_M1005_b N_A_27_115#_c_289_n 0.0015601f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_36 N_GND_c_2_p N_A_27_115#_c_289_n 0.00735421f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_37 N_GND_c_4_p N_A_27_115#_c_289_n 0.00476028f $X=1.7 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_38 N_GND_M1005_d N_A_27_115#_c_292_n 0.00542913f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.16
cc_39 N_GND_c_3_p N_A_27_115#_c_292_n 0.0135055f $X=0.69 $Y=0.74 $X2=1.035
+ $Y2=1.16
cc_40 N_GND_M1005_b N_A_27_115#_c_294_n 0.0476186f $X=-0.045 $Y=0 $X2=1.895
+ $Y2=0.56
cc_41 N_GND_c_4_p N_A_27_115#_c_294_n 0.0197787f $X=1.7 $Y=0.19 $X2=1.895
+ $Y2=0.56
cc_42 N_GND_M1005_b N_A_27_115#_c_296_n 0.0145317f $X=-0.045 $Y=0 $X2=1.205
+ $Y2=0.56
cc_43 N_GND_c_3_p N_A_27_115#_c_296_n 0.0062002f $X=0.69 $Y=0.74 $X2=1.205
+ $Y2=0.56
cc_44 N_GND_c_4_p N_A_27_115#_c_296_n 0.00506617f $X=1.7 $Y=0.19 $X2=1.205
+ $Y2=0.56
cc_45 N_GND_M1005_b N_A_27_115#_c_299_n 0.0170548f $X=-0.045 $Y=0 $X2=1.98
+ $Y2=0.56
cc_46 N_GND_c_4_p N_A_27_115#_c_299_n 0.00495178f $X=1.7 $Y=0.19 $X2=1.98
+ $Y2=0.56
cc_47 N_VDD_M1001_b N_A0_M1001_g 0.0208474f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_48 N_VDD_c_48_p N_A0_M1001_g 0.00751602f $X=0.26 $Y=3.885 $X2=0.475 $Y2=3.825
cc_49 N_VDD_c_49_p N_A0_M1001_g 0.00496961f $X=1.825 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_50 N_VDD_c_50_p N_A0_M1001_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.475 $Y2=3.825
cc_51 N_VDD_M1001_b N_A0_c_78_n 0.0059005f $X=-0.045 $Y=2.645 $X2=0.415 $Y2=2.5
cc_52 N_VDD_M1001_s N_A0_c_80_n 0.00849866f $X=0.135 $Y=2.825 $X2=0.415 $Y2=2.5
cc_53 N_VDD_M1001_b N_A0_c_80_n 0.00549657f $X=-0.045 $Y=2.645 $X2=0.415 $Y2=2.5
cc_54 N_VDD_c_48_p N_A0_c_80_n 2.89251e-19 $X=0.26 $Y=3.885 $X2=0.415 $Y2=2.5
cc_55 N_VDD_M1001_s A0 0.0139414f $X=0.135 $Y=2.825 $X2=0.415 $Y2=3.07
cc_56 N_VDD_c_48_p A0 0.00289954f $X=0.26 $Y=3.885 $X2=0.415 $Y2=3.07
cc_57 N_VDD_M1001_b N_A1_M1007_g 0.019001f $X=-0.045 $Y=2.645 $X2=0.835
+ $Y2=3.825
cc_58 N_VDD_c_49_p N_A1_M1007_g 0.00496961f $X=1.825 $Y=5.397 $X2=0.835
+ $Y2=3.825
cc_59 N_VDD_c_50_p N_A1_M1007_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.835 $Y2=3.825
cc_60 N_VDD_M1001_b N_A1_c_115_n 0.00395559f $X=-0.045 $Y=2.645 $X2=0.895
+ $Y2=2.7
cc_61 N_VDD_M1001_b A1 0.00722999f $X=-0.045 $Y=2.645 $X2=0.895 $Y2=2.7
cc_62 N_VDD_M1001_b N_B0_M1003_g 0.0209279f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=3.825
cc_63 N_VDD_c_49_p N_B0_M1003_g 0.00496961f $X=1.825 $Y=5.397 $X2=1.335
+ $Y2=3.825
cc_64 N_VDD_c_50_p N_B0_M1003_g 0.00429146f $X=1.7 $Y=5.36 $X2=1.335 $Y2=3.825
cc_65 N_VDD_M1001_b N_B1_c_213_n 0.0286771f $X=-0.045 $Y=2.645 $X2=1.73 $Y2=2.7
cc_66 N_VDD_c_49_p N_B1_c_213_n 0.00496961f $X=1.825 $Y=5.397 $X2=1.73 $Y2=2.7
cc_67 N_VDD_c_67_p N_B1_c_213_n 0.00751602f $X=1.91 $Y=3.885 $X2=1.73 $Y2=2.7
cc_68 N_VDD_c_50_p N_B1_c_213_n 0.00429146f $X=1.7 $Y=5.36 $X2=1.73 $Y2=2.7
cc_69 N_VDD_M1001_b N_Y_c_246_n 0.00201035f $X=-0.045 $Y=2.645 $X2=1.085
+ $Y2=3.545
cc_70 N_VDD_c_49_p N_Y_c_246_n 0.00454108f $X=1.825 $Y=5.397 $X2=1.085 $Y2=3.545
cc_71 N_VDD_c_50_p N_Y_c_246_n 0.00436053f $X=1.7 $Y=5.36 $X2=1.085 $Y2=3.545
cc_72 N_VDD_M1001_b N_Y_c_242_n 0.00136067f $X=-0.045 $Y=2.645 $X2=1.665
+ $Y2=1.59
cc_73 N_A0_c_78_n N_A1_M1007_g 0.157986f $X=0.415 $Y=2.5 $X2=0.835 $Y2=3.825
cc_74 N_A0_c_79_n N_A1_M1007_g 0.00799469f $X=0.415 $Y=2.335 $X2=0.835 $Y2=3.825
cc_75 N_A0_c_80_n N_A1_M1007_g 0.00302464f $X=0.415 $Y=2.5 $X2=0.835 $Y2=3.825
cc_76 A0 N_A1_M1007_g 0.00376364f $X=0.415 $Y=3.07 $X2=0.835 $Y2=3.825
cc_77 N_A0_c_73_n N_A1_M1000_g 0.0354622f $X=0.475 $Y=1.44 $X2=0.905 $Y2=0.945
cc_78 N_A0_c_79_n N_A1_M1000_g 0.00744899f $X=0.415 $Y=2.335 $X2=0.905 $Y2=0.945
cc_79 N_A0_c_79_n N_A1_c_113_n 0.0167307f $X=0.415 $Y=2.335 $X2=0.815 $Y2=1.96
cc_80 N_A0_c_78_n N_A1_c_114_n 0.00128494f $X=0.415 $Y=2.5 $X2=0.815 $Y2=1.96
cc_81 N_A0_c_79_n N_A1_c_114_n 0.00640175f $X=0.415 $Y=2.335 $X2=0.815 $Y2=1.96
cc_82 N_A0_c_80_n N_A1_c_114_n 0.0241512f $X=0.415 $Y=2.5 $X2=0.815 $Y2=1.96
cc_83 N_A0_M1001_g N_A1_c_115_n 0.00128494f $X=0.475 $Y=3.825 $X2=0.895 $Y2=2.7
cc_84 N_A0_M1001_g A1 4.3358e-19 $X=0.475 $Y=3.825 $X2=0.895 $Y2=2.7
cc_85 N_A0_c_80_n A1 0.00249278f $X=0.415 $Y=2.5 $X2=0.895 $Y2=2.7
cc_86 A0 A_110_565# 0.0129699f $X=0.415 $Y=3.07 $X2=0.55 $Y2=2.825
cc_87 N_A0_c_80_n N_Y_c_250_n 0.00152664f $X=0.415 $Y=2.5 $X2=1.17 $Y2=3.155
cc_88 A0 N_Y_c_250_n 0.00392194f $X=0.415 $Y=3.07 $X2=1.17 $Y2=3.155
cc_89 N_A0_c_73_n N_A_27_115#_c_292_n 0.0200828f $X=0.475 $Y=1.44 $X2=1.035
+ $Y2=1.16
cc_90 N_A0_c_77_n N_A_27_115#_c_302_n 0.00299014f $X=0.475 $Y=1.515 $X2=0.345
+ $Y2=1.16
cc_91 N_A1_M1000_g N_B0_M1002_g 0.0275149f $X=0.905 $Y=0.945 $X2=1.335 $Y2=0.945
cc_92 N_A1_M1007_g N_B0_M1003_g 0.0467845f $X=0.835 $Y=3.825 $X2=1.335 $Y2=3.825
cc_93 N_A1_M1000_g N_B0_M1003_g 0.0122699f $X=0.905 $Y=0.945 $X2=1.335 $Y2=3.825
cc_94 N_A1_c_114_n N_B0_M1003_g 0.00184175f $X=0.815 $Y=1.96 $X2=1.335 $Y2=3.825
cc_95 N_A1_c_115_n N_B0_M1003_g 0.00125927f $X=0.895 $Y=2.7 $X2=1.335 $Y2=3.825
cc_96 A1 N_B0_M1003_g 0.0039398f $X=0.895 $Y=2.7 $X2=1.335 $Y2=3.825
cc_97 N_A1_M1000_g N_B0_c_164_n 0.0194178f $X=0.905 $Y=0.945 $X2=1.325 $Y2=1.64
cc_98 N_A1_M1007_g N_B0_c_165_n 0.00190813f $X=0.835 $Y=3.825 $X2=1.2 $Y2=2.33
cc_99 N_A1_M1000_g N_B0_c_165_n 0.00207047f $X=0.905 $Y=0.945 $X2=1.2 $Y2=2.33
cc_100 N_A1_c_114_n N_B0_c_165_n 0.0340786f $X=0.815 $Y=1.96 $X2=1.2 $Y2=2.33
cc_101 N_A1_M1000_g N_B0_c_166_n 0.00747606f $X=0.905 $Y=0.945 $X2=1.325
+ $Y2=1.64
cc_102 N_A1_c_114_n N_B0_c_166_n 5.67333e-19 $X=0.815 $Y=1.96 $X2=1.325 $Y2=1.64
cc_103 N_A1_M1007_g B0 0.00416458f $X=0.835 $Y=3.825 $X2=1.2 $Y2=2.33
cc_104 N_A1_c_113_n B0 0.00100952f $X=0.815 $Y=1.96 $X2=1.2 $Y2=2.33
cc_105 N_A1_c_114_n B0 0.00821238f $X=0.815 $Y=1.96 $X2=1.2 $Y2=2.33
cc_106 N_A1_c_115_n B0 2.4196e-19 $X=0.895 $Y=2.7 $X2=1.2 $Y2=2.33
cc_107 A1 B0 0.0191116f $X=0.895 $Y=2.7 $X2=1.2 $Y2=2.33
cc_108 N_A1_M1007_g N_Y_c_246_n 0.0178366f $X=0.835 $Y=3.825 $X2=1.085 $Y2=3.545
cc_109 N_A1_M1007_g N_Y_c_250_n 0.00383489f $X=0.835 $Y=3.825 $X2=1.17 $Y2=3.155
cc_110 A1 N_Y_c_250_n 0.00669635f $X=0.895 $Y=2.7 $X2=1.17 $Y2=3.155
cc_111 N_A1_c_115_n N_Y_c_242_n 0.00278415f $X=0.895 $Y=2.7 $X2=1.665 $Y2=1.59
cc_112 A1 N_Y_c_242_n 0.00663666f $X=0.895 $Y=2.7 $X2=1.665 $Y2=1.59
cc_113 N_A1_M1000_g N_A_27_115#_c_292_n 0.0176257f $X=0.905 $Y=0.945 $X2=1.035
+ $Y2=1.16
cc_114 N_A1_c_113_n N_A_27_115#_c_292_n 0.0022598f $X=0.815 $Y=1.96 $X2=1.035
+ $Y2=1.16
cc_115 N_A1_c_114_n N_A_27_115#_c_292_n 0.0046765f $X=0.815 $Y=1.96 $X2=1.035
+ $Y2=1.16
cc_116 N_A1_M1000_g N_A_27_115#_c_296_n 0.0012781f $X=0.905 $Y=0.945 $X2=1.205
+ $Y2=0.56
cc_117 N_B0_M1002_g N_B1_M1006_g 0.0284495f $X=1.335 $Y=0.945 $X2=1.765
+ $Y2=0.945
cc_118 N_B0_c_164_n N_B1_M1006_g 0.0181174f $X=1.325 $Y=1.64 $X2=1.765 $Y2=0.945
cc_119 N_B0_c_166_n N_B1_M1006_g 4.38138e-19 $X=1.325 $Y=1.64 $X2=1.765
+ $Y2=0.945
cc_120 N_B0_M1003_g N_B1_c_213_n 0.143903f $X=1.335 $Y=3.825 $X2=1.73 $Y2=2.7
cc_121 N_B0_M1003_g N_B1_c_214_n 0.0302551f $X=1.335 $Y=3.825 $X2=2.005
+ $Y2=1.965
cc_122 N_B0_c_165_n N_B1_c_214_n 6.71671e-19 $X=1.2 $Y=2.33 $X2=2.005 $Y2=1.965
cc_123 N_B0_M1003_g N_Y_c_246_n 0.0178366f $X=1.335 $Y=3.825 $X2=1.085 $Y2=3.545
cc_124 N_B0_M1003_g N_Y_c_258_n 0.018662f $X=1.335 $Y=3.825 $X2=1.58 $Y2=3.155
cc_125 N_B0_c_165_n N_Y_c_258_n 0.00149445f $X=1.2 $Y=2.33 $X2=1.58 $Y2=3.155
cc_126 N_B0_c_165_n N_Y_c_250_n 9.67274e-19 $X=1.2 $Y=2.33 $X2=1.17 $Y2=3.155
cc_127 N_B0_M1003_g N_Y_c_242_n 0.0112817f $X=1.335 $Y=3.825 $X2=1.665 $Y2=1.59
cc_128 N_B0_c_164_n N_Y_c_242_n 0.0017101f $X=1.325 $Y=1.64 $X2=1.665 $Y2=1.59
cc_129 N_B0_c_165_n N_Y_c_242_n 0.0251114f $X=1.2 $Y=2.33 $X2=1.665 $Y2=1.59
cc_130 N_B0_c_166_n N_Y_c_242_n 0.0203888f $X=1.325 $Y=1.64 $X2=1.665 $Y2=1.59
cc_131 B0 N_Y_c_242_n 0.00640554f $X=1.2 $Y=2.33 $X2=1.665 $Y2=1.59
cc_132 N_B0_M1002_g N_Y_c_243_n 0.00182993f $X=1.335 $Y=0.945 $X2=1.665
+ $Y2=1.475
cc_133 N_B0_M1002_g N_Y_c_244_n 4.93282e-19 $X=1.335 $Y=0.945 $X2=1.665 $Y2=1.22
cc_134 N_B0_c_164_n Y 0.00379994f $X=1.325 $Y=1.64 $X2=1.665 $Y2=1.59
cc_135 N_B0_c_166_n Y 0.00757027f $X=1.325 $Y=1.64 $X2=1.665 $Y2=1.59
cc_136 N_B0_c_164_n N_A_27_115#_c_292_n 3.3129e-19 $X=1.325 $Y=1.64 $X2=1.035
+ $Y2=1.16
cc_137 N_B0_c_166_n N_A_27_115#_c_292_n 0.00613522f $X=1.325 $Y=1.64 $X2=1.035
+ $Y2=1.16
cc_138 N_B0_M1002_g N_A_27_115#_c_294_n 0.0133229f $X=1.335 $Y=0.945 $X2=1.895
+ $Y2=0.56
cc_139 N_B1_c_213_n N_Y_c_258_n 0.0176551f $X=1.73 $Y=2.7 $X2=1.58 $Y2=3.155
cc_140 N_B1_M1006_g N_Y_c_242_n 0.0109199f $X=1.765 $Y=0.945 $X2=1.665 $Y2=1.59
cc_141 N_B1_c_212_n N_Y_c_242_n 0.0207198f $X=1.73 $Y=2.55 $X2=1.665 $Y2=1.59
cc_142 N_B1_c_213_n N_Y_c_242_n 0.0284849f $X=1.73 $Y=2.7 $X2=1.665 $Y2=1.59
cc_143 N_B1_c_214_n N_Y_c_242_n 0.00825017f $X=2.005 $Y=1.965 $X2=1.665 $Y2=1.59
cc_144 N_B1_c_215_n N_Y_c_242_n 0.0203078f $X=2.005 $Y=1.965 $X2=1.665 $Y2=1.59
cc_145 B1 N_Y_c_242_n 0.00704472f $X=2.005 $Y=1.965 $X2=1.665 $Y2=1.59
cc_146 N_B1_M1006_g N_Y_c_277_n 0.00669883f $X=1.765 $Y=0.945 $X2=1.665 $Y2=1.22
cc_147 N_B1_M1006_g N_Y_c_243_n 0.00517857f $X=1.765 $Y=0.945 $X2=1.665
+ $Y2=1.475
cc_148 N_B1_M1006_g N_Y_c_244_n 0.0106956f $X=1.765 $Y=0.945 $X2=1.665 $Y2=1.22
cc_149 N_B1_M1006_g Y 0.00959656f $X=1.765 $Y=0.945 $X2=1.665 $Y2=1.59
cc_150 B1 Y 0.00540133f $X=2.005 $Y=1.965 $X2=1.665 $Y2=1.59
cc_151 N_B1_M1006_g N_A_27_115#_c_294_n 0.0106313f $X=1.765 $Y=0.945 $X2=1.895
+ $Y2=0.56
cc_152 N_B1_M1006_g N_A_27_115#_c_299_n 8.86565e-19 $X=1.765 $Y=0.945 $X2=1.98
+ $Y2=0.56
cc_153 N_Y_c_258_n A_282_565# 0.00732587f $X=1.58 $Y=3.155 $X2=1.41 $Y2=2.825
cc_154 N_Y_c_244_n N_A_27_115#_c_292_n 0.00102777f $X=1.665 $Y=1.22 $X2=1.035
+ $Y2=1.16
cc_155 N_Y_M1002_d N_A_27_115#_c_294_n 0.00177252f $X=1.41 $Y=0.575 $X2=1.895
+ $Y2=0.56
cc_156 N_Y_c_285_p N_A_27_115#_c_294_n 0.0113096f $X=1.55 $Y=0.99 $X2=1.895
+ $Y2=0.56
cc_157 N_Y_c_277_n N_A_27_115#_c_294_n 0.00131309f $X=1.665 $Y=1.22 $X2=1.895
+ $Y2=0.56
cc_158 N_Y_c_244_n N_A_27_115#_c_294_n 0.0049508f $X=1.665 $Y=1.22 $X2=1.895
+ $Y2=0.56
