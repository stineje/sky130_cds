* File: sky130_osu_sc_12T_ms__and2_8.pex.spice
* Created: Fri Nov 12 15:20:43 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__AND2_8%GND 1 2 3 4 5 63 65 73 75 82 84 91 93
+ 100 102 110 123 125
r146 123 125 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r147 108 110 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.56 $Y2=0.755
r148 102 108 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.475
+ $Y=0.152 $X2=4.56 $Y2=0.305
r149 98 100 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.755
r150 94 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r151 89 116 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r152 89 91 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.755
r153 85 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r154 84 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r155 80 115 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r156 80 82 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r157 75 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r158 71 73 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.755
r159 63 125 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r160 63 123 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r161 63 98 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.7 $Y2=0.305
r162 63 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.615 $Y2=0.152
r163 63 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.785 $Y2=0.152
r164 63 71 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r165 63 65 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r166 63 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r167 63 102 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.475 $Y2=0.152
r168 63 103 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=3.785 $Y2=0.152
r169 63 93 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r170 63 94 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r171 63 84 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r172 63 85 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r173 63 75 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r174 63 76 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r175 63 65 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r176 5 110 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.575 $X2=4.56 $Y2=0.755
r177 4 100 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.755
r178 3 91 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.7 $Y=0.575
+ $X2=2.84 $Y2=0.755
r179 2 82 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.755
r180 1 73 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_8%VDD 1 2 3 4 5 6 53 57 59 65 67 73 77 83
+ 87 93 97 104 117 121
r87 117 121 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=4.42 $Y2=4.287
r88 109 117 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r89 104 107 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.56 $Y=2.955
+ $X2=4.56 $Y2=3.635
r90 102 107 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.56 $Y=4.135
+ $X2=4.56 $Y2=3.635
r91 100 121 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=4.25
+ $X2=4.42 $Y2=4.25
r92 98 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=4.287
+ $X2=3.7 $Y2=4.287
r93 98 100 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=4.287
+ $X2=4.42 $Y2=4.287
r94 97 102 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.475 $Y=4.287
+ $X2=4.56 $Y2=4.135
r95 97 100 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.475 $Y=4.287
+ $X2=4.42 $Y2=4.287
r96 93 96 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=2.955 $X2=3.7
+ $Y2=3.635
r97 91 115 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.7 $Y=4.135
+ $X2=3.7 $Y2=4.287
r98 91 96 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.7 $Y=4.135 $X2=3.7
+ $Y2=3.635
r99 88 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=4.287
+ $X2=2.84 $Y2=4.287
r100 88 90 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=4.287
+ $X2=3.06 $Y2=4.287
r101 87 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=4.287
+ $X2=3.7 $Y2=4.287
r102 87 90 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=4.287
+ $X2=3.06 $Y2=4.287
r103 83 86 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=2.955
+ $X2=2.84 $Y2=3.635
r104 81 113 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=4.135
+ $X2=2.84 $Y2=4.287
r105 81 86 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.84 $Y=4.135
+ $X2=2.84 $Y2=3.635
r106 78 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=1.98 $Y2=4.287
r107 78 80 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=2.38 $Y2=4.287
r108 77 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.84 $Y2=4.287
r109 77 80 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.38 $Y2=4.287
r110 73 76 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r111 71 112 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=4.287
r112 71 76 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=3.635
r113 68 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r114 68 70 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r115 67 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.287
r116 67 70 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r117 63 111 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r118 63 65 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.295
r119 60 109 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r120 60 62 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r121 59 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r122 59 62 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r123 55 109 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r124 55 57 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r125 53 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=4.135 $X2=4.42 $Y2=4.22
r126 53 115 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r127 53 90 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r128 53 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r129 53 70 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r130 53 62 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r131 53 109 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r132 6 107 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=2.605 $X2=4.56 $Y2=3.635
r133 6 104 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=2.605 $X2=4.56 $Y2=2.955
r134 5 96 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=3.635
r135 5 93 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=2.955
r136 4 86 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=3.635
r137 4 83 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=2.955
r138 3 76 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r139 3 73 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r140 2 65 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.295
r141 1 57 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_8%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=2.85
+ $X2=0.275 $Y2=2.85
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.85
+ $X2=0.27 $Y2=2.85
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.285
+ $X2=0.27 $Y2=2.85
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.285 $X2=0.27 $Y2=2.285
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.285
+ $X2=0.475 $Y2=2.285
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.45
+ $X2=0.475 $Y2=2.285
r38 5 7 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.475 $Y=2.45
+ $X2=0.475 $Y2=3.235
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=2.285
r40 1 3 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_8%B 3 7 10 14 22
c41 7 0 1.37149e-19 $X=0.905 $Y=3.235
r42 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.48
+ $X2=0.955 $Y2=2.48
r43 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.48
+ $X2=0.95 $Y2=2.48
r44 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=1.945
+ $X2=0.95 $Y2=2.48
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.945 $X2=0.95 $Y2=1.945
r46 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=1.945
+ $X2=0.922 $Y2=2.11
r47 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=1.945
+ $X2=0.922 $Y2=1.78
r48 7 12 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.11
r49 3 11 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.835 $Y=0.835
+ $X2=0.835 $Y2=1.78
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_8%A_27_115# 1 3 11 13 15 17 18 22 24 26 27
+ 28 29 33 35 37 38 40 44 46 48 49 51 55 58 59 61 62 64 68 70 72 73 75 79 81 83
+ 84 86 90 92 94 95 101 102 103 104 105 106 107 108 109 110 111 114 116 117 122
+ 126 128 129 130
c243 68 0 1.33323e-19 $X=3.485 $Y=0.835
c244 55 0 1.33323e-19 $X=3.055 $Y=0.835
c245 44 0 1.33323e-19 $X=2.625 $Y=0.835
c246 33 0 1.33323e-19 $X=2.195 $Y=0.835
c247 22 0 1.33323e-19 $X=1.765 $Y=0.835
r248 129 130 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.065
+ $X2=0.65 $Y2=3.235
r249 124 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.455
+ $X2=0.61 $Y2=1.455
r250 124 126 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.455
+ $X2=1.43 $Y2=1.455
r251 122 130 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.69 $Y=3.295
+ $X2=0.69 $Y2=3.235
r252 118 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=1.455
r253 118 129 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=3.065
r254 116 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.455
+ $X2=0.61 $Y2=1.455
r255 116 117 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.455
+ $X2=0.345 $Y2=1.455
r256 112 117 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.345 $Y2=1.455
r257 112 114 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r258 99 126 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.455 $X2=1.43 $Y2=1.455
r259 97 99 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.455
+ $X2=1.43 $Y2=1.455
r260 96 97 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.455
+ $X2=1.37 $Y2=1.455
r261 92 94 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=4.345 $Y=2.48
+ $X2=4.345 $Y2=3.235
r262 88 90 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.345 $Y=1.29
+ $X2=4.345 $Y2=0.835
r263 87 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=2.405
+ $X2=3.915 $Y2=2.405
r264 86 92 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=2.405
+ $X2=4.345 $Y2=2.48
r265 86 87 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=2.405
+ $X2=3.99 $Y2=2.405
r266 85 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.365
+ $X2=3.915 $Y2=1.365
r267 84 88 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=1.365
+ $X2=4.345 $Y2=1.29
r268 84 85 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.365
+ $X2=3.99 $Y2=1.365
r269 81 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=2.48
+ $X2=3.915 $Y2=2.405
r270 81 83 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.915 $Y=2.48
+ $X2=3.915 $Y2=3.235
r271 77 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=1.29
+ $X2=3.915 $Y2=1.365
r272 77 79 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.915 $Y=1.29
+ $X2=3.915 $Y2=0.835
r273 76 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.405
+ $X2=3.485 $Y2=2.405
r274 75 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.405
+ $X2=3.915 $Y2=2.405
r275 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.405
+ $X2=3.56 $Y2=2.405
r276 74 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.365
+ $X2=3.485 $Y2=1.365
r277 73 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.365
+ $X2=3.915 $Y2=1.365
r278 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.365
+ $X2=3.56 $Y2=1.365
r279 70 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.48
+ $X2=3.485 $Y2=2.405
r280 70 72 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.485 $Y=2.48
+ $X2=3.485 $Y2=3.235
r281 66 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.29
+ $X2=3.485 $Y2=1.365
r282 66 68 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.485 $Y=1.29
+ $X2=3.485 $Y2=0.835
r283 65 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.405
+ $X2=3.055 $Y2=2.405
r284 64 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.405
+ $X2=3.485 $Y2=2.405
r285 64 65 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.405
+ $X2=3.13 $Y2=2.405
r286 63 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.365
+ $X2=3.055 $Y2=1.365
r287 62 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.365
+ $X2=3.485 $Y2=1.365
r288 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.365
+ $X2=3.13 $Y2=1.365
r289 59 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.48
+ $X2=3.055 $Y2=2.405
r290 59 61 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.055 $Y=2.48
+ $X2=3.055 $Y2=3.235
r291 58 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.33
+ $X2=3.055 $Y2=2.405
r292 57 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=1.365
r293 57 58 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=2.33
r294 53 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.29
+ $X2=3.055 $Y2=1.365
r295 53 55 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.055 $Y=1.29
+ $X2=3.055 $Y2=0.835
r296 52 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.405
+ $X2=2.625 $Y2=2.405
r297 51 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.405
+ $X2=3.055 $Y2=2.405
r298 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.405
+ $X2=2.7 $Y2=2.405
r299 50 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.365
+ $X2=2.625 $Y2=1.365
r300 49 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.365
+ $X2=3.055 $Y2=1.365
r301 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.365
+ $X2=2.7 $Y2=1.365
r302 46 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=2.405
r303 46 48 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=3.235
r304 42 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.29
+ $X2=2.625 $Y2=1.365
r305 42 44 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.625 $Y=1.29
+ $X2=2.625 $Y2=0.835
r306 41 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.405
+ $X2=2.195 $Y2=2.405
r307 40 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.625 $Y2=2.405
r308 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.27 $Y2=2.405
r309 39 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.365
+ $X2=2.195 $Y2=1.365
r310 38 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.365
+ $X2=2.625 $Y2=1.365
r311 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.365
+ $X2=2.27 $Y2=1.365
r312 35 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=2.405
r313 35 37 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=3.235
r314 31 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=1.365
r315 31 33 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=0.835
r316 30 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.405
+ $X2=1.765 $Y2=2.405
r317 29 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=2.195 $Y2=2.405
r318 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=1.84 $Y2=2.405
r319 27 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=2.195 $Y2=1.365
r320 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=1.84 $Y2=1.365
r321 24 101 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=2.405
r322 24 26 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r323 20 28 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.84 $Y2=1.365
r324 20 99 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.43 $Y2=1.455
r325 20 22 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=0.835
r326 19 95 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.405
+ $X2=1.352 $Y2=2.405
r327 18 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.405
r328 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.445 $Y2=2.405
r329 17 95 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.33
+ $X2=1.352 $Y2=2.405
r330 16 97 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=1.455
r331 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=2.33
r332 13 95 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.352 $Y2=2.405
r333 13 15 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r334 9 96 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=1.455
r335 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.835
r336 3 122 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.295
r337 1 114 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68
+ 76 82 89 90 92 94 96 99 100 101 102 103 104 105 106 107 110 111 125
c171 110 0 1.33323e-19 $X=4.13 $Y=1.115
c172 104 0 1.33323e-19 $X=3.27 $Y=1.115
c173 101 0 2.66647e-19 $X=2.555 $Y=1
c174 89 0 1.33323e-19 $X=1.55 $Y=1.115
c175 40 0 1.37149e-19 $X=1.55 $Y=2.11
r176 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.995
+ $X2=4.13 $Y2=2.11
r177 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.115
+ $X2=4.13 $Y2=1
r178 110 111 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=4.13 $Y=1.115
+ $X2=4.13 $Y2=1.995
r179 107 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=2.11
+ $X2=3.27 $Y2=2.11
r180 106 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=2.11
+ $X2=4.13 $Y2=2.11
r181 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=2.11
+ $X2=3.415 $Y2=2.11
r182 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.995
+ $X2=3.27 $Y2=2.11
r183 104 121 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.115
+ $X2=3.27 $Y2=1
r184 104 105 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=3.27 $Y=1.115
+ $X2=3.27 $Y2=1.995
r185 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.11
+ $X2=2.41 $Y2=2.11
r186 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.11
+ $X2=3.27 $Y2=2.11
r187 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.11
+ $X2=2.555 $Y2=2.11
r188 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1
+ $X2=2.41 $Y2=1
r189 100 121 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1
+ $X2=3.27 $Y2=1
r190 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1
+ $X2=2.555 $Y2=1
r191 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.995
+ $X2=2.41 $Y2=2.11
r192 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=1
r193 98 99 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=1.995
r194 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.11
+ $X2=1.55 $Y2=2.11
r195 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.11
+ $X2=2.41 $Y2=2.11
r196 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.11
+ $X2=1.695 $Y2=2.11
r197 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1
+ $X2=1.55 $Y2=1
r198 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=2.41 $Y2=1
r199 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=1.695 $Y2=1
r200 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=2.11
r201 90 92 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=1.74
r202 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r203 89 92 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.74
r204 85 87 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.13 $Y=2.955
+ $X2=4.13 $Y2=3.635
r205 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=2.11
+ $X2=4.13 $Y2=2.11
r206 82 85 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=4.13 $Y=2.11
+ $X2=4.13 $Y2=2.955
r207 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=1 $X2=4.13
+ $Y2=1
r208 76 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.13 $Y=0.755
+ $X2=4.13 $Y2=1
r209 71 73 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=2.955
+ $X2=3.27 $Y2=3.635
r210 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.11
+ $X2=3.27 $Y2=2.11
r211 68 71 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.27 $Y=2.11
+ $X2=3.27 $Y2=2.955
r212 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1 $X2=3.27
+ $Y2=1
r213 62 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.27 $Y=0.755
+ $X2=3.27 $Y2=1
r214 57 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=2.955
+ $X2=2.41 $Y2=3.635
r215 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.11
+ $X2=2.41 $Y2=2.11
r216 54 57 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.41 $Y=2.11
+ $X2=2.41 $Y2=2.955
r217 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1 $X2=2.41
+ $Y2=1
r218 48 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.41 $Y=0.755
+ $X2=2.41 $Y2=1
r219 43 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r220 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.11
r221 40 43 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.955
r222 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r223 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r224 12 87 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.605 $X2=4.13 $Y2=3.635
r225 12 85 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.605 $X2=4.13 $Y2=2.955
r226 11 73 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=3.635
r227 11 71 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=2.955
r228 10 59 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=3.635
r229 10 57 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=2.955
r230 9 45 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r231 9 43 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r232 4 76 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.755
r233 3 62 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.755
r234 2 48 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.755
r235 1 34 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
.ends

