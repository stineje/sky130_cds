* File: sky130_osu_sc_12T_hs__and2_4.spice
* Created: Fri Nov 12 15:07:01 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__and2_4.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_4  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 A_110_115# N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_B_M1002_g A_110_115# N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75002 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.09625 PD=0.83 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1001_d N_A_27_115#_M1009_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1010 N_Y_M1010_d N_A_27_115#_M1010_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1010_d N_A_27_115#_M1011_g N_GND_M1011_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1007 N_VDD_M1007_d N_B_M1007_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1007_d N_A_27_115#_M1003_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_27_115#_M1005_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1005_d N_A_27_115#_M1006_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_VDD_M1008_d N_A_27_115#_M1008_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_8 A A PROBETYPE=1
pX14_noxref noxref_9 B B PROBETYPE=1
pX15_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_4.pxi.spice"
*
.ends
*
*
