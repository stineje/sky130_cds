* File: sky130_osu_sc_15T_ms__and2_1.spice
* Created: Fri Nov 12 14:40:03 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__and2_1.pex.spice"
.subckt sky130_osu_sc_15T_ms__and2_1  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 A_110_115# N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1004_b NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.0777 PD=1.09 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1001_d N_GND_M1004_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1295 PD=2.01 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_115#_M1005_d N_A_M1005_g N_VDD_M1005_s N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1002 N_VDD_M1002_d N_B_M1002_g N_A_27_115#_M1005_d N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_VDD_M1002_d N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1005_b NWDIODE A=5.64925 P=9.73
pX7_noxref noxref_8 A A PROBETYPE=1
pX8_noxref noxref_9 B B PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__and2_1.pxi.spice"
*
.ends
*
*
