* File: sky130_osu_sc_12T_ls__dffs_1.pxi.spice
* Created: Fri Nov 12 15:36:23 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%GND N_GND_M1000_d N_GND_M1001_s N_GND_M1021_d
+ N_GND_M1006_d N_GND_M1025_d N_GND_M1008_d N_GND_M1012_b N_GND_c_2_p
+ N_GND_c_24_p N_GND_c_25_p N_GND_c_26_p N_GND_c_27_p N_GND_c_28_p N_GND_c_29_p
+ N_GND_c_30_p N_GND_c_6_p N_GND_c_7_p N_GND_c_33_p N_GND_c_157_p GND
+ N_GND_c_3_p PM_SKY130_OSU_SC_12T_LS__DFFS_1%GND
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%VDD N_VDD_M1009_s N_VDD_M1020_d N_VDD_M1007_s
+ N_VDD_M1014_d N_VDD_M1026_d N_VDD_M1024_s N_VDD_M1016_d N_VDD_M1029_d
+ N_VDD_M1009_b N_VDD_c_218_p N_VDD_c_219_p N_VDD_c_227_p N_VDD_c_228_p
+ N_VDD_c_238_p N_VDD_c_263_p N_VDD_c_248_p N_VDD_c_252_p N_VDD_c_253_p
+ N_VDD_c_254_p N_VDD_c_222_p N_VDD_c_223_p N_VDD_c_293_p N_VDD_c_294_p
+ N_VDD_c_315_p VDD N_VDD_c_220_p PM_SKY130_OSU_SC_12T_LS__DFFS_1%VDD
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%SN N_SN_M1012_g N_SN_M1009_g N_SN_c_334_n
+ N_SN_M1025_g N_SN_M1016_g N_SN_c_339_n N_SN_c_340_n N_SN_c_342_n N_SN_c_343_n
+ N_SN_c_345_n N_SN_c_346_n N_SN_c_363_n SN PM_SKY130_OSU_SC_12T_LS__DFFS_1%SN
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_152_89# N_A_152_89#_M1023_d
+ N_A_152_89#_M1011_d N_A_152_89#_M1000_g N_A_152_89#_M1020_g
+ N_A_152_89#_c_484_n N_A_152_89#_c_485_n N_A_152_89#_c_486_n
+ N_A_152_89#_c_489_n N_A_152_89#_c_501_n N_A_152_89#_c_505_n
+ N_A_152_89#_c_491_n N_A_152_89#_c_507_n N_A_152_89#_c_492_n
+ PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_152_89#
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%D N_D_M1001_g N_D_M1007_g N_D_c_575_n
+ N_D_c_576_n D PM_SKY130_OSU_SC_12T_LS__DFFS_1%D
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%CK N_CK_M1011_g N_CK_M1018_g N_CK_M1010_g
+ N_CK_M1028_g N_CK_M1003_g N_CK_c_611_n N_CK_M1017_g N_CK_c_612_n N_CK_c_613_n
+ N_CK_c_614_n N_CK_c_615_n N_CK_c_618_n N_CK_c_619_n N_CK_c_622_n N_CK_c_623_n
+ N_CK_c_627_n N_CK_c_628_n N_CK_c_629_n N_CK_c_630_n N_CK_c_631_n N_CK_c_632_n
+ N_CK_c_633_n N_CK_c_634_n N_CK_c_635_n N_CK_c_636_n N_CK_c_637_n N_CK_c_638_n
+ N_CK_c_639_n CK PM_SKY130_OSU_SC_12T_LS__DFFS_1%CK
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_27_115# N_A_27_115#_M1012_s
+ N_A_27_115#_M1009_d N_A_27_115#_M1021_g N_A_27_115#_M1014_g
+ N_A_27_115#_c_848_n N_A_27_115#_c_850_n N_A_27_115#_c_851_n
+ N_A_27_115#_c_852_n N_A_27_115#_M1013_g N_A_27_115#_M1005_g
+ N_A_27_115#_c_857_n N_A_27_115#_c_860_n N_A_27_115#_c_861_n
+ N_A_27_115#_c_862_n N_A_27_115#_c_865_n N_A_27_115#_c_867_n
+ N_A_27_115#_c_868_n N_A_27_115#_c_869_n N_A_27_115#_c_870_n
+ N_A_27_115#_c_913_n PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_27_115#
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_428_89# N_A_428_89#_M1003_d
+ N_A_428_89#_M1017_d N_A_428_89#_c_984_n N_A_428_89#_M1023_g
+ N_A_428_89#_c_987_n N_A_428_89#_c_988_n N_A_428_89#_c_989_n
+ N_A_428_89#_M1015_g N_A_428_89#_c_991_n N_A_428_89#_M1022_g
+ N_A_428_89#_c_993_n N_A_428_89#_M1002_g N_A_428_89#_c_997_n
+ N_A_428_89#_c_998_n N_A_428_89#_c_999_n N_A_428_89#_c_1000_n
+ N_A_428_89#_c_1001_n N_A_428_89#_c_1002_n N_A_428_89#_c_1017_n
+ N_A_428_89#_c_1006_n N_A_428_89#_c_1022_n N_A_428_89#_c_1007_n
+ N_A_428_89#_c_1008_n N_A_428_89#_c_1009_n N_A_428_89#_c_1010_n
+ PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_428_89#
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_970_89# N_A_970_89#_M1004_s
+ N_A_970_89#_M1024_d N_A_970_89#_M1006_g N_A_970_89#_M1026_g
+ N_A_970_89#_M1008_g N_A_970_89#_M1029_g N_A_970_89#_c_1185_n
+ N_A_970_89#_c_1187_n N_A_970_89#_c_1188_n N_A_970_89#_c_1189_n
+ N_A_970_89#_c_1194_n N_A_970_89#_c_1195_n N_A_970_89#_c_1196_n
+ N_A_970_89#_c_1197_n N_A_970_89#_c_1198_n N_A_970_89#_c_1201_n
+ N_A_970_89#_c_1202_n N_A_970_89#_c_1203_n N_A_970_89#_c_1204_n
+ N_A_970_89#_c_1207_n N_A_970_89#_c_1208_n N_A_970_89#_c_1209_n
+ N_A_970_89#_c_1210_n N_A_970_89#_c_1211_n N_A_970_89#_c_1212_n
+ N_A_970_89#_c_1213_n PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_970_89#
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_808_115# N_A_808_115#_M1010_d
+ N_A_808_115#_M1022_d N_A_808_115#_M1004_g N_A_808_115#_M1024_g
+ N_A_808_115#_c_1382_n N_A_808_115#_c_1383_n N_A_808_115#_c_1426_n
+ N_A_808_115#_c_1459_n N_A_808_115#_c_1400_n N_A_808_115#_c_1384_n
+ N_A_808_115#_c_1385_n N_A_808_115#_c_1386_n N_A_808_115#_c_1389_n
+ N_A_808_115#_c_1390_n N_A_808_115#_c_1391_n N_A_808_115#_c_1393_n
+ N_A_808_115#_c_1394_n PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_808_115#
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%QN N_QN_M1008_s N_QN_M1029_s N_QN_M1027_g
+ N_QN_M1019_g N_QN_c_1527_n N_QN_c_1528_n N_QN_c_1532_n N_QN_c_1533_n
+ N_QN_c_1535_n N_QN_c_1536_n N_QN_c_1537_n N_QN_c_1538_n QN
+ PM_SKY130_OSU_SC_12T_LS__DFFS_1%QN
x_PM_SKY130_OSU_SC_12T_LS__DFFS_1%Q N_Q_M1027_d N_Q_M1019_d N_Q_c_1610_n
+ N_Q_c_1614_n N_Q_c_1612_n N_Q_c_1613_n N_Q_c_1618_n Q
+ PM_SKY130_OSU_SC_12T_LS__DFFS_1%Q
cc_1 N_GND_M1012_b N_SN_M1012_g 0.0374026f $X=-0.055 $Y=0 $X2=0.475 $Y2=0.755
cc_2 N_GND_c_2_p N_SN_M1012_g 0.00454486f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.755
cc_3 N_GND_c_3_p N_SN_M1012_g 0.00468827f $X=7.815 $Y=0.19 $X2=0.475 $Y2=0.755
cc_4 N_GND_M1012_b N_SN_M1009_g 0.0619433f $X=-0.055 $Y=0 $X2=0.475 $Y2=3.445
cc_5 N_GND_M1012_b N_SN_c_334_n 0.0170242f $X=-0.055 $Y=0 $X2=6.665 $Y2=1.04
cc_6 N_GND_c_6_p N_SN_c_334_n 0.00591263f $X=6.795 $Y=0.152 $X2=6.665 $Y2=1.04
cc_7 N_GND_c_7_p N_SN_c_334_n 0.00502587f $X=6.88 $Y=0.74 $X2=6.665 $Y2=1.04
cc_8 N_GND_c_3_p N_SN_c_334_n 0.00468827f $X=7.815 $Y=0.19 $X2=6.665 $Y2=1.04
cc_9 N_GND_M1012_b N_SN_M1016_g 0.0694085f $X=-0.055 $Y=0 $X2=6.735 $Y2=3.445
cc_10 N_GND_M1012_b N_SN_c_339_n 0.0438182f $X=-0.055 $Y=0 $X2=0.32 $Y2=1.47
cc_11 N_GND_M1012_b N_SN_c_340_n 0.0530634f $X=-0.055 $Y=0 $X2=6.735 $Y2=1.232
cc_12 N_GND_c_7_p N_SN_c_340_n 0.00328003f $X=6.88 $Y=0.74 $X2=6.735 $Y2=1.232
cc_13 N_GND_M1012_b N_SN_c_342_n 0.00303389f $X=-0.055 $Y=0 $X2=0.32 $Y2=1.47
cc_14 N_GND_M1012_b N_SN_c_343_n 0.00373713f $X=-0.055 $Y=0 $X2=6.94 $Y2=1.165
cc_15 N_GND_c_7_p N_SN_c_343_n 0.0112653f $X=6.88 $Y=0.74 $X2=6.94 $Y2=1.165
cc_16 N_GND_M1012_b N_SN_c_345_n 0.00899939f $X=-0.055 $Y=0 $X2=0.32 $Y2=1.415
cc_17 N_GND_M1000_d N_SN_c_346_n 0.00250063f $X=0.91 $Y=0.575 $X2=1.405
+ $Y2=0.985
cc_18 N_GND_M1001_s N_SN_c_346_n 0.00261163f $X=1.515 $Y=0.575 $X2=1.405
+ $Y2=0.985
cc_19 N_GND_M1021_d N_SN_c_346_n 0.00717371f $X=3.25 $Y=0.575 $X2=1.405
+ $Y2=0.985
cc_20 N_GND_M1006_d N_SN_c_346_n 0.0037916f $X=5 $Y=0.575 $X2=1.405 $Y2=0.985
cc_21 N_GND_M1025_d N_SN_c_346_n 0.00269126f $X=6.74 $Y=0.575 $X2=1.405
+ $Y2=0.985
cc_22 N_GND_M1012_b N_SN_c_346_n 0.0213084f $X=-0.055 $Y=0 $X2=1.405 $Y2=0.985
cc_23 N_GND_c_2_p N_SN_c_346_n 0.00267702f $X=0.965 $Y=0.152 $X2=1.405 $Y2=0.985
cc_24 N_GND_c_24_p N_SN_c_346_n 0.00586327f $X=1.05 $Y=0.74 $X2=1.405 $Y2=0.985
cc_25 N_GND_c_25_p N_SN_c_346_n 0.0069593f $X=1.555 $Y=0.152 $X2=1.405 $Y2=0.985
cc_26 N_GND_c_26_p N_SN_c_346_n 0.011817f $X=1.64 $Y=0.755 $X2=1.405 $Y2=0.985
cc_27 N_GND_c_27_p N_SN_c_346_n 0.0191206f $X=3.305 $Y=0.152 $X2=1.405 $Y2=0.985
cc_28 N_GND_c_28_p N_SN_c_346_n 0.00706915f $X=3.39 $Y=0.74 $X2=1.405 $Y2=0.985
cc_29 N_GND_c_29_p N_SN_c_346_n 0.0191175f $X=5.055 $Y=0.152 $X2=1.405 $Y2=0.985
cc_30 N_GND_c_30_p N_SN_c_346_n 0.0140066f $X=5.14 $Y=0.755 $X2=1.405 $Y2=0.985
cc_31 N_GND_c_6_p N_SN_c_346_n 0.0141329f $X=6.795 $Y=0.152 $X2=1.405 $Y2=0.985
cc_32 N_GND_c_7_p N_SN_c_346_n 0.00625311f $X=6.88 $Y=0.74 $X2=1.405 $Y2=0.985
cc_33 N_GND_c_33_p N_SN_c_346_n 0.00117416f $X=7.815 $Y=0.152 $X2=1.405
+ $Y2=0.985
cc_34 N_GND_M1012_b N_SN_c_363_n 0.00243402f $X=-0.055 $Y=0 $X2=0.405 $Y2=0.985
cc_35 N_GND_c_2_p N_SN_c_363_n 0.00122396f $X=0.965 $Y=0.152 $X2=0.405 $Y2=0.985
cc_36 N_GND_M1012_b SN 0.0179639f $X=-0.055 $Y=0 $X2=0.32 $Y2=1.535
cc_37 N_GND_M1012_b N_A_152_89#_M1000_g 0.0571285f $X=-0.055 $Y=0 $X2=0.835
+ $Y2=0.755
cc_38 N_GND_c_2_p N_A_152_89#_M1000_g 0.00591263f $X=0.965 $Y=0.152 $X2=0.835
+ $Y2=0.755
cc_39 N_GND_c_24_p N_A_152_89#_M1000_g 0.00502587f $X=1.05 $Y=0.74 $X2=0.835
+ $Y2=0.755
cc_40 N_GND_c_3_p N_A_152_89#_M1000_g 0.00468827f $X=7.815 $Y=0.19 $X2=0.835
+ $Y2=0.755
cc_41 N_GND_M1012_b N_A_152_89#_M1020_g 0.0211692f $X=-0.055 $Y=0 $X2=0.905
+ $Y2=3.445
cc_42 N_GND_M1012_b N_A_152_89#_c_484_n 0.0441133f $X=-0.055 $Y=0 $X2=1.03
+ $Y2=1.925
cc_43 N_GND_M1012_b N_A_152_89#_c_485_n 0.0134726f $X=-0.055 $Y=0 $X2=1.03
+ $Y2=1.925
cc_44 N_GND_M1012_b N_A_152_89#_c_486_n 0.0259206f $X=-0.055 $Y=0 $X2=2.33
+ $Y2=1.285
cc_45 N_GND_c_24_p N_A_152_89#_c_486_n 6.10944e-19 $X=1.05 $Y=0.74 $X2=2.33
+ $Y2=1.285
cc_46 N_GND_c_26_p N_A_152_89#_c_486_n 0.00677569f $X=1.64 $Y=0.755 $X2=2.33
+ $Y2=1.285
cc_47 N_GND_M1012_b N_A_152_89#_c_489_n 0.00339036f $X=-0.055 $Y=0 $X2=1.115
+ $Y2=1.285
cc_48 N_GND_c_24_p N_A_152_89#_c_489_n 0.00546659f $X=1.05 $Y=0.74 $X2=1.115
+ $Y2=1.285
cc_49 N_GND_M1012_b N_A_152_89#_c_491_n 0.00198494f $X=-0.055 $Y=0 $X2=2.415
+ $Y2=1.2
cc_50 N_GND_M1012_b N_A_152_89#_c_492_n 0.00311983f $X=-0.055 $Y=0 $X2=2.415
+ $Y2=0.755
cc_51 N_GND_c_27_p N_A_152_89#_c_492_n 0.0146229f $X=3.305 $Y=0.152 $X2=2.415
+ $Y2=0.755
cc_52 N_GND_c_3_p N_A_152_89#_c_492_n 0.0098977f $X=7.815 $Y=0.19 $X2=2.415
+ $Y2=0.755
cc_53 N_GND_M1012_b N_D_M1001_g 0.0421748f $X=-0.055 $Y=0 $X2=1.855 $Y2=0.835
cc_54 N_GND_c_26_p N_D_M1001_g 0.00509529f $X=1.64 $Y=0.755 $X2=1.855 $Y2=0.835
cc_55 N_GND_c_27_p N_D_M1001_g 0.00606474f $X=3.305 $Y=0.152 $X2=1.855 $Y2=0.835
cc_56 N_GND_c_3_p N_D_M1001_g 0.00468827f $X=7.815 $Y=0.19 $X2=1.855 $Y2=0.835
cc_57 N_GND_M1012_b N_D_M1007_g 0.0365658f $X=-0.055 $Y=0 $X2=1.855 $Y2=3.235
cc_58 N_GND_M1012_b N_D_c_575_n 0.0315489f $X=-0.055 $Y=0 $X2=1.915 $Y2=1.74
cc_59 N_GND_M1012_b N_D_c_576_n 0.00311208f $X=-0.055 $Y=0 $X2=1.915 $Y2=1.74
cc_60 N_GND_M1012_b D 0.0139986f $X=-0.055 $Y=0 $X2=1.915 $Y2=1.74
cc_61 N_GND_M1012_b N_CK_c_611_n 0.030775f $X=-0.055 $Y=0 $X2=5.355 $Y2=2.45
cc_62 N_GND_M1012_b N_CK_c_612_n 0.0444354f $X=-0.055 $Y=0 $X2=5.41 $Y2=2.12
cc_63 N_GND_M1012_b N_CK_c_613_n 0.0244095f $X=-0.055 $Y=0 $X2=2.275 $Y2=2.285
cc_64 N_GND_M1012_b N_CK_c_614_n 0.0254608f $X=-0.055 $Y=0 $X2=2.755 $Y2=1.37
cc_65 N_GND_M1012_b N_CK_c_615_n 0.0173906f $X=-0.055 $Y=0 $X2=2.755 $Y2=1.205
cc_66 N_GND_c_27_p N_CK_c_615_n 0.00606474f $X=3.305 $Y=0.152 $X2=2.755
+ $Y2=1.205
cc_67 N_GND_c_3_p N_CK_c_615_n 0.00468827f $X=7.815 $Y=0.19 $X2=2.755 $Y2=1.205
cc_68 N_GND_M1012_b N_CK_c_618_n 0.026814f $X=-0.055 $Y=0 $X2=4.025 $Y2=1.37
cc_69 N_GND_M1012_b N_CK_c_619_n 0.0174883f $X=-0.055 $Y=0 $X2=4.025 $Y2=1.205
cc_70 N_GND_c_29_p N_CK_c_619_n 0.00606474f $X=5.055 $Y=0.152 $X2=4.025
+ $Y2=1.205
cc_71 N_GND_c_3_p N_CK_c_619_n 0.00468827f $X=7.815 $Y=0.19 $X2=4.025 $Y2=1.205
cc_72 N_GND_M1012_b N_CK_c_622_n 0.0218864f $X=-0.055 $Y=0 $X2=4.505 $Y2=2.285
cc_73 N_GND_M1012_b N_CK_c_623_n 0.0206446f $X=-0.055 $Y=0 $X2=5.382 $Y2=1.205
cc_74 N_GND_c_30_p N_CK_c_623_n 0.00311745f $X=5.14 $Y=0.755 $X2=5.382 $Y2=1.205
cc_75 N_GND_c_6_p N_CK_c_623_n 0.00606474f $X=6.795 $Y=0.152 $X2=5.382 $Y2=1.205
cc_76 N_GND_c_3_p N_CK_c_623_n 0.00468827f $X=7.815 $Y=0.19 $X2=5.382 $Y2=1.205
cc_77 N_GND_M1012_b N_CK_c_627_n 0.0132119f $X=-0.055 $Y=0 $X2=5.382 $Y2=1.355
cc_78 N_GND_M1012_b N_CK_c_628_n 0.00609317f $X=-0.055 $Y=0 $X2=2.67 $Y2=2.11
cc_79 N_GND_M1012_b N_CK_c_629_n 0.00922239f $X=-0.055 $Y=0 $X2=2.755 $Y2=1.37
cc_80 N_GND_M1012_b N_CK_c_630_n 0.00776632f $X=-0.055 $Y=0 $X2=4.025 $Y2=1.37
cc_81 N_GND_M1012_b N_CK_c_631_n 0.00482391f $X=-0.055 $Y=0 $X2=4.42 $Y2=2.11
cc_82 N_GND_M1012_b N_CK_c_632_n 5.00459e-19 $X=-0.055 $Y=0 $X2=4.11 $Y2=2.11
cc_83 N_GND_M1012_b N_CK_c_633_n 6.56762e-19 $X=-0.055 $Y=0 $X2=5.5 $Y2=2.11
cc_84 N_GND_M1012_b N_CK_c_634_n 0.00276905f $X=-0.055 $Y=0 $X2=2.275 $Y2=2.11
cc_85 N_GND_M1012_b N_CK_c_635_n 0.00120157f $X=-0.055 $Y=0 $X2=4.505 $Y2=2.11
cc_86 N_GND_M1012_b N_CK_c_636_n 0.033889f $X=-0.055 $Y=0 $X2=4.36 $Y2=2.11
cc_87 N_GND_M1012_b N_CK_c_637_n 0.00714094f $X=-0.055 $Y=0 $X2=2.42 $Y2=2.11
cc_88 N_GND_M1012_b N_CK_c_638_n 0.013834f $X=-0.055 $Y=0 $X2=5.355 $Y2=2.11
cc_89 N_GND_M1012_b N_CK_c_639_n 0.00256396f $X=-0.055 $Y=0 $X2=4.65 $Y2=2.11
cc_90 N_GND_M1012_b CK 0.00137114f $X=-0.055 $Y=0 $X2=5.5 $Y2=2.11
cc_91 N_GND_M1012_b N_A_27_115#_M1021_g 0.0171926f $X=-0.055 $Y=0 $X2=3.175
+ $Y2=0.835
cc_92 N_GND_c_27_p N_A_27_115#_M1021_g 0.00606474f $X=3.305 $Y=0.152 $X2=3.175
+ $Y2=0.835
cc_93 N_GND_c_28_p N_A_27_115#_M1021_g 0.00308284f $X=3.39 $Y=0.74 $X2=3.175
+ $Y2=0.835
cc_94 N_GND_c_3_p N_A_27_115#_M1021_g 0.00468827f $X=7.815 $Y=0.19 $X2=3.175
+ $Y2=0.835
cc_95 N_GND_M1012_b N_A_27_115#_c_848_n 0.0241659f $X=-0.055 $Y=0 $X2=3.53
+ $Y2=1.37
cc_96 N_GND_c_28_p N_A_27_115#_c_848_n 9.93645e-19 $X=3.39 $Y=0.74 $X2=3.53
+ $Y2=1.37
cc_97 N_GND_M1012_b N_A_27_115#_c_850_n 0.0105855f $X=-0.055 $Y=0 $X2=3.25
+ $Y2=1.37
cc_98 N_GND_M1012_b N_A_27_115#_c_851_n 0.0232417f $X=-0.055 $Y=0 $X2=3.53
+ $Y2=2.285
cc_99 N_GND_M1012_b N_A_27_115#_c_852_n 0.0105265f $X=-0.055 $Y=0 $X2=3.25
+ $Y2=2.285
cc_100 N_GND_M1012_b N_A_27_115#_M1013_g 0.0171936f $X=-0.055 $Y=0 $X2=3.605
+ $Y2=0.835
cc_101 N_GND_c_28_p N_A_27_115#_M1013_g 0.00308284f $X=3.39 $Y=0.74 $X2=3.605
+ $Y2=0.835
cc_102 N_GND_c_29_p N_A_27_115#_M1013_g 0.00606474f $X=5.055 $Y=0.152 $X2=3.605
+ $Y2=0.835
cc_103 N_GND_c_3_p N_A_27_115#_M1013_g 0.00468827f $X=7.815 $Y=0.19 $X2=3.605
+ $Y2=0.835
cc_104 N_GND_M1012_b N_A_27_115#_c_857_n 0.0010023f $X=-0.055 $Y=0 $X2=0.605
+ $Y2=0.91
cc_105 N_GND_c_2_p N_A_27_115#_c_857_n 0.00681706f $X=0.965 $Y=0.152 $X2=0.605
+ $Y2=0.91
cc_106 N_GND_c_3_p N_A_27_115#_c_857_n 0.00992214f $X=7.815 $Y=0.19 $X2=0.605
+ $Y2=0.91
cc_107 N_GND_M1012_b N_A_27_115#_c_860_n 0.0144521f $X=-0.055 $Y=0 $X2=0.69
+ $Y2=1.905
cc_108 N_GND_M1012_b N_A_27_115#_c_861_n 0.00871176f $X=-0.055 $Y=0 $X2=3.345
+ $Y2=2.285
cc_109 N_GND_M1012_b N_A_27_115#_c_862_n 0.00471684f $X=-0.055 $Y=0 $X2=0.26
+ $Y2=0.74
cc_110 N_GND_c_2_p N_A_27_115#_c_862_n 0.00710526f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_111 N_GND_c_3_p N_A_27_115#_c_862_n 0.00469007f $X=7.815 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_112 N_GND_M1012_b N_A_27_115#_c_865_n 0.0022123f $X=-0.055 $Y=0 $X2=3.345
+ $Y2=1.37
cc_113 N_GND_c_28_p N_A_27_115#_c_865_n 0.0044459f $X=3.39 $Y=0.74 $X2=3.345
+ $Y2=1.37
cc_114 N_GND_M1012_b N_A_27_115#_c_867_n 0.00267544f $X=-0.055 $Y=0 $X2=0.69
+ $Y2=1.79
cc_115 N_GND_M1012_b N_A_27_115#_c_868_n 0.0342377f $X=-0.055 $Y=0 $X2=3.11
+ $Y2=1.37
cc_116 N_GND_M1012_b N_A_27_115#_c_869_n 6.95759e-19 $X=-0.055 $Y=0 $X2=0.775
+ $Y2=1.37
cc_117 N_GND_M1012_b N_A_27_115#_c_870_n 0.00409378f $X=-0.055 $Y=0 $X2=0.69
+ $Y2=1.905
cc_118 N_GND_M1012_b N_A_428_89#_c_984_n 0.0173059f $X=-0.055 $Y=0 $X2=2.215
+ $Y2=1.205
cc_119 N_GND_c_27_p N_A_428_89#_c_984_n 0.00606474f $X=3.305 $Y=0.152 $X2=2.215
+ $Y2=1.205
cc_120 N_GND_c_3_p N_A_428_89#_c_984_n 0.00468827f $X=7.815 $Y=0.19 $X2=2.215
+ $Y2=1.205
cc_121 N_GND_M1012_b N_A_428_89#_c_987_n 0.0203057f $X=-0.055 $Y=0 $X2=2.335
+ $Y2=1.745
cc_122 N_GND_M1012_b N_A_428_89#_c_988_n 0.0207095f $X=-0.055 $Y=0 $X2=2.74
+ $Y2=1.82
cc_123 N_GND_M1012_b N_A_428_89#_c_989_n 0.00755029f $X=-0.055 $Y=0 $X2=2.41
+ $Y2=1.82
cc_124 N_GND_M1012_b N_A_428_89#_M1015_g 0.032457f $X=-0.055 $Y=0 $X2=2.815
+ $Y2=3.235
cc_125 N_GND_M1012_b N_A_428_89#_c_991_n 0.0559794f $X=-0.055 $Y=0 $X2=3.89
+ $Y2=1.82
cc_126 N_GND_M1012_b N_A_428_89#_M1022_g 0.0313037f $X=-0.055 $Y=0 $X2=3.965
+ $Y2=3.235
cc_127 N_GND_M1012_b N_A_428_89#_c_993_n 0.021099f $X=-0.055 $Y=0 $X2=4.37
+ $Y2=1.825
cc_128 N_GND_M1012_b N_A_428_89#_M1002_g 0.0348938f $X=-0.055 $Y=0 $X2=4.565
+ $Y2=0.835
cc_129 N_GND_c_29_p N_A_428_89#_M1002_g 0.00606474f $X=5.055 $Y=0.152 $X2=4.565
+ $Y2=0.835
cc_130 N_GND_c_3_p N_A_428_89#_M1002_g 0.00468827f $X=7.815 $Y=0.19 $X2=4.565
+ $Y2=0.835
cc_131 N_GND_M1012_b N_A_428_89#_c_997_n 0.0141736f $X=-0.055 $Y=0 $X2=2.335
+ $Y2=1.28
cc_132 N_GND_M1012_b N_A_428_89#_c_998_n 0.00426512f $X=-0.055 $Y=0 $X2=2.815
+ $Y2=1.82
cc_133 N_GND_M1012_b N_A_428_89#_c_999_n 0.00467948f $X=-0.055 $Y=0 $X2=3.965
+ $Y2=1.825
cc_134 N_GND_M1012_b N_A_428_89#_c_1000_n 0.0269513f $X=-0.055 $Y=0 $X2=4.505
+ $Y2=1.74
cc_135 N_GND_M1012_b N_A_428_89#_c_1001_n 0.00260727f $X=-0.055 $Y=0 $X2=4.505
+ $Y2=1.74
cc_136 N_GND_M1012_b N_A_428_89#_c_1002_n 0.0147565f $X=-0.055 $Y=0 $X2=5.57
+ $Y2=0.755
cc_137 N_GND_c_30_p N_A_428_89#_c_1002_n 4.65312e-19 $X=5.14 $Y=0.755 $X2=5.57
+ $Y2=0.755
cc_138 N_GND_c_6_p N_A_428_89#_c_1002_n 0.00747016f $X=6.795 $Y=0.152 $X2=5.57
+ $Y2=0.755
cc_139 N_GND_c_3_p N_A_428_89#_c_1002_n 0.00476261f $X=7.815 $Y=0.19 $X2=5.57
+ $Y2=0.755
cc_140 N_GND_M1012_b N_A_428_89#_c_1006_n 0.0117092f $X=-0.055 $Y=0 $X2=5.845
+ $Y2=2.62
cc_141 N_GND_M1012_b N_A_428_89#_c_1007_n 0.0097904f $X=-0.055 $Y=0 $X2=5.57
+ $Y2=1.755
cc_142 N_GND_M1012_b N_A_428_89#_c_1008_n 0.00759032f $X=-0.055 $Y=0 $X2=5.405
+ $Y2=1.74
cc_143 N_GND_M1012_b N_A_428_89#_c_1009_n 9.17297e-19 $X=-0.055 $Y=0 $X2=4.65
+ $Y2=1.74
cc_144 N_GND_M1012_b N_A_428_89#_c_1010_n 0.00142162f $X=-0.055 $Y=0 $X2=5.52
+ $Y2=1.74
cc_145 N_GND_M1012_b N_A_970_89#_M1006_g 0.0321276f $X=-0.055 $Y=0 $X2=4.925
+ $Y2=0.835
cc_146 N_GND_c_29_p N_A_970_89#_M1006_g 0.00606474f $X=5.055 $Y=0.152 $X2=4.925
+ $Y2=0.835
cc_147 N_GND_c_30_p N_A_970_89#_M1006_g 0.00315235f $X=5.14 $Y=0.755 $X2=4.925
+ $Y2=0.835
cc_148 N_GND_c_3_p N_A_970_89#_M1006_g 0.00468827f $X=7.815 $Y=0.19 $X2=4.925
+ $Y2=0.835
cc_149 N_GND_M1012_b N_A_970_89#_M1026_g 0.0300755f $X=-0.055 $Y=0 $X2=4.925
+ $Y2=3.235
cc_150 N_GND_M1012_b N_A_970_89#_c_1185_n 0.0259647f $X=-0.055 $Y=0 $X2=4.985
+ $Y2=1.71
cc_151 N_GND_c_30_p N_A_970_89#_c_1185_n 0.00109087f $X=5.14 $Y=0.755 $X2=4.985
+ $Y2=1.71
cc_152 N_GND_M1012_b N_A_970_89#_c_1187_n 0.0292185f $X=-0.055 $Y=0 $X2=7.57
+ $Y2=1.71
cc_153 N_GND_M1012_b N_A_970_89#_c_1188_n 0.0147409f $X=-0.055 $Y=0 $X2=7.572
+ $Y2=1.545
cc_154 N_GND_M1012_b N_A_970_89#_c_1189_n 0.0169275f $X=-0.055 $Y=0 $X2=7.66
+ $Y2=1.17
cc_155 N_GND_c_7_p N_A_970_89#_c_1189_n 0.00344579f $X=6.88 $Y=0.74 $X2=7.66
+ $Y2=1.17
cc_156 N_GND_c_33_p N_A_970_89#_c_1189_n 0.00606474f $X=7.815 $Y=0.152 $X2=7.66
+ $Y2=1.17
cc_157 N_GND_c_157_p N_A_970_89#_c_1189_n 0.00308284f $X=7.9 $Y=0.74 $X2=7.66
+ $Y2=1.17
cc_158 N_GND_c_3_p N_A_970_89#_c_1189_n 0.00468827f $X=7.815 $Y=0.19 $X2=7.66
+ $Y2=1.17
cc_159 N_GND_M1012_b N_A_970_89#_c_1194_n 0.0136411f $X=-0.055 $Y=0 $X2=7.66
+ $Y2=1.32
cc_160 N_GND_M1012_b N_A_970_89#_c_1195_n 0.0365245f $X=-0.055 $Y=0 $X2=7.66
+ $Y2=2.375
cc_161 N_GND_M1012_b N_A_970_89#_c_1196_n 0.00495925f $X=-0.055 $Y=0 $X2=7.66
+ $Y2=2.525
cc_162 N_GND_M1012_b N_A_970_89#_c_1197_n 0.00491423f $X=-0.055 $Y=0 $X2=4.985
+ $Y2=1.71
cc_163 N_GND_M1012_b N_A_970_89#_c_1198_n 9.87353e-19 $X=-0.055 $Y=0 $X2=6.435
+ $Y2=0.91
cc_164 N_GND_c_6_p N_A_970_89#_c_1198_n 0.00658268f $X=6.795 $Y=0.152 $X2=6.435
+ $Y2=0.91
cc_165 N_GND_c_3_p N_A_970_89#_c_1198_n 0.00992214f $X=7.815 $Y=0.19 $X2=6.435
+ $Y2=0.91
cc_166 N_GND_M1012_b N_A_970_89#_c_1201_n 0.00666412f $X=-0.055 $Y=0 $X2=6.52
+ $Y2=1.625
cc_167 N_GND_M1012_b N_A_970_89#_c_1202_n 0.0133983f $X=-0.055 $Y=0 $X2=6.52
+ $Y2=3.615
cc_168 N_GND_M1012_b N_A_970_89#_c_1203_n 0.0176905f $X=-0.055 $Y=0 $X2=7.57
+ $Y2=1.71
cc_169 N_GND_M1012_b N_A_970_89#_c_1204_n 0.00292206f $X=-0.055 $Y=0 $X2=6.09
+ $Y2=0.74
cc_170 N_GND_c_6_p N_A_970_89#_c_1204_n 0.00732079f $X=6.795 $Y=0.152 $X2=6.09
+ $Y2=0.74
cc_171 N_GND_c_3_p N_A_970_89#_c_1204_n 0.00469007f $X=7.815 $Y=0.19 $X2=6.09
+ $Y2=0.74
cc_172 N_GND_M1012_b N_A_970_89#_c_1207_n 0.00194787f $X=-0.055 $Y=0 $X2=6.52
+ $Y2=1.71
cc_173 N_GND_M1012_b N_A_970_89#_c_1208_n 0.00282652f $X=-0.055 $Y=0 $X2=5.785
+ $Y2=2.48
cc_174 N_GND_M1012_b N_A_970_89#_c_1209_n 0.00123753f $X=-0.055 $Y=0 $X2=5.13
+ $Y2=2.48
cc_175 N_GND_M1012_b N_A_970_89#_c_1210_n 0.00597518f $X=-0.055 $Y=0 $X2=5.882
+ $Y2=2.39
cc_176 N_GND_M1012_b N_A_970_89#_c_1211_n 0.0505983f $X=-0.055 $Y=0 $X2=7.425
+ $Y2=1.71
cc_177 N_GND_M1012_b N_A_970_89#_c_1212_n 0.00133099f $X=-0.055 $Y=0 $X2=5.96
+ $Y2=1.71
cc_178 N_GND_M1012_b N_A_970_89#_c_1213_n 0.00173636f $X=-0.055 $Y=0 $X2=7.57
+ $Y2=1.71
cc_179 N_GND_M1012_b N_A_808_115#_M1004_g 0.0302349f $X=-0.055 $Y=0 $X2=6.305
+ $Y2=0.755
cc_180 N_GND_c_6_p N_A_808_115#_M1004_g 0.00454486f $X=6.795 $Y=0.152 $X2=6.305
+ $Y2=0.755
cc_181 N_GND_c_3_p N_A_808_115#_M1004_g 0.00468827f $X=7.815 $Y=0.19 $X2=6.305
+ $Y2=0.755
cc_182 N_GND_M1012_b N_A_808_115#_M1024_g 0.0548993f $X=-0.055 $Y=0 $X2=6.305
+ $Y2=3.445
cc_183 N_GND_M1012_b N_A_808_115#_c_1382_n 0.0439803f $X=-0.055 $Y=0 $X2=6.305
+ $Y2=1.37
cc_184 N_GND_M1012_b N_A_808_115#_c_1383_n 0.0111437f $X=-0.055 $Y=0 $X2=3.685
+ $Y2=1.37
cc_185 N_GND_M1012_b N_A_808_115#_c_1384_n 0.00915481f $X=-0.055 $Y=0 $X2=4.365
+ $Y2=1.37
cc_186 N_GND_M1012_b N_A_808_115#_c_1385_n 0.00162209f $X=-0.055 $Y=0 $X2=6.1
+ $Y2=1.37
cc_187 N_GND_M1012_b N_A_808_115#_c_1386_n 0.00312748f $X=-0.055 $Y=0 $X2=4.265
+ $Y2=0.755
cc_188 N_GND_c_29_p N_A_808_115#_c_1386_n 0.0150533f $X=5.055 $Y=0.152 $X2=4.265
+ $Y2=0.755
cc_189 N_GND_c_3_p N_A_808_115#_c_1386_n 0.00994746f $X=7.815 $Y=0.19 $X2=4.265
+ $Y2=0.755
cc_190 N_GND_M1012_b N_A_808_115#_c_1389_n 0.00267903f $X=-0.055 $Y=0 $X2=4.245
+ $Y2=1.37
cc_191 N_GND_M1012_b N_A_808_115#_c_1390_n 0.00201489f $X=-0.055 $Y=0 $X2=3.83
+ $Y2=1.37
cc_192 N_GND_M1012_b N_A_808_115#_c_1391_n 0.0123881f $X=-0.055 $Y=0 $X2=5.955
+ $Y2=1.37
cc_193 N_GND_c_30_p N_A_808_115#_c_1391_n 8.8332e-19 $X=5.14 $Y=0.755 $X2=5.955
+ $Y2=1.37
cc_194 N_GND_M1012_b N_A_808_115#_c_1393_n 0.0027147f $X=-0.055 $Y=0 $X2=4.48
+ $Y2=1.37
cc_195 N_GND_M1012_b N_A_808_115#_c_1394_n 6.75279e-19 $X=-0.055 $Y=0 $X2=6.1
+ $Y2=1.37
cc_196 N_GND_M1012_b N_QN_M1027_g 0.0561552f $X=-0.055 $Y=0 $X2=8.115 $Y2=0.835
cc_197 N_GND_c_157_p N_QN_M1027_g 0.00308284f $X=7.9 $Y=0.74 $X2=8.115 $Y2=0.835
cc_198 N_GND_c_3_p N_QN_M1027_g 0.00468827f $X=7.815 $Y=0.19 $X2=8.115 $Y2=0.835
cc_199 N_GND_M1012_b N_QN_M1019_g 0.0186095f $X=-0.055 $Y=0 $X2=8.115 $Y2=3.235
cc_200 N_GND_M1012_b N_QN_c_1527_n 0.0291912f $X=-0.055 $Y=0 $X2=8.055 $Y2=1.915
cc_201 N_GND_M1012_b N_QN_c_1528_n 0.00453751f $X=-0.055 $Y=0 $X2=7.47 $Y2=0.74
cc_202 N_GND_c_7_p N_QN_c_1528_n 0.0124968f $X=6.88 $Y=0.74 $X2=7.47 $Y2=0.74
cc_203 N_GND_c_33_p N_QN_c_1528_n 0.00757793f $X=7.815 $Y=0.152 $X2=7.47
+ $Y2=0.74
cc_204 N_GND_c_3_p N_QN_c_1528_n 0.00476261f $X=7.815 $Y=0.19 $X2=7.47 $Y2=0.74
cc_205 N_GND_M1012_b N_QN_c_1532_n 0.00138285f $X=-0.055 $Y=0 $X2=7.47 $Y2=2.48
cc_206 N_GND_M1012_b N_QN_c_1533_n 0.0134237f $X=-0.055 $Y=0 $X2=7.97 $Y2=1.37
cc_207 N_GND_c_157_p N_QN_c_1533_n 0.00779875f $X=7.9 $Y=0.74 $X2=7.97 $Y2=1.37
cc_208 N_GND_M1012_b N_QN_c_1535_n 0.0029714f $X=-0.055 $Y=0 $X2=7.555 $Y2=1.37
cc_209 N_GND_M1012_b N_QN_c_1536_n 0.0138424f $X=-0.055 $Y=0 $X2=7.97 $Y2=2.285
cc_210 N_GND_M1012_b N_QN_c_1537_n 0.00426693f $X=-0.055 $Y=0 $X2=7.555
+ $Y2=2.285
cc_211 N_GND_M1012_b N_QN_c_1538_n 0.0034889f $X=-0.055 $Y=0 $X2=8.055 $Y2=1.915
cc_212 N_GND_M1012_b QN 0.00291738f $X=-0.055 $Y=0 $X2=7.475 $Y2=2.48
cc_213 N_GND_M1012_b N_Q_c_1610_n 0.00880645f $X=-0.055 $Y=0 $X2=8.33 $Y2=0.74
cc_214 N_GND_c_3_p N_Q_c_1610_n 0.00467398f $X=7.815 $Y=0.19 $X2=8.33 $Y2=0.74
cc_215 N_GND_M1012_b N_Q_c_1612_n 0.0625704f $X=-0.055 $Y=0 $X2=8.445 $Y2=2.68
cc_216 N_GND_M1012_b N_Q_c_1613_n 0.0152652f $X=-0.055 $Y=0 $X2=8.445 $Y2=1.035
cc_217 N_VDD_M1009_b N_SN_M1009_g 0.0602812f $X=-0.055 $Y=2.815 $X2=0.475
+ $Y2=3.445
cc_218 N_VDD_c_218_p N_SN_M1009_g 0.00713292f $X=0.26 $Y=3.615 $X2=0.475
+ $Y2=3.445
cc_219 N_VDD_c_219_p N_SN_M1009_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475
+ $Y2=3.445
cc_220 N_VDD_c_220_p N_SN_M1009_g 0.00468827f $X=7.815 $Y=4.25 $X2=0.475
+ $Y2=3.445
cc_221 N_VDD_M1009_b N_SN_M1016_g 0.0498528f $X=-0.055 $Y=2.815 $X2=6.735
+ $Y2=3.445
cc_222 N_VDD_c_222_p N_SN_M1016_g 0.00606474f $X=6.865 $Y=4.287 $X2=6.735
+ $Y2=3.445
cc_223 N_VDD_c_223_p N_SN_M1016_g 0.00713292f $X=6.95 $Y=3.615 $X2=6.735
+ $Y2=3.445
cc_224 N_VDD_c_220_p N_SN_M1016_g 0.00468827f $X=7.815 $Y=4.25 $X2=6.735
+ $Y2=3.445
cc_225 N_VDD_M1009_b N_A_152_89#_M1020_g 0.0535193f $X=-0.055 $Y=2.815 $X2=0.905
+ $Y2=3.445
cc_226 N_VDD_c_219_p N_A_152_89#_M1020_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905
+ $Y2=3.445
cc_227 N_VDD_c_227_p N_A_152_89#_M1020_g 0.00713292f $X=1.12 $Y=3.615 $X2=0.905
+ $Y2=3.445
cc_228 N_VDD_c_228_p N_A_152_89#_M1020_g 0.00802793f $X=1.64 $Y=3.295 $X2=0.905
+ $Y2=3.445
cc_229 N_VDD_c_220_p N_A_152_89#_M1020_g 0.00468827f $X=7.815 $Y=4.25 $X2=0.905
+ $Y2=3.445
cc_230 N_VDD_M1009_b N_A_152_89#_c_485_n 0.00286294f $X=-0.055 $Y=2.815 $X2=1.03
+ $Y2=1.925
cc_231 N_VDD_M1007_s N_A_152_89#_c_501_n 0.0125004f $X=1.515 $Y=2.605 $X2=2.345
+ $Y2=2.705
cc_232 N_VDD_M1009_b N_A_152_89#_c_501_n 0.0269258f $X=-0.055 $Y=2.815 $X2=2.345
+ $Y2=2.705
cc_233 N_VDD_c_227_p N_A_152_89#_c_501_n 0.00302899f $X=1.12 $Y=3.615 $X2=2.345
+ $Y2=2.705
cc_234 N_VDD_c_228_p N_A_152_89#_c_501_n 0.00952036f $X=1.64 $Y=3.295 $X2=2.345
+ $Y2=2.705
cc_235 N_VDD_M1009_b N_A_152_89#_c_505_n 0.00352946f $X=-0.055 $Y=2.815
+ $X2=1.115 $Y2=2.705
cc_236 N_VDD_c_227_p N_A_152_89#_c_505_n 0.00296793f $X=1.12 $Y=3.615 $X2=1.115
+ $Y2=2.705
cc_237 N_VDD_M1009_b N_A_152_89#_c_507_n 0.00313975f $X=-0.055 $Y=2.815
+ $X2=2.515 $Y2=2.955
cc_238 N_VDD_c_238_p N_A_152_89#_c_507_n 0.0149461f $X=3.305 $Y=4.287 $X2=2.515
+ $Y2=2.955
cc_239 N_VDD_c_220_p N_A_152_89#_c_507_n 0.00958198f $X=7.815 $Y=4.25 $X2=2.515
+ $Y2=2.955
cc_240 N_VDD_M1009_b N_D_M1007_g 0.0222869f $X=-0.055 $Y=2.815 $X2=1.855
+ $Y2=3.235
cc_241 N_VDD_c_228_p N_D_M1007_g 0.00636672f $X=1.64 $Y=3.295 $X2=1.855
+ $Y2=3.235
cc_242 N_VDD_c_238_p N_D_M1007_g 0.00606474f $X=3.305 $Y=4.287 $X2=1.855
+ $Y2=3.235
cc_243 N_VDD_c_220_p N_D_M1007_g 0.00468827f $X=7.815 $Y=4.25 $X2=1.855
+ $Y2=3.235
cc_244 N_VDD_M1009_b N_CK_M1011_g 0.020128f $X=-0.055 $Y=2.815 $X2=2.215
+ $Y2=3.235
cc_245 N_VDD_c_238_p N_CK_M1011_g 0.00606474f $X=3.305 $Y=4.287 $X2=2.215
+ $Y2=3.235
cc_246 N_VDD_c_220_p N_CK_M1011_g 0.00468827f $X=7.815 $Y=4.25 $X2=2.215
+ $Y2=3.235
cc_247 N_VDD_M1009_b N_CK_M1028_g 0.0201163f $X=-0.055 $Y=2.815 $X2=4.565
+ $Y2=3.235
cc_248 N_VDD_c_248_p N_CK_M1028_g 0.00606474f $X=5.055 $Y=4.287 $X2=4.565
+ $Y2=3.235
cc_249 N_VDD_c_220_p N_CK_M1028_g 0.00468827f $X=7.815 $Y=4.25 $X2=4.565
+ $Y2=3.235
cc_250 N_VDD_M1009_b N_CK_c_611_n 0.007968f $X=-0.055 $Y=2.815 $X2=5.355
+ $Y2=2.45
cc_251 N_VDD_M1009_b N_CK_M1017_g 0.0218804f $X=-0.055 $Y=2.815 $X2=5.355
+ $Y2=3.235
cc_252 N_VDD_c_252_p N_CK_M1017_g 0.00409291f $X=5.14 $Y=3.21 $X2=5.355
+ $Y2=3.235
cc_253 N_VDD_c_253_p N_CK_M1017_g 0.00606474f $X=6.005 $Y=4.287 $X2=5.355
+ $Y2=3.235
cc_254 N_VDD_c_254_p N_CK_M1017_g 0.00394336f $X=6.09 $Y=3.615 $X2=5.355
+ $Y2=3.235
cc_255 N_VDD_c_220_p N_CK_M1017_g 0.00468827f $X=7.815 $Y=4.25 $X2=5.355
+ $Y2=3.235
cc_256 N_VDD_M1009_b N_CK_c_613_n 0.00487135f $X=-0.055 $Y=2.815 $X2=2.275
+ $Y2=2.285
cc_257 N_VDD_M1009_b N_CK_c_622_n 0.00486793f $X=-0.055 $Y=2.815 $X2=4.505
+ $Y2=2.285
cc_258 N_VDD_M1009_b N_CK_c_633_n 0.0010436f $X=-0.055 $Y=2.815 $X2=5.5 $Y2=2.11
cc_259 N_VDD_M1009_b N_CK_c_634_n 6.42499e-19 $X=-0.055 $Y=2.815 $X2=2.275
+ $Y2=2.11
cc_260 N_VDD_M1009_b N_CK_c_635_n 0.0022456f $X=-0.055 $Y=2.815 $X2=4.505
+ $Y2=2.11
cc_261 N_VDD_M1009_b N_A_27_115#_M1014_g 0.0192219f $X=-0.055 $Y=2.815 $X2=3.175
+ $Y2=3.235
cc_262 N_VDD_c_238_p N_A_27_115#_M1014_g 0.00606474f $X=3.305 $Y=4.287 $X2=3.175
+ $Y2=3.235
cc_263 N_VDD_c_263_p N_A_27_115#_M1014_g 0.00337744f $X=3.39 $Y=3.295 $X2=3.175
+ $Y2=3.235
cc_264 N_VDD_c_220_p N_A_27_115#_M1014_g 0.00468827f $X=7.815 $Y=4.25 $X2=3.175
+ $Y2=3.235
cc_265 N_VDD_c_263_p N_A_27_115#_c_851_n 8.24975e-19 $X=3.39 $Y=3.295 $X2=3.53
+ $Y2=2.285
cc_266 N_VDD_M1009_b N_A_27_115#_M1005_g 0.0181098f $X=-0.055 $Y=2.815 $X2=3.605
+ $Y2=3.235
cc_267 N_VDD_c_263_p N_A_27_115#_M1005_g 0.00337744f $X=3.39 $Y=3.295 $X2=3.605
+ $Y2=3.235
cc_268 N_VDD_c_248_p N_A_27_115#_M1005_g 0.00606474f $X=5.055 $Y=4.287 $X2=3.605
+ $Y2=3.235
cc_269 N_VDD_c_220_p N_A_27_115#_M1005_g 0.00468827f $X=7.815 $Y=4.25 $X2=3.605
+ $Y2=3.235
cc_270 N_VDD_M1009_b N_A_27_115#_c_860_n 0.0147746f $X=-0.055 $Y=2.815 $X2=0.69
+ $Y2=1.905
cc_271 N_VDD_c_219_p N_A_27_115#_c_860_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69
+ $Y2=1.905
cc_272 N_VDD_c_220_p N_A_27_115#_c_860_n 0.00475776f $X=7.815 $Y=4.25 $X2=0.69
+ $Y2=1.905
cc_273 N_VDD_M1009_b N_A_27_115#_c_861_n 0.00424346f $X=-0.055 $Y=2.815
+ $X2=3.345 $Y2=2.285
cc_274 N_VDD_c_263_p N_A_27_115#_c_861_n 0.004428f $X=3.39 $Y=3.295 $X2=3.345
+ $Y2=2.285
cc_275 N_VDD_M1009_b N_A_428_89#_M1015_g 0.0215131f $X=-0.055 $Y=2.815 $X2=2.815
+ $Y2=3.235
cc_276 N_VDD_c_238_p N_A_428_89#_M1015_g 0.00606474f $X=3.305 $Y=4.287 $X2=2.815
+ $Y2=3.235
cc_277 N_VDD_c_220_p N_A_428_89#_M1015_g 0.00468827f $X=7.815 $Y=4.25 $X2=2.815
+ $Y2=3.235
cc_278 N_VDD_M1009_b N_A_428_89#_M1022_g 0.0214821f $X=-0.055 $Y=2.815 $X2=3.965
+ $Y2=3.235
cc_279 N_VDD_c_248_p N_A_428_89#_M1022_g 0.00606474f $X=5.055 $Y=4.287 $X2=3.965
+ $Y2=3.235
cc_280 N_VDD_c_220_p N_A_428_89#_M1022_g 0.00468827f $X=7.815 $Y=4.25 $X2=3.965
+ $Y2=3.235
cc_281 N_VDD_M1009_b N_A_428_89#_c_1017_n 0.00156053f $X=-0.055 $Y=2.815
+ $X2=5.57 $Y2=2.955
cc_282 N_VDD_c_253_p N_A_428_89#_c_1017_n 0.00747016f $X=6.005 $Y=4.287 $X2=5.57
+ $Y2=2.955
cc_283 N_VDD_c_254_p N_A_428_89#_c_1017_n 0.0213592f $X=6.09 $Y=3.615 $X2=5.57
+ $Y2=2.955
cc_284 N_VDD_c_220_p N_A_428_89#_c_1017_n 0.00476261f $X=7.815 $Y=4.25 $X2=5.57
+ $Y2=2.955
cc_285 N_VDD_M1009_b N_A_428_89#_c_1006_n 0.00552543f $X=-0.055 $Y=2.815
+ $X2=5.845 $Y2=2.62
cc_286 N_VDD_M1009_b N_A_428_89#_c_1022_n 0.0123356f $X=-0.055 $Y=2.815
+ $X2=5.845 $Y2=2.705
cc_287 N_VDD_M1009_b N_A_970_89#_M1026_g 0.0178558f $X=-0.055 $Y=2.815 $X2=4.925
+ $Y2=3.235
cc_288 N_VDD_c_248_p N_A_970_89#_M1026_g 0.00606474f $X=5.055 $Y=4.287 $X2=4.925
+ $Y2=3.235
cc_289 N_VDD_c_252_p N_A_970_89#_M1026_g 0.00409291f $X=5.14 $Y=3.21 $X2=4.925
+ $Y2=3.235
cc_290 N_VDD_c_220_p N_A_970_89#_M1026_g 0.00468827f $X=7.815 $Y=4.25 $X2=4.925
+ $Y2=3.235
cc_291 N_VDD_M1009_b N_A_970_89#_c_1196_n 0.0266934f $X=-0.055 $Y=2.815 $X2=7.66
+ $Y2=2.525
cc_292 N_VDD_c_223_p N_A_970_89#_c_1196_n 0.00394336f $X=6.95 $Y=3.615 $X2=7.66
+ $Y2=2.525
cc_293 N_VDD_c_293_p N_A_970_89#_c_1196_n 0.00606474f $X=7.815 $Y=4.287 $X2=7.66
+ $Y2=2.525
cc_294 N_VDD_c_294_p N_A_970_89#_c_1196_n 0.00480838f $X=7.9 $Y=3.265 $X2=7.66
+ $Y2=2.525
cc_295 N_VDD_c_220_p N_A_970_89#_c_1196_n 0.00468827f $X=7.815 $Y=4.25 $X2=7.66
+ $Y2=2.525
cc_296 N_VDD_M1009_b N_A_970_89#_c_1197_n 0.00242843f $X=-0.055 $Y=2.815
+ $X2=4.985 $Y2=1.71
cc_297 N_VDD_c_252_p N_A_970_89#_c_1197_n 4.62798e-19 $X=5.14 $Y=3.21 $X2=4.985
+ $Y2=1.71
cc_298 N_VDD_M1009_b N_A_970_89#_c_1202_n 0.0151745f $X=-0.055 $Y=2.815 $X2=6.52
+ $Y2=3.615
cc_299 N_VDD_c_222_p N_A_970_89#_c_1202_n 0.00734006f $X=6.865 $Y=4.287 $X2=6.52
+ $Y2=3.615
cc_300 N_VDD_c_220_p N_A_970_89#_c_1202_n 0.00475776f $X=7.815 $Y=4.25 $X2=6.52
+ $Y2=3.615
cc_301 N_VDD_M1009_b N_A_970_89#_c_1208_n 0.00919639f $X=-0.055 $Y=2.815
+ $X2=5.785 $Y2=2.48
cc_302 N_VDD_c_252_p N_A_970_89#_c_1208_n 0.00425473f $X=5.14 $Y=3.21 $X2=5.785
+ $Y2=2.48
cc_303 N_VDD_M1009_b N_A_970_89#_c_1209_n 0.00604093f $X=-0.055 $Y=2.815
+ $X2=5.13 $Y2=2.48
cc_304 N_VDD_c_252_p N_A_970_89#_c_1209_n 0.003295f $X=5.14 $Y=3.21 $X2=5.13
+ $Y2=2.48
cc_305 N_VDD_M1009_b N_A_808_115#_M1024_g 0.047909f $X=-0.055 $Y=2.815 $X2=6.305
+ $Y2=3.445
cc_306 N_VDD_c_254_p N_A_808_115#_M1024_g 0.00713292f $X=6.09 $Y=3.615 $X2=6.305
+ $Y2=3.445
cc_307 N_VDD_c_222_p N_A_808_115#_M1024_g 0.00606474f $X=6.865 $Y=4.287
+ $X2=6.305 $Y2=3.445
cc_308 N_VDD_c_220_p N_A_808_115#_M1024_g 0.00468827f $X=7.815 $Y=4.25 $X2=6.305
+ $Y2=3.445
cc_309 N_VDD_M1009_b N_A_808_115#_c_1383_n 0.00168314f $X=-0.055 $Y=2.815
+ $X2=3.685 $Y2=1.37
cc_310 N_VDD_M1009_b N_A_808_115#_c_1400_n 0.00313975f $X=-0.055 $Y=2.815
+ $X2=4.265 $Y2=3.295
cc_311 N_VDD_c_248_p N_A_808_115#_c_1400_n 0.014959f $X=5.055 $Y=4.287 $X2=4.265
+ $Y2=3.295
cc_312 N_VDD_c_220_p N_A_808_115#_c_1400_n 0.00958198f $X=7.815 $Y=4.25
+ $X2=4.265 $Y2=3.295
cc_313 N_VDD_M1009_b N_QN_M1019_g 0.0248218f $X=-0.055 $Y=2.815 $X2=8.115
+ $Y2=3.235
cc_314 N_VDD_c_294_p N_QN_M1019_g 0.00480838f $X=7.9 $Y=3.265 $X2=8.115
+ $Y2=3.235
cc_315 N_VDD_c_315_p N_QN_M1019_g 0.00606474f $X=7.815 $Y=4.25 $X2=8.115
+ $Y2=3.235
cc_316 N_VDD_c_220_p N_QN_M1019_g 0.00468827f $X=7.815 $Y=4.25 $X2=8.115
+ $Y2=3.235
cc_317 N_VDD_M1009_b N_QN_c_1532_n 0.00648064f $X=-0.055 $Y=2.815 $X2=7.47
+ $Y2=2.48
cc_318 N_VDD_c_223_p N_QN_c_1532_n 0.0213592f $X=6.95 $Y=3.615 $X2=7.47 $Y2=2.48
cc_319 N_VDD_c_293_p N_QN_c_1532_n 0.00757793f $X=7.815 $Y=4.287 $X2=7.47
+ $Y2=2.48
cc_320 N_VDD_c_220_p N_QN_c_1532_n 0.00476261f $X=7.815 $Y=4.25 $X2=7.47
+ $Y2=2.48
cc_321 N_VDD_c_294_p N_QN_c_1536_n 0.00818856f $X=7.9 $Y=3.265 $X2=7.97
+ $Y2=2.285
cc_322 N_VDD_M1009_b QN 0.0108749f $X=-0.055 $Y=2.815 $X2=7.475 $Y2=2.48
cc_323 N_VDD_M1009_b N_Q_c_1614_n 0.00156053f $X=-0.055 $Y=2.815 $X2=8.33
+ $Y2=3.265
cc_324 N_VDD_c_315_p N_Q_c_1614_n 0.00757793f $X=7.815 $Y=4.25 $X2=8.33
+ $Y2=3.265
cc_325 N_VDD_c_220_p N_Q_c_1614_n 0.00476261f $X=7.815 $Y=4.25 $X2=8.33
+ $Y2=3.265
cc_326 N_VDD_M1009_b N_Q_c_1612_n 0.0117744f $X=-0.055 $Y=2.815 $X2=8.445
+ $Y2=2.68
cc_327 N_VDD_M1009_b N_Q_c_1618_n 0.0093035f $X=-0.055 $Y=2.815 $X2=8.33
+ $Y2=2.807
cc_328 N_VDD_M1009_b Q 0.00503768f $X=-0.055 $Y=2.815 $X2=8.325 $Y2=2.85
cc_329 N_VDD_c_294_p Q 0.00675808f $X=7.9 $Y=3.265 $X2=8.325 $Y2=2.85
cc_330 N_SN_c_346_n N_A_152_89#_M1023_d 0.00331296f $X=1.405 $Y=0.985 $X2=2.29
+ $Y2=0.575
cc_331 N_SN_M1012_g N_A_152_89#_M1000_g 0.0505158f $X=0.475 $Y=0.755 $X2=0.835
+ $Y2=0.755
cc_332 N_SN_c_342_n N_A_152_89#_M1000_g 3.99631e-19 $X=0.32 $Y=1.47 $X2=0.835
+ $Y2=0.755
cc_333 N_SN_c_346_n N_A_152_89#_M1000_g 0.00552757f $X=1.405 $Y=0.985 $X2=0.835
+ $Y2=0.755
cc_334 N_SN_M1009_g N_A_152_89#_M1020_g 0.0538406f $X=0.475 $Y=3.445 $X2=0.905
+ $Y2=3.445
cc_335 N_SN_c_339_n N_A_152_89#_c_484_n 0.0505158f $X=0.32 $Y=1.47 $X2=1.03
+ $Y2=1.925
cc_336 N_SN_c_346_n N_A_152_89#_c_486_n 0.0286687f $X=1.405 $Y=0.985 $X2=2.33
+ $Y2=1.285
cc_337 N_SN_c_346_n N_A_152_89#_c_489_n 0.00229619f $X=1.405 $Y=0.985 $X2=1.115
+ $Y2=1.285
cc_338 N_SN_c_346_n N_A_152_89#_c_491_n 0.0132104f $X=1.405 $Y=0.985 $X2=2.415
+ $Y2=1.2
cc_339 N_SN_c_346_n N_A_152_89#_c_492_n 0.0130964f $X=1.405 $Y=0.985 $X2=2.415
+ $Y2=0.755
cc_340 N_SN_c_346_n N_D_M1001_g 0.00615654f $X=1.405 $Y=0.985 $X2=1.855
+ $Y2=0.835
cc_341 N_SN_c_346_n N_CK_c_614_n 7.97906e-19 $X=1.405 $Y=0.985 $X2=2.755
+ $Y2=1.37
cc_342 N_SN_c_346_n N_CK_c_615_n 0.00594264f $X=1.405 $Y=0.985 $X2=2.755
+ $Y2=1.205
cc_343 N_SN_c_346_n N_CK_c_618_n 7.97906e-19 $X=1.405 $Y=0.985 $X2=4.025
+ $Y2=1.37
cc_344 N_SN_c_346_n N_CK_c_619_n 0.00589873f $X=1.405 $Y=0.985 $X2=4.025
+ $Y2=1.205
cc_345 N_SN_c_346_n N_CK_c_623_n 0.00650745f $X=1.405 $Y=0.985 $X2=5.382
+ $Y2=1.205
cc_346 N_SN_c_346_n N_CK_c_627_n 0.00106638f $X=1.405 $Y=0.985 $X2=5.382
+ $Y2=1.355
cc_347 N_SN_c_346_n N_CK_c_629_n 0.00482442f $X=1.405 $Y=0.985 $X2=2.755
+ $Y2=1.37
cc_348 N_SN_c_346_n N_CK_c_630_n 0.0048224f $X=1.405 $Y=0.985 $X2=4.025 $Y2=1.37
cc_349 N_SN_c_346_n N_A_27_115#_M1021_g 0.00567f $X=1.405 $Y=0.985 $X2=3.175
+ $Y2=0.835
cc_350 N_SN_c_346_n N_A_27_115#_c_848_n 2.33608e-19 $X=1.405 $Y=0.985 $X2=3.53
+ $Y2=1.37
cc_351 N_SN_c_346_n N_A_27_115#_M1013_g 0.00592874f $X=1.405 $Y=0.985 $X2=3.605
+ $Y2=0.835
cc_352 N_SN_M1012_g N_A_27_115#_c_857_n 0.0113757f $X=0.475 $Y=0.755 $X2=0.605
+ $Y2=0.91
cc_353 N_SN_c_339_n N_A_27_115#_c_857_n 2.9588e-19 $X=0.32 $Y=1.47 $X2=0.605
+ $Y2=0.91
cc_354 N_SN_c_342_n N_A_27_115#_c_857_n 0.0021045f $X=0.32 $Y=1.47 $X2=0.605
+ $Y2=0.91
cc_355 N_SN_c_346_n N_A_27_115#_c_857_n 0.0152444f $X=1.405 $Y=0.985 $X2=0.605
+ $Y2=0.91
cc_356 N_SN_c_363_n N_A_27_115#_c_857_n 0.00261497f $X=0.405 $Y=0.985 $X2=0.605
+ $Y2=0.91
cc_357 SN N_A_27_115#_c_857_n 7.12685e-19 $X=0.32 $Y=1.535 $X2=0.605 $Y2=0.91
cc_358 N_SN_M1012_g N_A_27_115#_c_860_n 0.0424099f $X=0.475 $Y=0.755 $X2=0.69
+ $Y2=1.905
cc_359 N_SN_c_342_n N_A_27_115#_c_860_n 0.018845f $X=0.32 $Y=1.47 $X2=0.69
+ $Y2=1.905
cc_360 N_SN_c_345_n N_A_27_115#_c_860_n 0.00994822f $X=0.32 $Y=1.415 $X2=0.69
+ $Y2=1.905
cc_361 N_SN_c_346_n N_A_27_115#_c_860_n 0.0074124f $X=1.405 $Y=0.985 $X2=0.69
+ $Y2=1.905
cc_362 SN N_A_27_115#_c_860_n 8.35233e-19 $X=0.32 $Y=1.535 $X2=0.69 $Y2=1.905
cc_363 N_SN_M1012_g N_A_27_115#_c_862_n 5.28354e-19 $X=0.475 $Y=0.755 $X2=0.26
+ $Y2=0.74
cc_364 N_SN_c_339_n N_A_27_115#_c_862_n 0.00243073f $X=0.32 $Y=1.47 $X2=0.26
+ $Y2=0.74
cc_365 N_SN_c_342_n N_A_27_115#_c_862_n 0.00395258f $X=0.32 $Y=1.47 $X2=0.26
+ $Y2=0.74
cc_366 N_SN_c_363_n N_A_27_115#_c_862_n 0.0089299f $X=0.405 $Y=0.985 $X2=0.26
+ $Y2=0.74
cc_367 SN N_A_27_115#_c_862_n 0.00224014f $X=0.32 $Y=1.535 $X2=0.26 $Y2=0.74
cc_368 N_SN_c_346_n N_A_27_115#_c_865_n 0.00463957f $X=1.405 $Y=0.985 $X2=3.345
+ $Y2=1.37
cc_369 N_SN_c_339_n N_A_27_115#_c_867_n 0.00179417f $X=0.32 $Y=1.47 $X2=0.69
+ $Y2=1.79
cc_370 N_SN_c_346_n N_A_27_115#_c_868_n 0.128323f $X=1.405 $Y=0.985 $X2=3.11
+ $Y2=1.37
cc_371 N_SN_M1012_g N_A_27_115#_c_869_n 0.00179417f $X=0.475 $Y=0.755 $X2=0.775
+ $Y2=1.37
cc_372 N_SN_c_342_n N_A_27_115#_c_869_n 0.00153176f $X=0.32 $Y=1.47 $X2=0.775
+ $Y2=1.37
cc_373 N_SN_c_345_n N_A_27_115#_c_869_n 0.0117425f $X=0.32 $Y=1.415 $X2=0.775
+ $Y2=1.37
cc_374 N_SN_c_346_n N_A_27_115#_c_869_n 0.0596473f $X=1.405 $Y=0.985 $X2=0.775
+ $Y2=1.37
cc_375 SN N_A_27_115#_c_869_n 0.0241465f $X=0.32 $Y=1.535 $X2=0.775 $Y2=1.37
cc_376 N_SN_M1009_g N_A_27_115#_c_870_n 0.0103038f $X=0.475 $Y=3.445 $X2=0.69
+ $Y2=1.905
cc_377 N_SN_c_346_n N_A_27_115#_c_913_n 0.0240989f $X=1.405 $Y=0.985 $X2=3.255
+ $Y2=1.37
cc_378 N_SN_c_346_n N_A_428_89#_M1003_d 0.00202099f $X=1.405 $Y=0.985 $X2=5.43
+ $Y2=0.575
cc_379 N_SN_c_346_n N_A_428_89#_c_984_n 0.00557192f $X=1.405 $Y=0.985 $X2=2.215
+ $Y2=1.205
cc_380 N_SN_c_346_n N_A_428_89#_M1002_g 0.00592686f $X=1.405 $Y=0.985 $X2=4.565
+ $Y2=0.835
cc_381 N_SN_c_346_n N_A_428_89#_c_1002_n 0.0167385f $X=1.405 $Y=0.985 $X2=5.57
+ $Y2=0.755
cc_382 N_SN_c_346_n N_A_970_89#_M1004_s 5.44275e-19 $X=1.405 $Y=0.985 $X2=5.965
+ $Y2=0.575
cc_383 N_SN_c_346_n N_A_970_89#_M1006_g 0.00549553f $X=1.405 $Y=0.985 $X2=4.925
+ $Y2=0.835
cc_384 N_SN_M1016_g N_A_970_89#_c_1187_n 0.00575596f $X=6.735 $Y=3.445 $X2=7.57
+ $Y2=1.71
cc_385 N_SN_c_340_n N_A_970_89#_c_1188_n 5.94331e-19 $X=6.735 $Y=1.232 $X2=7.572
+ $Y2=1.545
cc_386 N_SN_c_340_n N_A_970_89#_c_1189_n 0.00206122f $X=6.735 $Y=1.232 $X2=7.66
+ $Y2=1.17
cc_387 N_SN_c_340_n N_A_970_89#_c_1194_n 0.00399517f $X=6.735 $Y=1.232 $X2=7.66
+ $Y2=1.32
cc_388 N_SN_c_334_n N_A_970_89#_c_1198_n 0.00458594f $X=6.665 $Y=1.04 $X2=6.435
+ $Y2=0.91
cc_389 N_SN_c_346_n N_A_970_89#_c_1198_n 0.0168843f $X=1.405 $Y=0.985 $X2=6.435
+ $Y2=0.91
cc_390 N_SN_c_334_n N_A_970_89#_c_1201_n 0.00114006f $X=6.665 $Y=1.04 $X2=6.52
+ $Y2=1.625
cc_391 N_SN_M1016_g N_A_970_89#_c_1201_n 0.0047492f $X=6.735 $Y=3.445 $X2=6.52
+ $Y2=1.625
cc_392 N_SN_c_340_n N_A_970_89#_c_1201_n 0.0101217f $X=6.735 $Y=1.232 $X2=6.52
+ $Y2=1.625
cc_393 N_SN_c_343_n N_A_970_89#_c_1201_n 0.0158894f $X=6.94 $Y=1.165 $X2=6.52
+ $Y2=1.625
cc_394 N_SN_c_346_n N_A_970_89#_c_1201_n 0.0163452f $X=1.405 $Y=0.985 $X2=6.52
+ $Y2=1.625
cc_395 N_SN_M1016_g N_A_970_89#_c_1202_n 0.0312089f $X=6.735 $Y=3.445 $X2=6.52
+ $Y2=3.615
cc_396 N_SN_M1016_g N_A_970_89#_c_1203_n 0.0140658f $X=6.735 $Y=3.445 $X2=7.57
+ $Y2=1.71
cc_397 N_SN_c_340_n N_A_970_89#_c_1203_n 0.00568865f $X=6.735 $Y=1.232 $X2=7.57
+ $Y2=1.71
cc_398 N_SN_c_343_n N_A_970_89#_c_1203_n 0.0120162f $X=6.94 $Y=1.165 $X2=7.57
+ $Y2=1.71
cc_399 N_SN_c_346_n N_A_970_89#_c_1203_n 0.0038502f $X=1.405 $Y=0.985 $X2=7.57
+ $Y2=1.71
cc_400 N_SN_c_346_n N_A_970_89#_c_1204_n 0.00732645f $X=1.405 $Y=0.985 $X2=6.09
+ $Y2=0.74
cc_401 N_SN_M1016_g N_A_970_89#_c_1211_n 0.0113977f $X=6.735 $Y=3.445 $X2=7.425
+ $Y2=1.71
cc_402 N_SN_c_340_n N_A_970_89#_c_1211_n 0.00365839f $X=6.735 $Y=1.232 $X2=7.425
+ $Y2=1.71
cc_403 N_SN_c_343_n N_A_970_89#_c_1211_n 0.00262432f $X=6.94 $Y=1.165 $X2=7.425
+ $Y2=1.71
cc_404 N_SN_c_346_n N_A_970_89#_c_1211_n 0.019887f $X=1.405 $Y=0.985 $X2=7.425
+ $Y2=1.71
cc_405 N_SN_M1016_g N_A_970_89#_c_1213_n 7.50694e-19 $X=6.735 $Y=3.445 $X2=7.57
+ $Y2=1.71
cc_406 N_SN_c_346_n N_A_808_115#_M1010_d 0.0033686f $X=1.405 $Y=0.985 $X2=4.04
+ $Y2=0.575
cc_407 N_SN_c_334_n N_A_808_115#_M1004_g 0.0300902f $X=6.665 $Y=1.04 $X2=6.305
+ $Y2=0.755
cc_408 N_SN_c_346_n N_A_808_115#_M1004_g 0.00640862f $X=1.405 $Y=0.985 $X2=6.305
+ $Y2=0.755
cc_409 N_SN_M1016_g N_A_808_115#_c_1382_n 0.0795539f $X=6.735 $Y=3.445 $X2=6.305
+ $Y2=1.37
cc_410 N_SN_c_340_n N_A_808_115#_c_1382_n 0.0300902f $X=6.735 $Y=1.232 $X2=6.305
+ $Y2=1.37
cc_411 N_SN_c_346_n N_A_808_115#_c_1382_n 0.00408776f $X=1.405 $Y=0.985
+ $X2=6.305 $Y2=1.37
cc_412 N_SN_c_346_n N_A_808_115#_c_1383_n 0.00199877f $X=1.405 $Y=0.985
+ $X2=3.685 $Y2=1.37
cc_413 N_SN_c_346_n N_A_808_115#_c_1384_n 0.00457616f $X=1.405 $Y=0.985
+ $X2=4.365 $Y2=1.37
cc_414 N_SN_c_346_n N_A_808_115#_c_1385_n 0.00243761f $X=1.405 $Y=0.985 $X2=6.1
+ $Y2=1.37
cc_415 N_SN_c_346_n N_A_808_115#_c_1386_n 0.0225179f $X=1.405 $Y=0.985 $X2=4.265
+ $Y2=0.755
cc_416 N_SN_c_346_n N_A_808_115#_c_1389_n 0.0319494f $X=1.405 $Y=0.985 $X2=4.245
+ $Y2=1.37
cc_417 N_SN_c_346_n N_A_808_115#_c_1390_n 0.0241315f $X=1.405 $Y=0.985 $X2=3.83
+ $Y2=1.37
cc_418 N_SN_c_346_n N_A_808_115#_c_1391_n 0.115224f $X=1.405 $Y=0.985 $X2=5.955
+ $Y2=1.37
cc_419 N_SN_c_346_n N_A_808_115#_c_1393_n 0.0187045f $X=1.405 $Y=0.985 $X2=4.48
+ $Y2=1.37
cc_420 N_SN_c_346_n N_A_808_115#_c_1394_n 0.0261247f $X=1.405 $Y=0.985 $X2=6.1
+ $Y2=1.37
cc_421 N_SN_c_334_n N_QN_c_1528_n 0.00270711f $X=6.665 $Y=1.04 $X2=7.47 $Y2=0.74
cc_422 N_SN_c_340_n N_QN_c_1528_n 0.00162792f $X=6.735 $Y=1.232 $X2=7.47
+ $Y2=0.74
cc_423 N_SN_c_343_n N_QN_c_1528_n 0.00918877f $X=6.94 $Y=1.165 $X2=7.47 $Y2=0.74
cc_424 N_SN_c_346_n N_QN_c_1528_n 0.00925906f $X=1.405 $Y=0.985 $X2=7.47
+ $Y2=0.74
cc_425 N_SN_M1016_g N_QN_c_1532_n 0.0223105f $X=6.735 $Y=3.445 $X2=7.47 $Y2=2.48
cc_426 N_SN_M1016_g N_QN_c_1535_n 7.97934e-19 $X=6.735 $Y=3.445 $X2=7.555
+ $Y2=1.37
cc_427 N_SN_c_340_n N_QN_c_1535_n 0.00199491f $X=6.735 $Y=1.232 $X2=7.555
+ $Y2=1.37
cc_428 N_SN_c_343_n N_QN_c_1535_n 0.00417626f $X=6.94 $Y=1.165 $X2=7.555
+ $Y2=1.37
cc_429 N_SN_M1016_g N_QN_c_1537_n 0.00454519f $X=6.735 $Y=3.445 $X2=7.555
+ $Y2=2.285
cc_430 N_SN_M1016_g QN 0.00489905f $X=6.735 $Y=3.445 $X2=7.475 $Y2=2.48
cc_431 N_SN_c_346_n A_386_115# 0.00382239f $X=1.405 $Y=0.985 $X2=1.93 $Y2=0.575
cc_432 N_SN_c_346_n A_578_115# 0.00477583f $X=1.405 $Y=0.985 $X2=2.89 $Y2=0.575
cc_433 N_SN_c_346_n A_736_115# 0.00433937f $X=1.405 $Y=0.985 $X2=3.68 $Y2=0.575
cc_434 N_SN_c_346_n A_928_115# 0.00470365f $X=1.405 $Y=0.985 $X2=4.64 $Y2=0.575
cc_435 N_A_152_89#_c_485_n N_D_M1001_g 0.0067352f $X=1.03 $Y=1.925 $X2=1.855
+ $Y2=0.835
cc_436 N_A_152_89#_c_486_n N_D_M1001_g 0.0123567f $X=2.33 $Y=1.285 $X2=1.855
+ $Y2=0.835
cc_437 N_A_152_89#_c_485_n N_D_M1007_g 0.0108821f $X=1.03 $Y=1.925 $X2=1.855
+ $Y2=3.235
cc_438 N_A_152_89#_c_501_n N_D_M1007_g 0.0211938f $X=2.345 $Y=2.705 $X2=1.855
+ $Y2=3.235
cc_439 N_A_152_89#_c_484_n N_D_c_575_n 0.00665334f $X=1.03 $Y=1.925 $X2=1.915
+ $Y2=1.74
cc_440 N_A_152_89#_c_485_n N_D_c_575_n 0.00142467f $X=1.03 $Y=1.925 $X2=1.915
+ $Y2=1.74
cc_441 N_A_152_89#_c_486_n N_D_c_575_n 0.00207628f $X=2.33 $Y=1.285 $X2=1.915
+ $Y2=1.74
cc_442 N_A_152_89#_c_484_n N_D_c_576_n 9.56786e-19 $X=1.03 $Y=1.925 $X2=1.915
+ $Y2=1.74
cc_443 N_A_152_89#_c_486_n N_D_c_576_n 0.0086486f $X=2.33 $Y=1.285 $X2=1.915
+ $Y2=1.74
cc_444 N_A_152_89#_c_484_n D 0.00134429f $X=1.03 $Y=1.925 $X2=1.915 $Y2=1.74
cc_445 N_A_152_89#_c_486_n D 0.00200799f $X=2.33 $Y=1.285 $X2=1.915 $Y2=1.74
cc_446 N_A_152_89#_c_501_n N_CK_M1011_g 0.0153421f $X=2.345 $Y=2.705 $X2=2.215
+ $Y2=3.235
cc_447 N_A_152_89#_c_501_n N_CK_c_613_n 0.00150627f $X=2.345 $Y=2.705 $X2=2.275
+ $Y2=2.285
cc_448 N_A_152_89#_c_486_n N_CK_c_614_n 9.45214e-19 $X=2.33 $Y=1.285 $X2=2.755
+ $Y2=1.37
cc_449 N_A_152_89#_c_492_n N_CK_c_614_n 0.00165184f $X=2.415 $Y=0.755 $X2=2.755
+ $Y2=1.37
cc_450 N_A_152_89#_c_491_n N_CK_c_615_n 0.00476923f $X=2.415 $Y=1.2 $X2=2.755
+ $Y2=1.205
cc_451 N_A_152_89#_c_492_n N_CK_c_615_n 0.00243799f $X=2.415 $Y=0.755 $X2=2.755
+ $Y2=1.205
cc_452 N_A_152_89#_c_486_n N_CK_c_628_n 0.0019742f $X=2.33 $Y=1.285 $X2=2.67
+ $Y2=2.11
cc_453 N_A_152_89#_c_501_n N_CK_c_628_n 0.00883015f $X=2.345 $Y=2.705 $X2=2.67
+ $Y2=2.11
cc_454 N_A_152_89#_c_486_n N_CK_c_629_n 0.012316f $X=2.33 $Y=1.285 $X2=2.755
+ $Y2=1.37
cc_455 N_A_152_89#_c_492_n N_CK_c_629_n 5.6999e-19 $X=2.415 $Y=0.755 $X2=2.755
+ $Y2=1.37
cc_456 N_A_152_89#_c_486_n N_CK_c_634_n 0.00224443f $X=2.33 $Y=1.285 $X2=2.275
+ $Y2=2.11
cc_457 N_A_152_89#_c_501_n N_CK_c_634_n 0.0101098f $X=2.345 $Y=2.705 $X2=2.275
+ $Y2=2.11
cc_458 N_A_152_89#_c_501_n N_CK_c_636_n 0.00601583f $X=2.345 $Y=2.705 $X2=4.36
+ $Y2=2.11
cc_459 N_A_152_89#_c_501_n N_CK_c_637_n 0.00409373f $X=2.345 $Y=2.705 $X2=2.42
+ $Y2=2.11
cc_460 N_A_152_89#_M1000_g N_A_27_115#_c_857_n 0.00475296f $X=0.835 $Y=0.755
+ $X2=0.605 $Y2=0.91
cc_461 N_A_152_89#_M1000_g N_A_27_115#_c_860_n 0.0152082f $X=0.835 $Y=0.755
+ $X2=0.69 $Y2=1.905
cc_462 N_A_152_89#_M1020_g N_A_27_115#_c_860_n 0.0123669f $X=0.905 $Y=3.445
+ $X2=0.69 $Y2=1.905
cc_463 N_A_152_89#_c_484_n N_A_27_115#_c_860_n 0.005601f $X=1.03 $Y=1.925
+ $X2=0.69 $Y2=1.905
cc_464 N_A_152_89#_c_485_n N_A_27_115#_c_860_n 0.0829295f $X=1.03 $Y=1.925
+ $X2=0.69 $Y2=1.905
cc_465 N_A_152_89#_c_489_n N_A_27_115#_c_860_n 0.0125444f $X=1.115 $Y=1.285
+ $X2=0.69 $Y2=1.905
cc_466 N_A_152_89#_c_505_n N_A_27_115#_c_860_n 0.013584f $X=1.115 $Y=2.705
+ $X2=0.69 $Y2=1.905
cc_467 N_A_152_89#_M1000_g N_A_27_115#_c_867_n 0.00239999f $X=0.835 $Y=0.755
+ $X2=0.69 $Y2=1.79
cc_468 N_A_152_89#_c_484_n N_A_27_115#_c_867_n 2.36419e-19 $X=1.03 $Y=1.925
+ $X2=0.69 $Y2=1.79
cc_469 N_A_152_89#_c_485_n N_A_27_115#_c_867_n 0.00741295f $X=1.03 $Y=1.925
+ $X2=0.69 $Y2=1.79
cc_470 N_A_152_89#_M1000_g N_A_27_115#_c_868_n 0.00793273f $X=0.835 $Y=0.755
+ $X2=3.11 $Y2=1.37
cc_471 N_A_152_89#_c_484_n N_A_27_115#_c_868_n 0.00211509f $X=1.03 $Y=1.925
+ $X2=3.11 $Y2=1.37
cc_472 N_A_152_89#_c_485_n N_A_27_115#_c_868_n 0.00987249f $X=1.03 $Y=1.925
+ $X2=3.11 $Y2=1.37
cc_473 N_A_152_89#_c_486_n N_A_27_115#_c_868_n 0.0544147f $X=2.33 $Y=1.285
+ $X2=3.11 $Y2=1.37
cc_474 N_A_152_89#_c_489_n N_A_27_115#_c_868_n 0.00410183f $X=1.115 $Y=1.285
+ $X2=3.11 $Y2=1.37
cc_475 N_A_152_89#_c_492_n N_A_27_115#_c_868_n 9.30236e-19 $X=2.415 $Y=0.755
+ $X2=3.11 $Y2=1.37
cc_476 N_A_152_89#_c_484_n N_A_27_115#_c_870_n 0.00472146f $X=1.03 $Y=1.925
+ $X2=0.69 $Y2=1.905
cc_477 N_A_152_89#_c_485_n N_A_27_115#_c_870_n 0.0060239f $X=1.03 $Y=1.925
+ $X2=0.69 $Y2=1.905
cc_478 N_A_152_89#_c_486_n N_A_428_89#_c_984_n 0.00232293f $X=2.33 $Y=1.285
+ $X2=2.215 $Y2=1.205
cc_479 N_A_152_89#_c_491_n N_A_428_89#_c_984_n 0.00473574f $X=2.415 $Y=1.2
+ $X2=2.215 $Y2=1.205
cc_480 N_A_152_89#_c_492_n N_A_428_89#_c_984_n 0.00116801f $X=2.415 $Y=0.755
+ $X2=2.215 $Y2=1.205
cc_481 N_A_152_89#_c_486_n N_A_428_89#_c_987_n 0.00326059f $X=2.33 $Y=1.285
+ $X2=2.335 $Y2=1.745
cc_482 N_A_152_89#_c_486_n N_A_428_89#_c_988_n 0.00156949f $X=2.33 $Y=1.285
+ $X2=2.74 $Y2=1.82
cc_483 N_A_152_89#_c_486_n N_A_428_89#_c_997_n 0.00984832f $X=2.33 $Y=1.285
+ $X2=2.335 $Y2=1.28
cc_484 N_A_152_89#_c_501_n A_386_521# 0.00732587f $X=2.345 $Y=2.705 $X2=1.93
+ $Y2=2.605
cc_485 N_D_M1007_g N_CK_c_613_n 0.11474f $X=1.855 $Y=3.235 $X2=2.275 $Y2=2.285
cc_486 N_D_c_575_n N_CK_c_629_n 2.89615e-19 $X=1.915 $Y=1.74 $X2=2.755 $Y2=1.37
cc_487 N_D_c_576_n N_CK_c_629_n 0.00478177f $X=1.915 $Y=1.74 $X2=2.755 $Y2=1.37
cc_488 D N_CK_c_629_n 0.00551577f $X=1.915 $Y=1.74 $X2=2.755 $Y2=1.37
cc_489 N_D_M1007_g N_CK_c_634_n 0.00494364f $X=1.855 $Y=3.235 $X2=2.275 $Y2=2.11
cc_490 N_D_M1007_g N_CK_c_637_n 0.00515433f $X=1.855 $Y=3.235 $X2=2.42 $Y2=2.11
cc_491 D N_CK_c_637_n 0.00375733f $X=1.915 $Y=1.74 $X2=2.42 $Y2=2.11
cc_492 N_D_M1001_g N_A_27_115#_c_868_n 0.0030176f $X=1.855 $Y=0.835 $X2=3.11
+ $Y2=1.37
cc_493 N_D_c_575_n N_A_27_115#_c_868_n 7.9412e-19 $X=1.915 $Y=1.74 $X2=3.11
+ $Y2=1.37
cc_494 N_D_c_576_n N_A_27_115#_c_868_n 0.00111625f $X=1.915 $Y=1.74 $X2=3.11
+ $Y2=1.37
cc_495 D N_A_27_115#_c_868_n 0.0353362f $X=1.915 $Y=1.74 $X2=3.11 $Y2=1.37
cc_496 N_D_M1001_g N_A_428_89#_c_984_n 0.0565233f $X=1.855 $Y=0.835 $X2=2.215
+ $Y2=1.205
cc_497 N_D_M1001_g N_A_428_89#_c_987_n 0.00932846f $X=1.855 $Y=0.835 $X2=2.335
+ $Y2=1.745
cc_498 N_D_c_575_n N_A_428_89#_c_987_n 0.0210215f $X=1.915 $Y=1.74 $X2=2.335
+ $Y2=1.745
cc_499 N_D_c_576_n N_A_428_89#_c_987_n 0.00164409f $X=1.915 $Y=1.74 $X2=2.335
+ $Y2=1.745
cc_500 D N_A_428_89#_c_987_n 0.00342011f $X=1.915 $Y=1.74 $X2=2.335 $Y2=1.745
cc_501 D N_A_428_89#_c_989_n 4.62757e-19 $X=1.915 $Y=1.74 $X2=2.41 $Y2=1.82
cc_502 N_CK_c_615_n N_A_27_115#_M1021_g 0.0337508f $X=2.755 $Y=1.205 $X2=3.175
+ $Y2=0.835
cc_503 N_CK_c_629_n N_A_27_115#_M1021_g 0.00109079f $X=2.755 $Y=1.37 $X2=3.175
+ $Y2=0.835
cc_504 N_CK_c_618_n N_A_27_115#_c_848_n 0.0333348f $X=4.025 $Y=1.37 $X2=3.53
+ $Y2=1.37
cc_505 N_CK_c_630_n N_A_27_115#_c_848_n 3.18936e-19 $X=4.025 $Y=1.37 $X2=3.53
+ $Y2=1.37
cc_506 N_CK_c_614_n N_A_27_115#_c_850_n 0.0337508f $X=2.755 $Y=1.37 $X2=3.25
+ $Y2=1.37
cc_507 N_CK_c_636_n N_A_27_115#_c_851_n 0.00772879f $X=4.36 $Y=2.11 $X2=3.53
+ $Y2=2.285
cc_508 N_CK_c_636_n N_A_27_115#_c_852_n 0.00679967f $X=4.36 $Y=2.11 $X2=3.25
+ $Y2=2.285
cc_509 N_CK_c_619_n N_A_27_115#_M1013_g 0.0333348f $X=4.025 $Y=1.205 $X2=3.605
+ $Y2=0.835
cc_510 N_CK_c_614_n N_A_27_115#_c_861_n 7.30049e-19 $X=2.755 $Y=1.37 $X2=3.345
+ $Y2=2.285
cc_511 N_CK_c_628_n N_A_27_115#_c_861_n 0.00401809f $X=2.67 $Y=2.11 $X2=3.345
+ $Y2=2.285
cc_512 N_CK_c_629_n N_A_27_115#_c_861_n 0.0203851f $X=2.755 $Y=1.37 $X2=3.345
+ $Y2=2.285
cc_513 N_CK_c_636_n N_A_27_115#_c_861_n 0.0206884f $X=4.36 $Y=2.11 $X2=3.345
+ $Y2=2.285
cc_514 N_CK_c_614_n N_A_27_115#_c_865_n 7.18106e-19 $X=2.755 $Y=1.37 $X2=3.345
+ $Y2=1.37
cc_515 N_CK_c_629_n N_A_27_115#_c_865_n 0.00742068f $X=2.755 $Y=1.37 $X2=3.345
+ $Y2=1.37
cc_516 N_CK_c_630_n N_A_27_115#_c_865_n 0.00149326f $X=4.025 $Y=1.37 $X2=3.345
+ $Y2=1.37
cc_517 N_CK_c_636_n N_A_27_115#_c_865_n 0.00102309f $X=4.36 $Y=2.11 $X2=3.345
+ $Y2=1.37
cc_518 N_CK_c_614_n N_A_27_115#_c_868_n 0.00387031f $X=2.755 $Y=1.37 $X2=3.11
+ $Y2=1.37
cc_519 N_CK_c_628_n N_A_27_115#_c_868_n 0.00443421f $X=2.67 $Y=2.11 $X2=3.11
+ $Y2=1.37
cc_520 N_CK_c_629_n N_A_27_115#_c_868_n 0.0151309f $X=2.755 $Y=1.37 $X2=3.11
+ $Y2=1.37
cc_521 N_CK_c_634_n N_A_27_115#_c_868_n 7.12046e-19 $X=2.275 $Y=2.11 $X2=3.11
+ $Y2=1.37
cc_522 N_CK_c_637_n N_A_27_115#_c_868_n 0.0126164f $X=2.42 $Y=2.11 $X2=3.11
+ $Y2=1.37
cc_523 N_CK_c_614_n N_A_27_115#_c_913_n 3.3031e-19 $X=2.755 $Y=1.37 $X2=3.255
+ $Y2=1.37
cc_524 N_CK_c_629_n N_A_27_115#_c_913_n 0.00143592f $X=2.755 $Y=1.37 $X2=3.255
+ $Y2=1.37
cc_525 N_CK_c_636_n N_A_27_115#_c_913_n 0.0129652f $X=4.36 $Y=2.11 $X2=3.255
+ $Y2=1.37
cc_526 N_CK_c_615_n N_A_428_89#_c_984_n 0.0168419f $X=2.755 $Y=1.205 $X2=2.215
+ $Y2=1.205
cc_527 N_CK_c_629_n N_A_428_89#_c_987_n 0.00613747f $X=2.755 $Y=1.37 $X2=2.335
+ $Y2=1.745
cc_528 N_CK_c_614_n N_A_428_89#_c_988_n 0.0183603f $X=2.755 $Y=1.37 $X2=2.74
+ $Y2=1.82
cc_529 N_CK_c_629_n N_A_428_89#_c_988_n 0.00630484f $X=2.755 $Y=1.37 $X2=2.74
+ $Y2=1.82
cc_530 N_CK_c_636_n N_A_428_89#_c_988_n 0.00558832f $X=4.36 $Y=2.11 $X2=2.74
+ $Y2=1.82
cc_531 N_CK_c_613_n N_A_428_89#_c_989_n 0.00904036f $X=2.275 $Y=2.285 $X2=2.41
+ $Y2=1.82
cc_532 N_CK_c_628_n N_A_428_89#_c_989_n 0.00810782f $X=2.67 $Y=2.11 $X2=2.41
+ $Y2=1.82
cc_533 N_CK_c_634_n N_A_428_89#_c_989_n 0.00109468f $X=2.275 $Y=2.11 $X2=2.41
+ $Y2=1.82
cc_534 N_CK_c_637_n N_A_428_89#_c_989_n 0.00131242f $X=2.42 $Y=2.11 $X2=2.41
+ $Y2=1.82
cc_535 N_CK_M1011_g N_A_428_89#_M1015_g 0.0316011f $X=2.215 $Y=3.235 $X2=2.815
+ $Y2=3.235
cc_536 N_CK_c_613_n N_A_428_89#_M1015_g 0.0128384f $X=2.275 $Y=2.285 $X2=2.815
+ $Y2=3.235
cc_537 N_CK_c_628_n N_A_428_89#_M1015_g 0.0081071f $X=2.67 $Y=2.11 $X2=2.815
+ $Y2=3.235
cc_538 N_CK_c_629_n N_A_428_89#_M1015_g 0.00478024f $X=2.755 $Y=1.37 $X2=2.815
+ $Y2=3.235
cc_539 N_CK_c_634_n N_A_428_89#_M1015_g 0.00184124f $X=2.275 $Y=2.11 $X2=2.815
+ $Y2=3.235
cc_540 N_CK_c_636_n N_A_428_89#_M1015_g 0.00938974f $X=4.36 $Y=2.11 $X2=2.815
+ $Y2=3.235
cc_541 N_CK_c_637_n N_A_428_89#_M1015_g 4.2e-19 $X=2.42 $Y=2.11 $X2=2.815
+ $Y2=3.235
cc_542 N_CK_c_636_n N_A_428_89#_c_991_n 0.00607908f $X=4.36 $Y=2.11 $X2=3.89
+ $Y2=1.82
cc_543 N_CK_M1028_g N_A_428_89#_M1022_g 0.0316011f $X=4.565 $Y=3.235 $X2=3.965
+ $Y2=3.235
cc_544 N_CK_c_622_n N_A_428_89#_M1022_g 0.0118393f $X=4.505 $Y=2.285 $X2=3.965
+ $Y2=3.235
cc_545 N_CK_c_630_n N_A_428_89#_M1022_g 0.00368284f $X=4.025 $Y=1.37 $X2=3.965
+ $Y2=3.235
cc_546 N_CK_c_632_n N_A_428_89#_M1022_g 0.00654233f $X=4.11 $Y=2.11 $X2=3.965
+ $Y2=3.235
cc_547 N_CK_c_635_n N_A_428_89#_M1022_g 0.00128351f $X=4.505 $Y=2.11 $X2=3.965
+ $Y2=3.235
cc_548 N_CK_c_636_n N_A_428_89#_M1022_g 0.00497421f $X=4.36 $Y=2.11 $X2=3.965
+ $Y2=3.235
cc_549 N_CK_c_639_n N_A_428_89#_M1022_g 4.2e-19 $X=4.65 $Y=2.11 $X2=3.965
+ $Y2=3.235
cc_550 N_CK_c_630_n N_A_428_89#_c_993_n 0.00681452f $X=4.025 $Y=1.37 $X2=4.37
+ $Y2=1.825
cc_551 N_CK_c_631_n N_A_428_89#_c_993_n 0.00791191f $X=4.42 $Y=2.11 $X2=4.37
+ $Y2=1.825
cc_552 N_CK_c_636_n N_A_428_89#_c_993_n 0.00484158f $X=4.36 $Y=2.11 $X2=4.37
+ $Y2=1.825
cc_553 N_CK_c_639_n N_A_428_89#_c_993_n 0.0012566f $X=4.65 $Y=2.11 $X2=4.37
+ $Y2=1.825
cc_554 N_CK_c_618_n N_A_428_89#_M1002_g 0.0126057f $X=4.025 $Y=1.37 $X2=4.565
+ $Y2=0.835
cc_555 N_CK_c_619_n N_A_428_89#_M1002_g 0.0168302f $X=4.025 $Y=1.205 $X2=4.565
+ $Y2=0.835
cc_556 N_CK_c_630_n N_A_428_89#_M1002_g 0.00138616f $X=4.025 $Y=1.37 $X2=4.565
+ $Y2=0.835
cc_557 N_CK_c_614_n N_A_428_89#_c_997_n 0.0216263f $X=2.755 $Y=1.37 $X2=2.335
+ $Y2=1.28
cc_558 N_CK_c_634_n N_A_428_89#_c_997_n 2.45465e-19 $X=2.275 $Y=2.11 $X2=2.335
+ $Y2=1.28
cc_559 N_CK_c_629_n N_A_428_89#_c_998_n 0.00568091f $X=2.755 $Y=1.37 $X2=2.815
+ $Y2=1.82
cc_560 N_CK_c_618_n N_A_428_89#_c_999_n 0.0183777f $X=4.025 $Y=1.37 $X2=3.965
+ $Y2=1.825
cc_561 N_CK_c_630_n N_A_428_89#_c_999_n 0.00451735f $X=4.025 $Y=1.37 $X2=3.965
+ $Y2=1.825
cc_562 N_CK_c_622_n N_A_428_89#_c_1000_n 0.0173927f $X=4.505 $Y=2.285 $X2=4.505
+ $Y2=1.74
cc_563 N_CK_c_630_n N_A_428_89#_c_1000_n 0.00341807f $X=4.025 $Y=1.37 $X2=4.505
+ $Y2=1.74
cc_564 N_CK_c_635_n N_A_428_89#_c_1000_n 0.00108517f $X=4.505 $Y=2.11 $X2=4.505
+ $Y2=1.74
cc_565 N_CK_c_622_n N_A_428_89#_c_1001_n 7.72371e-19 $X=4.505 $Y=2.285 $X2=4.505
+ $Y2=1.74
cc_566 N_CK_c_630_n N_A_428_89#_c_1001_n 0.00896072f $X=4.025 $Y=1.37 $X2=4.505
+ $Y2=1.74
cc_567 N_CK_c_631_n N_A_428_89#_c_1001_n 0.00449061f $X=4.42 $Y=2.11 $X2=4.505
+ $Y2=1.74
cc_568 N_CK_c_635_n N_A_428_89#_c_1001_n 0.00979766f $X=4.505 $Y=2.11 $X2=4.505
+ $Y2=1.74
cc_569 N_CK_c_639_n N_A_428_89#_c_1001_n 0.00182452f $X=4.65 $Y=2.11 $X2=4.505
+ $Y2=1.74
cc_570 N_CK_c_623_n N_A_428_89#_c_1002_n 0.00779247f $X=5.382 $Y=1.205 $X2=5.57
+ $Y2=0.755
cc_571 N_CK_c_627_n N_A_428_89#_c_1002_n 0.0121392f $X=5.382 $Y=1.355 $X2=5.57
+ $Y2=0.755
cc_572 N_CK_c_611_n N_A_428_89#_c_1006_n 0.0031983f $X=5.355 $Y=2.45 $X2=5.845
+ $Y2=2.62
cc_573 N_CK_M1017_g N_A_428_89#_c_1006_n 0.00397698f $X=5.355 $Y=3.235 $X2=5.845
+ $Y2=2.62
cc_574 N_CK_c_612_n N_A_428_89#_c_1006_n 0.00565489f $X=5.41 $Y=2.12 $X2=5.845
+ $Y2=2.62
cc_575 N_CK_c_633_n N_A_428_89#_c_1006_n 0.0277249f $X=5.5 $Y=2.11 $X2=5.845
+ $Y2=2.62
cc_576 CK N_A_428_89#_c_1006_n 0.00230094f $X=5.5 $Y=2.11 $X2=5.845 $Y2=2.62
cc_577 N_CK_c_611_n N_A_428_89#_c_1022_n 0.00233394f $X=5.355 $Y=2.45 $X2=5.845
+ $Y2=2.705
cc_578 N_CK_c_633_n N_A_428_89#_c_1022_n 0.00601935f $X=5.5 $Y=2.11 $X2=5.845
+ $Y2=2.705
cc_579 N_CK_c_611_n N_A_428_89#_c_1007_n 0.00187011f $X=5.355 $Y=2.45 $X2=5.57
+ $Y2=1.755
cc_580 N_CK_c_612_n N_A_428_89#_c_1007_n 0.00802926f $X=5.41 $Y=2.12 $X2=5.57
+ $Y2=1.755
cc_581 N_CK_c_633_n N_A_428_89#_c_1007_n 0.0100792f $X=5.5 $Y=2.11 $X2=5.57
+ $Y2=1.755
cc_582 CK N_A_428_89#_c_1007_n 0.00100188f $X=5.5 $Y=2.11 $X2=5.57 $Y2=1.755
cc_583 N_CK_c_612_n N_A_428_89#_c_1008_n 0.00220085f $X=5.41 $Y=2.12 $X2=5.405
+ $Y2=1.74
cc_584 N_CK_c_627_n N_A_428_89#_c_1008_n 2.6895e-19 $X=5.382 $Y=1.355 $X2=5.405
+ $Y2=1.74
cc_585 N_CK_c_638_n N_A_428_89#_c_1008_n 0.0583359f $X=5.355 $Y=2.11 $X2=5.405
+ $Y2=1.74
cc_586 CK N_A_428_89#_c_1008_n 0.00451538f $X=5.5 $Y=2.11 $X2=5.405 $Y2=1.74
cc_587 N_CK_c_630_n N_A_428_89#_c_1009_n 0.00365074f $X=4.025 $Y=1.37 $X2=4.65
+ $Y2=1.74
cc_588 N_CK_c_635_n N_A_428_89#_c_1009_n 4.76324e-19 $X=4.505 $Y=2.11 $X2=4.65
+ $Y2=1.74
cc_589 N_CK_c_639_n N_A_428_89#_c_1009_n 0.0296305f $X=4.65 $Y=2.11 $X2=4.65
+ $Y2=1.74
cc_590 N_CK_c_612_n N_A_428_89#_c_1010_n 0.00214951f $X=5.41 $Y=2.12 $X2=5.52
+ $Y2=1.74
cc_591 N_CK_c_633_n N_A_428_89#_c_1010_n 6.27299e-19 $X=5.5 $Y=2.11 $X2=5.52
+ $Y2=1.74
cc_592 CK N_A_428_89#_c_1010_n 0.0237732f $X=5.5 $Y=2.11 $X2=5.52 $Y2=1.74
cc_593 N_CK_c_612_n N_A_970_89#_M1006_g 0.00751867f $X=5.41 $Y=2.12 $X2=4.925
+ $Y2=0.835
cc_594 N_CK_c_623_n N_A_970_89#_M1006_g 0.0241221f $X=5.382 $Y=1.205 $X2=4.925
+ $Y2=0.835
cc_595 N_CK_c_611_n N_A_970_89#_M1026_g 0.0406479f $X=5.355 $Y=2.45 $X2=4.925
+ $Y2=3.235
cc_596 N_CK_c_612_n N_A_970_89#_M1026_g 0.0149738f $X=5.41 $Y=2.12 $X2=4.925
+ $Y2=3.235
cc_597 N_CK_c_622_n N_A_970_89#_M1026_g 0.11306f $X=4.505 $Y=2.285 $X2=4.925
+ $Y2=3.235
cc_598 N_CK_c_633_n N_A_970_89#_M1026_g 5.92505e-19 $X=5.5 $Y=2.11 $X2=4.925
+ $Y2=3.235
cc_599 N_CK_c_635_n N_A_970_89#_M1026_g 0.0022769f $X=4.505 $Y=2.11 $X2=4.925
+ $Y2=3.235
cc_600 N_CK_c_638_n N_A_970_89#_M1026_g 0.0028722f $X=5.355 $Y=2.11 $X2=4.925
+ $Y2=3.235
cc_601 N_CK_c_639_n N_A_970_89#_M1026_g 0.00113587f $X=4.65 $Y=2.11 $X2=4.925
+ $Y2=3.235
cc_602 N_CK_c_612_n N_A_970_89#_c_1185_n 0.0207577f $X=5.41 $Y=2.12 $X2=4.985
+ $Y2=1.71
cc_603 N_CK_c_638_n N_A_970_89#_c_1185_n 7.89968e-19 $X=5.355 $Y=2.11 $X2=4.985
+ $Y2=1.71
cc_604 N_CK_c_611_n N_A_970_89#_c_1197_n 0.00273823f $X=5.355 $Y=2.45 $X2=4.985
+ $Y2=1.71
cc_605 N_CK_c_612_n N_A_970_89#_c_1197_n 0.00560687f $X=5.41 $Y=2.12 $X2=4.985
+ $Y2=1.71
cc_606 N_CK_c_622_n N_A_970_89#_c_1197_n 0.00225319f $X=4.505 $Y=2.285 $X2=4.985
+ $Y2=1.71
cc_607 N_CK_c_633_n N_A_970_89#_c_1197_n 0.0147178f $X=5.5 $Y=2.11 $X2=4.985
+ $Y2=1.71
cc_608 N_CK_c_635_n N_A_970_89#_c_1197_n 0.0150823f $X=4.505 $Y=2.11 $X2=4.985
+ $Y2=1.71
cc_609 N_CK_c_638_n N_A_970_89#_c_1197_n 0.0137913f $X=5.355 $Y=2.11 $X2=4.985
+ $Y2=1.71
cc_610 N_CK_c_639_n N_A_970_89#_c_1197_n 0.00206138f $X=4.65 $Y=2.11 $X2=4.985
+ $Y2=1.71
cc_611 CK N_A_970_89#_c_1197_n 0.00189954f $X=5.5 $Y=2.11 $X2=4.985 $Y2=1.71
cc_612 N_CK_c_611_n N_A_970_89#_c_1208_n 0.00430081f $X=5.355 $Y=2.45 $X2=5.785
+ $Y2=2.48
cc_613 N_CK_M1017_g N_A_970_89#_c_1208_n 0.00886028f $X=5.355 $Y=3.235 $X2=5.785
+ $Y2=2.48
cc_614 N_CK_c_633_n N_A_970_89#_c_1208_n 0.00644495f $X=5.5 $Y=2.11 $X2=5.785
+ $Y2=2.48
cc_615 N_CK_c_638_n N_A_970_89#_c_1208_n 0.0190773f $X=5.355 $Y=2.11 $X2=5.785
+ $Y2=2.48
cc_616 CK N_A_970_89#_c_1208_n 0.025144f $X=5.5 $Y=2.11 $X2=5.785 $Y2=2.48
cc_617 N_CK_c_611_n N_A_970_89#_c_1209_n 4.83733e-19 $X=5.355 $Y=2.45 $X2=5.13
+ $Y2=2.48
cc_618 N_CK_M1017_g N_A_970_89#_c_1209_n 4.63789e-19 $X=5.355 $Y=3.235 $X2=5.13
+ $Y2=2.48
cc_619 N_CK_c_622_n N_A_970_89#_c_1209_n 0.00405956f $X=4.505 $Y=2.285 $X2=5.13
+ $Y2=2.48
cc_620 N_CK_c_633_n N_A_970_89#_c_1209_n 7.98697e-19 $X=5.5 $Y=2.11 $X2=5.13
+ $Y2=2.48
cc_621 N_CK_c_635_n N_A_970_89#_c_1209_n 0.0025579f $X=4.505 $Y=2.11 $X2=5.13
+ $Y2=2.48
cc_622 N_CK_c_638_n N_A_970_89#_c_1209_n 0.0253115f $X=5.355 $Y=2.11 $X2=5.13
+ $Y2=2.48
cc_623 N_CK_c_633_n N_A_970_89#_c_1210_n 0.00132196f $X=5.5 $Y=2.11 $X2=5.882
+ $Y2=2.39
cc_624 CK N_A_970_89#_c_1210_n 0.0218354f $X=5.5 $Y=2.11 $X2=5.882 $Y2=2.39
cc_625 N_CK_c_611_n N_A_808_115#_M1024_g 0.00467255f $X=5.355 $Y=2.45 $X2=6.305
+ $Y2=3.445
cc_626 N_CK_c_627_n N_A_808_115#_c_1382_n 0.00712865f $X=5.382 $Y=1.355
+ $X2=6.305 $Y2=1.37
cc_627 N_CK_c_618_n N_A_808_115#_c_1383_n 0.00187586f $X=4.025 $Y=1.37 $X2=3.685
+ $Y2=1.37
cc_628 N_CK_c_630_n N_A_808_115#_c_1383_n 0.0535471f $X=4.025 $Y=1.37 $X2=3.685
+ $Y2=1.37
cc_629 N_CK_c_632_n N_A_808_115#_c_1383_n 0.0116326f $X=4.11 $Y=2.11 $X2=3.685
+ $Y2=1.37
cc_630 N_CK_c_635_n N_A_808_115#_c_1383_n 0.00613815f $X=4.505 $Y=2.11 $X2=3.685
+ $Y2=1.37
cc_631 N_CK_c_636_n N_A_808_115#_c_1383_n 0.020361f $X=4.36 $Y=2.11 $X2=3.685
+ $Y2=1.37
cc_632 N_CK_c_639_n N_A_808_115#_c_1383_n 6.61118e-19 $X=4.65 $Y=2.11 $X2=3.685
+ $Y2=1.37
cc_633 N_CK_c_622_n N_A_808_115#_c_1426_n 0.00150627f $X=4.505 $Y=2.285
+ $X2=4.095 $Y2=2.705
cc_634 N_CK_c_631_n N_A_808_115#_c_1426_n 0.00843004f $X=4.42 $Y=2.11 $X2=4.095
+ $Y2=2.705
cc_635 N_CK_c_632_n N_A_808_115#_c_1426_n 0.00323798f $X=4.11 $Y=2.11 $X2=4.095
+ $Y2=2.705
cc_636 N_CK_c_635_n N_A_808_115#_c_1426_n 0.00103871f $X=4.505 $Y=2.11 $X2=4.095
+ $Y2=2.705
cc_637 N_CK_c_636_n N_A_808_115#_c_1426_n 0.012754f $X=4.36 $Y=2.11 $X2=4.095
+ $Y2=2.705
cc_638 N_CK_c_639_n N_A_808_115#_c_1426_n 0.00146098f $X=4.65 $Y=2.11 $X2=4.095
+ $Y2=2.705
cc_639 N_CK_c_618_n N_A_808_115#_c_1384_n 0.00154744f $X=4.025 $Y=1.37 $X2=4.365
+ $Y2=1.37
cc_640 N_CK_c_619_n N_A_808_115#_c_1384_n 0.00334187f $X=4.025 $Y=1.205
+ $X2=4.365 $Y2=1.37
cc_641 N_CK_c_630_n N_A_808_115#_c_1384_n 0.016958f $X=4.025 $Y=1.37 $X2=4.365
+ $Y2=1.37
cc_642 N_CK_c_631_n N_A_808_115#_c_1384_n 0.00112312f $X=4.42 $Y=2.11 $X2=4.365
+ $Y2=1.37
cc_643 N_CK_c_636_n N_A_808_115#_c_1384_n 2.80397e-19 $X=4.36 $Y=2.11 $X2=4.365
+ $Y2=1.37
cc_644 N_CK_c_618_n N_A_808_115#_c_1386_n 0.00191034f $X=4.025 $Y=1.37 $X2=4.265
+ $Y2=0.755
cc_645 N_CK_c_619_n N_A_808_115#_c_1386_n 0.00389012f $X=4.025 $Y=1.205
+ $X2=4.265 $Y2=0.755
cc_646 N_CK_c_630_n N_A_808_115#_c_1386_n 9.06033e-19 $X=4.025 $Y=1.37 $X2=4.265
+ $Y2=0.755
cc_647 N_CK_c_618_n N_A_808_115#_c_1389_n 0.00424711f $X=4.025 $Y=1.37 $X2=4.245
+ $Y2=1.37
cc_648 N_CK_c_630_n N_A_808_115#_c_1389_n 0.0125093f $X=4.025 $Y=1.37 $X2=4.245
+ $Y2=1.37
cc_649 N_CK_c_631_n N_A_808_115#_c_1389_n 0.00222579f $X=4.42 $Y=2.11 $X2=4.245
+ $Y2=1.37
cc_650 N_CK_c_618_n N_A_808_115#_c_1390_n 3.96626e-19 $X=4.025 $Y=1.37 $X2=3.83
+ $Y2=1.37
cc_651 N_CK_c_630_n N_A_808_115#_c_1390_n 6.47111e-19 $X=4.025 $Y=1.37 $X2=3.83
+ $Y2=1.37
cc_652 N_CK_c_636_n N_A_808_115#_c_1390_n 0.0128239f $X=4.36 $Y=2.11 $X2=3.83
+ $Y2=1.37
cc_653 N_CK_c_612_n N_A_808_115#_c_1391_n 0.00311774f $X=5.41 $Y=2.12 $X2=5.955
+ $Y2=1.37
cc_654 N_CK_c_627_n N_A_808_115#_c_1391_n 0.00385755f $X=5.382 $Y=1.355
+ $X2=5.955 $Y2=1.37
cc_655 N_CK_c_618_n N_A_808_115#_c_1393_n 4.32425e-19 $X=4.025 $Y=1.37 $X2=4.48
+ $Y2=1.37
cc_656 N_CK_c_630_n N_A_808_115#_c_1393_n 0.00112437f $X=4.025 $Y=1.37 $X2=4.48
+ $Y2=1.37
cc_657 N_CK_c_631_n N_A_808_115#_c_1393_n 5.56901e-19 $X=4.42 $Y=2.11 $X2=4.48
+ $Y2=1.37
cc_658 N_CK_c_636_n N_A_808_115#_c_1393_n 0.00585497f $X=4.36 $Y=2.11 $X2=4.48
+ $Y2=1.37
cc_659 N_A_27_115#_c_868_n N_A_428_89#_c_987_n 0.00253253f $X=3.11 $Y=1.37
+ $X2=2.335 $Y2=1.745
cc_660 N_A_27_115#_c_868_n N_A_428_89#_c_988_n 0.004711f $X=3.11 $Y=1.37
+ $X2=2.74 $Y2=1.82
cc_661 N_A_27_115#_c_852_n N_A_428_89#_M1015_g 0.114035f $X=3.25 $Y=2.285
+ $X2=2.815 $Y2=3.235
cc_662 N_A_27_115#_c_861_n N_A_428_89#_M1015_g 0.00486364f $X=3.345 $Y=2.285
+ $X2=2.815 $Y2=3.235
cc_663 N_A_27_115#_c_850_n N_A_428_89#_c_991_n 0.0342351f $X=3.25 $Y=1.37
+ $X2=3.89 $Y2=1.82
cc_664 N_A_27_115#_c_852_n N_A_428_89#_c_991_n 0.0307748f $X=3.25 $Y=2.285
+ $X2=3.89 $Y2=1.82
cc_665 N_A_27_115#_c_861_n N_A_428_89#_c_991_n 0.0113171f $X=3.345 $Y=2.285
+ $X2=3.89 $Y2=1.82
cc_666 N_A_27_115#_c_865_n N_A_428_89#_c_991_n 8.69982e-19 $X=3.345 $Y=1.37
+ $X2=3.89 $Y2=1.82
cc_667 N_A_27_115#_c_868_n N_A_428_89#_c_991_n 0.00486036f $X=3.11 $Y=1.37
+ $X2=3.89 $Y2=1.82
cc_668 N_A_27_115#_c_913_n N_A_428_89#_c_991_n 4.12801e-19 $X=3.255 $Y=1.37
+ $X2=3.89 $Y2=1.82
cc_669 N_A_27_115#_c_851_n N_A_428_89#_M1022_g 0.110621f $X=3.53 $Y=2.285
+ $X2=3.965 $Y2=3.235
cc_670 N_A_27_115#_M1014_g N_A_808_115#_c_1383_n 9.36754e-19 $X=3.175 $Y=3.235
+ $X2=3.685 $Y2=1.37
cc_671 N_A_27_115#_c_848_n N_A_808_115#_c_1383_n 0.00757614f $X=3.53 $Y=1.37
+ $X2=3.685 $Y2=1.37
cc_672 N_A_27_115#_c_851_n N_A_808_115#_c_1383_n 0.00738718f $X=3.53 $Y=2.285
+ $X2=3.685 $Y2=1.37
cc_673 N_A_27_115#_M1005_g N_A_808_115#_c_1383_n 0.00479454f $X=3.605 $Y=3.235
+ $X2=3.685 $Y2=1.37
cc_674 N_A_27_115#_c_861_n N_A_808_115#_c_1383_n 0.0702347f $X=3.345 $Y=2.285
+ $X2=3.685 $Y2=1.37
cc_675 N_A_27_115#_c_865_n N_A_808_115#_c_1383_n 0.0122452f $X=3.345 $Y=1.37
+ $X2=3.685 $Y2=1.37
cc_676 N_A_27_115#_c_913_n N_A_808_115#_c_1383_n 4.18442e-19 $X=3.255 $Y=1.37
+ $X2=3.685 $Y2=1.37
cc_677 N_A_27_115#_M1014_g N_A_808_115#_c_1459_n 9.13132e-19 $X=3.175 $Y=3.235
+ $X2=3.77 $Y2=2.705
cc_678 N_A_27_115#_M1005_g N_A_808_115#_c_1459_n 0.0096885f $X=3.605 $Y=3.235
+ $X2=3.77 $Y2=2.705
cc_679 N_A_27_115#_c_848_n N_A_808_115#_c_1390_n 0.00311393f $X=3.53 $Y=1.37
+ $X2=3.83 $Y2=1.37
cc_680 N_A_27_115#_c_865_n N_A_808_115#_c_1390_n 0.0012094f $X=3.345 $Y=1.37
+ $X2=3.83 $Y2=1.37
cc_681 N_A_27_115#_c_913_n N_A_808_115#_c_1390_n 0.0241863f $X=3.255 $Y=1.37
+ $X2=3.83 $Y2=1.37
cc_682 N_A_27_115#_c_857_n A_110_115# 0.00176584f $X=0.605 $Y=0.91 $X2=0.55
+ $Y2=0.575
cc_683 N_A_428_89#_M1002_g N_A_970_89#_M1006_g 0.0469043f $X=4.565 $Y=0.835
+ $X2=4.925 $Y2=0.835
cc_684 N_A_428_89#_c_1000_n N_A_970_89#_c_1185_n 0.0469043f $X=4.505 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_685 N_A_428_89#_c_1001_n N_A_970_89#_c_1185_n 7.65216e-19 $X=4.505 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_686 N_A_428_89#_c_1007_n N_A_970_89#_c_1185_n 6.62226e-19 $X=5.57 $Y=1.755
+ $X2=4.985 $Y2=1.71
cc_687 N_A_428_89#_c_1008_n N_A_970_89#_c_1185_n 0.00324237f $X=5.405 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_688 N_A_428_89#_c_1009_n N_A_970_89#_c_1185_n 8.85796e-19 $X=4.65 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_689 N_A_428_89#_c_1010_n N_A_970_89#_c_1185_n 3.05538e-19 $X=5.52 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_690 N_A_428_89#_M1002_g N_A_970_89#_c_1197_n 6.69335e-19 $X=4.565 $Y=0.835
+ $X2=4.985 $Y2=1.71
cc_691 N_A_428_89#_c_1000_n N_A_970_89#_c_1197_n 8.11022e-19 $X=4.505 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_692 N_A_428_89#_c_1001_n N_A_970_89#_c_1197_n 0.00843011f $X=4.505 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_693 N_A_428_89#_c_1002_n N_A_970_89#_c_1197_n 0.00363008f $X=5.57 $Y=0.755
+ $X2=4.985 $Y2=1.71
cc_694 N_A_428_89#_c_1007_n N_A_970_89#_c_1197_n 0.00504343f $X=5.57 $Y=1.755
+ $X2=4.985 $Y2=1.71
cc_695 N_A_428_89#_c_1008_n N_A_970_89#_c_1197_n 0.012434f $X=5.405 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_696 N_A_428_89#_c_1009_n N_A_970_89#_c_1197_n 0.00248328f $X=4.65 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_697 N_A_428_89#_c_1010_n N_A_970_89#_c_1197_n 0.00129444f $X=5.52 $Y=1.74
+ $X2=4.985 $Y2=1.71
cc_698 N_A_428_89#_c_1006_n N_A_970_89#_c_1202_n 0.0172245f $X=5.845 $Y=2.62
+ $X2=6.52 $Y2=3.615
cc_699 N_A_428_89#_c_1022_n N_A_970_89#_c_1202_n 0.00644034f $X=5.845 $Y=2.705
+ $X2=6.52 $Y2=3.615
cc_700 N_A_428_89#_c_1007_n N_A_970_89#_c_1202_n 0.00131397f $X=5.57 $Y=1.755
+ $X2=6.52 $Y2=3.615
cc_701 N_A_428_89#_c_1002_n N_A_970_89#_c_1204_n 0.0171447f $X=5.57 $Y=0.755
+ $X2=6.09 $Y2=0.74
cc_702 N_A_428_89#_c_1007_n N_A_970_89#_c_1207_n 0.00245266f $X=5.57 $Y=1.755
+ $X2=6.52 $Y2=1.71
cc_703 N_A_428_89#_c_1006_n N_A_970_89#_c_1208_n 0.0142483f $X=5.845 $Y=2.62
+ $X2=5.785 $Y2=2.48
cc_704 N_A_428_89#_c_1022_n N_A_970_89#_c_1208_n 0.0135048f $X=5.845 $Y=2.705
+ $X2=5.785 $Y2=2.48
cc_705 N_A_428_89#_c_1007_n N_A_970_89#_c_1208_n 0.00314001f $X=5.57 $Y=1.755
+ $X2=5.785 $Y2=2.48
cc_706 N_A_428_89#_c_1010_n N_A_970_89#_c_1208_n 9.06726e-19 $X=5.52 $Y=1.74
+ $X2=5.785 $Y2=2.48
cc_707 N_A_428_89#_c_1006_n N_A_970_89#_c_1210_n 0.0193217f $X=5.845 $Y=2.62
+ $X2=5.882 $Y2=2.39
cc_708 N_A_428_89#_c_1007_n N_A_970_89#_c_1210_n 0.00221219f $X=5.57 $Y=1.755
+ $X2=5.882 $Y2=2.39
cc_709 N_A_428_89#_c_1002_n N_A_970_89#_c_1212_n 2.51414e-19 $X=5.57 $Y=0.755
+ $X2=5.96 $Y2=1.71
cc_710 N_A_428_89#_c_1007_n N_A_970_89#_c_1212_n 0.00850958f $X=5.57 $Y=1.755
+ $X2=5.96 $Y2=1.71
cc_711 N_A_428_89#_c_1010_n N_A_970_89#_c_1212_n 0.0236753f $X=5.52 $Y=1.74
+ $X2=5.96 $Y2=1.71
cc_712 N_A_428_89#_c_1002_n N_A_808_115#_M1004_g 0.00411661f $X=5.57 $Y=0.755
+ $X2=6.305 $Y2=0.755
cc_713 N_A_428_89#_c_1002_n N_A_808_115#_M1024_g 0.00240207f $X=5.57 $Y=0.755
+ $X2=6.305 $Y2=3.445
cc_714 N_A_428_89#_c_1017_n N_A_808_115#_M1024_g 0.0139389f $X=5.57 $Y=2.955
+ $X2=6.305 $Y2=3.445
cc_715 N_A_428_89#_c_1006_n N_A_808_115#_M1024_g 0.0106651f $X=5.845 $Y=2.62
+ $X2=6.305 $Y2=3.445
cc_716 N_A_428_89#_c_1022_n N_A_808_115#_M1024_g 0.00343288f $X=5.845 $Y=2.705
+ $X2=6.305 $Y2=3.445
cc_717 N_A_428_89#_c_1007_n N_A_808_115#_M1024_g 0.00307177f $X=5.57 $Y=1.755
+ $X2=6.305 $Y2=3.445
cc_718 N_A_428_89#_c_1010_n N_A_808_115#_M1024_g 2.03588e-19 $X=5.52 $Y=1.74
+ $X2=6.305 $Y2=3.445
cc_719 N_A_428_89#_c_1002_n N_A_808_115#_c_1382_n 0.00361086f $X=5.57 $Y=0.755
+ $X2=6.305 $Y2=1.37
cc_720 N_A_428_89#_c_991_n N_A_808_115#_c_1383_n 0.0122693f $X=3.89 $Y=1.82
+ $X2=3.685 $Y2=1.37
cc_721 N_A_428_89#_c_999_n N_A_808_115#_c_1383_n 0.0112175f $X=3.965 $Y=1.825
+ $X2=3.685 $Y2=1.37
cc_722 N_A_428_89#_M1022_g N_A_808_115#_c_1426_n 0.0162544f $X=3.965 $Y=3.235
+ $X2=4.095 $Y2=2.705
cc_723 N_A_428_89#_c_993_n N_A_808_115#_c_1384_n 0.0013046f $X=4.37 $Y=1.825
+ $X2=4.365 $Y2=1.37
cc_724 N_A_428_89#_c_1000_n N_A_808_115#_c_1384_n 0.0019411f $X=4.505 $Y=1.74
+ $X2=4.365 $Y2=1.37
cc_725 N_A_428_89#_c_1001_n N_A_808_115#_c_1384_n 0.00640334f $X=4.505 $Y=1.74
+ $X2=4.365 $Y2=1.37
cc_726 N_A_428_89#_c_1009_n N_A_808_115#_c_1384_n 2.54388e-19 $X=4.65 $Y=1.74
+ $X2=4.365 $Y2=1.37
cc_727 N_A_428_89#_c_1002_n N_A_808_115#_c_1385_n 0.00736723f $X=5.57 $Y=0.755
+ $X2=6.1 $Y2=1.37
cc_728 N_A_428_89#_M1002_g N_A_808_115#_c_1386_n 0.0129399f $X=4.565 $Y=0.835
+ $X2=4.265 $Y2=0.755
cc_729 N_A_428_89#_c_991_n N_A_808_115#_c_1389_n 0.00156696f $X=3.89 $Y=1.82
+ $X2=4.245 $Y2=1.37
cc_730 N_A_428_89#_c_993_n N_A_808_115#_c_1389_n 0.00173579f $X=4.37 $Y=1.825
+ $X2=4.245 $Y2=1.37
cc_731 N_A_428_89#_c_999_n N_A_808_115#_c_1389_n 5.21392e-19 $X=3.965 $Y=1.825
+ $X2=4.245 $Y2=1.37
cc_732 N_A_428_89#_c_991_n N_A_808_115#_c_1390_n 0.00120486f $X=3.89 $Y=1.82
+ $X2=3.83 $Y2=1.37
cc_733 N_A_428_89#_M1002_g N_A_808_115#_c_1391_n 0.00522039f $X=4.565 $Y=0.835
+ $X2=5.955 $Y2=1.37
cc_734 N_A_428_89#_c_1001_n N_A_808_115#_c_1391_n 0.00245278f $X=4.505 $Y=1.74
+ $X2=5.955 $Y2=1.37
cc_735 N_A_428_89#_c_1002_n N_A_808_115#_c_1391_n 0.0167319f $X=5.57 $Y=0.755
+ $X2=5.955 $Y2=1.37
cc_736 N_A_428_89#_c_1007_n N_A_808_115#_c_1391_n 0.00799344f $X=5.57 $Y=1.755
+ $X2=5.955 $Y2=1.37
cc_737 N_A_428_89#_c_1008_n N_A_808_115#_c_1391_n 0.0632121f $X=5.405 $Y=1.74
+ $X2=5.955 $Y2=1.37
cc_738 N_A_428_89#_c_1009_n N_A_808_115#_c_1391_n 0.0154865f $X=4.65 $Y=1.74
+ $X2=5.955 $Y2=1.37
cc_739 N_A_428_89#_c_1010_n N_A_808_115#_c_1391_n 0.0223158f $X=5.52 $Y=1.74
+ $X2=5.955 $Y2=1.37
cc_740 N_A_428_89#_c_993_n N_A_808_115#_c_1393_n 0.00133981f $X=4.37 $Y=1.825
+ $X2=4.48 $Y2=1.37
cc_741 N_A_428_89#_M1002_g N_A_808_115#_c_1393_n 9.98441e-19 $X=4.565 $Y=0.835
+ $X2=4.48 $Y2=1.37
cc_742 N_A_428_89#_c_1000_n N_A_808_115#_c_1393_n 0.00176044f $X=4.505 $Y=1.74
+ $X2=4.48 $Y2=1.37
cc_743 N_A_428_89#_c_1001_n N_A_808_115#_c_1393_n 0.00106749f $X=4.505 $Y=1.74
+ $X2=4.48 $Y2=1.37
cc_744 N_A_428_89#_c_1009_n N_A_808_115#_c_1393_n 0.012288f $X=4.65 $Y=1.74
+ $X2=4.48 $Y2=1.37
cc_745 N_A_428_89#_c_1002_n N_A_808_115#_c_1394_n 0.00257549f $X=5.57 $Y=0.755
+ $X2=6.1 $Y2=1.37
cc_746 N_A_970_89#_c_1198_n N_A_808_115#_M1004_g 0.0111108f $X=6.435 $Y=0.91
+ $X2=6.305 $Y2=0.755
cc_747 N_A_970_89#_c_1201_n N_A_808_115#_M1004_g 0.0118289f $X=6.52 $Y=1.625
+ $X2=6.305 $Y2=0.755
cc_748 N_A_970_89#_c_1204_n N_A_808_115#_M1004_g 5.28354e-19 $X=6.09 $Y=0.74
+ $X2=6.305 $Y2=0.755
cc_749 N_A_970_89#_c_1202_n N_A_808_115#_M1024_g 0.0187082f $X=6.52 $Y=3.615
+ $X2=6.305 $Y2=3.445
cc_750 N_A_970_89#_c_1207_n N_A_808_115#_M1024_g 0.00262846f $X=6.52 $Y=1.71
+ $X2=6.305 $Y2=3.445
cc_751 N_A_970_89#_c_1210_n N_A_808_115#_M1024_g 0.0144812f $X=5.882 $Y=2.39
+ $X2=6.305 $Y2=3.445
cc_752 N_A_970_89#_c_1211_n N_A_808_115#_M1024_g 0.0155115f $X=7.425 $Y=1.71
+ $X2=6.305 $Y2=3.445
cc_753 N_A_970_89#_c_1198_n N_A_808_115#_c_1382_n 0.00120425f $X=6.435 $Y=0.91
+ $X2=6.305 $Y2=1.37
cc_754 N_A_970_89#_c_1204_n N_A_808_115#_c_1382_n 0.00373221f $X=6.09 $Y=0.74
+ $X2=6.305 $Y2=1.37
cc_755 N_A_970_89#_c_1211_n N_A_808_115#_c_1382_n 0.0041429f $X=7.425 $Y=1.71
+ $X2=6.305 $Y2=1.37
cc_756 N_A_970_89#_c_1198_n N_A_808_115#_c_1385_n 0.00328408f $X=6.435 $Y=0.91
+ $X2=6.1 $Y2=1.37
cc_757 N_A_970_89#_c_1201_n N_A_808_115#_c_1385_n 0.0115453f $X=6.52 $Y=1.625
+ $X2=6.1 $Y2=1.37
cc_758 N_A_970_89#_c_1204_n N_A_808_115#_c_1385_n 0.0065907f $X=6.09 $Y=0.74
+ $X2=6.1 $Y2=1.37
cc_759 N_A_970_89#_c_1211_n N_A_808_115#_c_1385_n 7.75828e-19 $X=7.425 $Y=1.71
+ $X2=6.1 $Y2=1.37
cc_760 N_A_970_89#_c_1212_n N_A_808_115#_c_1385_n 0.0043276f $X=5.96 $Y=1.71
+ $X2=6.1 $Y2=1.37
cc_761 N_A_970_89#_M1006_g N_A_808_115#_c_1391_n 0.00582363f $X=4.925 $Y=0.835
+ $X2=5.955 $Y2=1.37
cc_762 N_A_970_89#_c_1185_n N_A_808_115#_c_1391_n 8.23686e-19 $X=4.985 $Y=1.71
+ $X2=5.955 $Y2=1.37
cc_763 N_A_970_89#_c_1197_n N_A_808_115#_c_1391_n 0.00523454f $X=4.985 $Y=1.71
+ $X2=5.955 $Y2=1.37
cc_764 N_A_970_89#_c_1212_n N_A_808_115#_c_1391_n 0.0148546f $X=5.96 $Y=1.71
+ $X2=5.955 $Y2=1.37
cc_765 N_A_970_89#_c_1198_n N_A_808_115#_c_1394_n 2.40329e-19 $X=6.435 $Y=0.91
+ $X2=6.1 $Y2=1.37
cc_766 N_A_970_89#_c_1201_n N_A_808_115#_c_1394_n 0.00353745f $X=6.52 $Y=1.625
+ $X2=6.1 $Y2=1.37
cc_767 N_A_970_89#_c_1204_n N_A_808_115#_c_1394_n 5.23046e-19 $X=6.09 $Y=0.74
+ $X2=6.1 $Y2=1.37
cc_768 N_A_970_89#_c_1212_n N_A_808_115#_c_1394_n 0.0291049f $X=5.96 $Y=1.71
+ $X2=6.1 $Y2=1.37
cc_769 N_A_970_89#_c_1188_n N_QN_M1027_g 0.0153129f $X=7.572 $Y=1.545 $X2=8.115
+ $Y2=0.835
cc_770 N_A_970_89#_c_1189_n N_QN_M1027_g 0.0210474f $X=7.66 $Y=1.17 $X2=8.115
+ $Y2=0.835
cc_771 N_A_970_89#_c_1203_n N_QN_M1027_g 4.79563e-19 $X=7.57 $Y=1.71 $X2=8.115
+ $Y2=0.835
cc_772 N_A_970_89#_c_1195_n N_QN_M1019_g 0.0102953f $X=7.66 $Y=2.375 $X2=8.115
+ $Y2=3.235
cc_773 N_A_970_89#_c_1196_n N_QN_M1019_g 0.0339596f $X=7.66 $Y=2.525 $X2=8.115
+ $Y2=3.235
cc_774 N_A_970_89#_c_1187_n N_QN_c_1527_n 0.021196f $X=7.57 $Y=1.71 $X2=8.055
+ $Y2=1.915
cc_775 N_A_970_89#_c_1203_n N_QN_c_1527_n 3.0115e-19 $X=7.57 $Y=1.71 $X2=8.055
+ $Y2=1.915
cc_776 N_A_970_89#_c_1213_n N_QN_c_1527_n 4.60229e-19 $X=7.57 $Y=1.71 $X2=8.055
+ $Y2=1.915
cc_777 N_A_970_89#_c_1189_n N_QN_c_1528_n 0.00439872f $X=7.66 $Y=1.17 $X2=7.47
+ $Y2=0.74
cc_778 N_A_970_89#_c_1194_n N_QN_c_1528_n 0.00327645f $X=7.66 $Y=1.32 $X2=7.47
+ $Y2=0.74
cc_779 N_A_970_89#_c_1195_n N_QN_c_1532_n 0.00567875f $X=7.66 $Y=2.375 $X2=7.47
+ $Y2=2.48
cc_780 N_A_970_89#_c_1196_n N_QN_c_1532_n 0.0128273f $X=7.66 $Y=2.525 $X2=7.47
+ $Y2=2.48
cc_781 N_A_970_89#_c_1188_n N_QN_c_1533_n 0.00749228f $X=7.572 $Y=1.545 $X2=7.97
+ $Y2=1.37
cc_782 N_A_970_89#_c_1194_n N_QN_c_1533_n 0.0108281f $X=7.66 $Y=1.32 $X2=7.97
+ $Y2=1.37
cc_783 N_A_970_89#_c_1203_n N_QN_c_1533_n 0.0110498f $X=7.57 $Y=1.71 $X2=7.97
+ $Y2=1.37
cc_784 N_A_970_89#_c_1213_n N_QN_c_1533_n 0.00387586f $X=7.57 $Y=1.71 $X2=7.97
+ $Y2=1.37
cc_785 N_A_970_89#_c_1187_n N_QN_c_1535_n 0.00308111f $X=7.57 $Y=1.71 $X2=7.555
+ $Y2=1.37
cc_786 N_A_970_89#_c_1203_n N_QN_c_1535_n 0.0120703f $X=7.57 $Y=1.71 $X2=7.555
+ $Y2=1.37
cc_787 N_A_970_89#_c_1211_n N_QN_c_1535_n 0.0010572f $X=7.425 $Y=1.71 $X2=7.555
+ $Y2=1.37
cc_788 N_A_970_89#_c_1213_n N_QN_c_1535_n 0.00336135f $X=7.57 $Y=1.71 $X2=7.555
+ $Y2=1.37
cc_789 N_A_970_89#_c_1195_n N_QN_c_1536_n 0.016126f $X=7.66 $Y=2.375 $X2=7.97
+ $Y2=2.285
cc_790 N_A_970_89#_c_1196_n N_QN_c_1536_n 0.00248624f $X=7.66 $Y=2.525 $X2=7.97
+ $Y2=2.285
cc_791 N_A_970_89#_c_1203_n N_QN_c_1536_n 0.00426371f $X=7.57 $Y=1.71 $X2=7.97
+ $Y2=2.285
cc_792 N_A_970_89#_c_1213_n N_QN_c_1536_n 0.00253233f $X=7.57 $Y=1.71 $X2=7.97
+ $Y2=2.285
cc_793 N_A_970_89#_c_1187_n N_QN_c_1537_n 0.00265611f $X=7.57 $Y=1.71 $X2=7.555
+ $Y2=2.285
cc_794 N_A_970_89#_c_1203_n N_QN_c_1537_n 0.00471962f $X=7.57 $Y=1.71 $X2=7.555
+ $Y2=2.285
cc_795 N_A_970_89#_c_1211_n N_QN_c_1537_n 9.40773e-19 $X=7.425 $Y=1.71 $X2=7.555
+ $Y2=2.285
cc_796 N_A_970_89#_c_1213_n N_QN_c_1537_n 0.00140341f $X=7.57 $Y=1.71 $X2=7.555
+ $Y2=2.285
cc_797 N_A_970_89#_c_1187_n N_QN_c_1538_n 0.00216137f $X=7.57 $Y=1.71 $X2=8.055
+ $Y2=1.915
cc_798 N_A_970_89#_c_1188_n N_QN_c_1538_n 0.00323473f $X=7.572 $Y=1.545
+ $X2=8.055 $Y2=1.915
cc_799 N_A_970_89#_c_1195_n N_QN_c_1538_n 0.00226435f $X=7.66 $Y=2.375 $X2=8.055
+ $Y2=1.915
cc_800 N_A_970_89#_c_1203_n N_QN_c_1538_n 0.00987106f $X=7.57 $Y=1.71 $X2=8.055
+ $Y2=1.915
cc_801 N_A_970_89#_c_1213_n N_QN_c_1538_n 0.00377439f $X=7.57 $Y=1.71 $X2=8.055
+ $Y2=1.915
cc_802 N_A_970_89#_c_1196_n QN 0.00740862f $X=7.66 $Y=2.525 $X2=7.475 $Y2=2.48
cc_803 N_A_970_89#_c_1202_n QN 0.00567439f $X=6.52 $Y=3.615 $X2=7.475 $Y2=2.48
cc_804 N_A_970_89#_c_1203_n QN 0.00350993f $X=7.57 $Y=1.71 $X2=7.475 $Y2=2.48
cc_805 N_A_970_89#_c_1213_n QN 0.00842298f $X=7.57 $Y=1.71 $X2=7.475 $Y2=2.48
cc_806 N_A_970_89#_c_1198_n A_1276_115# 0.00176584f $X=6.435 $Y=0.91 $X2=6.38
+ $Y2=0.575
cc_807 N_A_808_115#_c_1426_n A_736_521# 0.00342591f $X=4.095 $Y=2.705 $X2=3.68
+ $Y2=2.605
cc_808 N_A_808_115#_c_1459_n A_736_521# 0.00144354f $X=3.77 $Y=2.705 $X2=3.68
+ $Y2=2.605
cc_809 N_QN_M1019_g N_Q_c_1614_n 0.0038009f $X=8.115 $Y=3.235 $X2=8.33 $Y2=3.265
cc_810 N_QN_M1027_g N_Q_c_1612_n 0.0383548f $X=8.115 $Y=0.835 $X2=8.445 $Y2=2.68
cc_811 N_QN_c_1533_n N_Q_c_1612_n 0.0111776f $X=7.97 $Y=1.37 $X2=8.445 $Y2=2.68
cc_812 N_QN_c_1536_n N_Q_c_1612_n 0.0111776f $X=7.97 $Y=2.285 $X2=8.445 $Y2=2.68
cc_813 N_QN_c_1538_n N_Q_c_1612_n 0.0438362f $X=8.055 $Y=1.915 $X2=8.445
+ $Y2=2.68
cc_814 N_QN_M1027_g N_Q_c_1613_n 0.00373219f $X=8.115 $Y=0.835 $X2=8.445
+ $Y2=1.035
cc_815 N_QN_M1019_g N_Q_c_1618_n 0.00474029f $X=8.115 $Y=3.235 $X2=8.33
+ $Y2=2.807
cc_816 N_QN_M1019_g Q 0.0131514f $X=8.115 $Y=3.235 $X2=8.325 $Y2=2.85
cc_817 N_QN_c_1536_n Q 0.00245821f $X=7.97 $Y=2.285 $X2=8.325 $Y2=2.85
