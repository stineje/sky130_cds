* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_18T_hs__buf_4
** N=7 EP=0 IP=0 FDC=13
M0 gnd A 4 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=575 $D=19
M1 Y 4 gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=575 $D=19
M2 gnd 4 Y gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=575 $D=19
M3 Y 4 gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=575 $D=19
M4 gnd 4 Y gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2120 $Y=575 $D=19
M5 vdd A 4 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=400 $Y=3085 $D=79
M6 Y 4 vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=830 $Y=3085 $D=79
M7 vdd 4 Y vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=1260 $Y=3085 $D=79
M8 Y 4 vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=1690 $Y=3085 $D=79
M9 vdd 4 Y vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=2120 $Y=3085 $D=79
X10 gnd vdd Dpar a=10.659 p=13.21 m=1 $[nwdiode] $X=-45 $Y=2905 $D=185
X11 6 A Probe probetype=1 $[A] $X=633 $Y=3328 $D=289
X12 7 Y Probe probetype=1 $[Y] $X=1053 $Y=2268 $D=289
.ENDS
***************************************
