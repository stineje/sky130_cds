magic
tech sky130A
magscale 1 2
timestamp 1640011036
<< nwell >>
rect 0 1336 255 1337
rect -269 763 1317 1336
rect -269 576 1310 763
<< nmoslvt >>
rect -180 110 -150 310
rect -94 110 -64 310
rect 96 110 126 310
rect 182 110 212 310
rect 254 110 284 310
rect 374 110 404 310
rect 446 110 476 310
rect 532 110 562 310
rect 740 110 770 310
rect 826 110 856 310
rect 1016 110 1046 310
rect 1102 110 1132 310
rect 1188 110 1218 310
<< pmos >>
rect -180 612 -150 1212
rect -108 612 -78 1212
rect 96 612 126 1212
rect 182 612 212 1212
rect 254 612 284 1212
rect 374 612 404 1212
rect 446 612 476 1212
rect 532 612 562 1212
rect 740 612 770 1212
rect 826 612 856 1212
rect 1016 612 1046 1212
rect 1102 612 1132 1212
rect 1188 612 1218 1212
<< ndiff >>
rect -233 262 -180 310
rect -233 126 -225 262
rect -191 126 -180 262
rect -233 110 -180 126
rect -150 262 -94 310
rect -150 126 -139 262
rect -105 126 -94 262
rect -150 110 -94 126
rect -64 262 -11 310
rect -64 126 -53 262
rect -19 126 -11 262
rect -64 110 -11 126
rect 43 262 96 310
rect 43 126 51 262
rect 85 126 96 262
rect 43 110 96 126
rect 126 262 182 310
rect 126 126 137 262
rect 171 126 182 262
rect 126 110 182 126
rect 212 110 254 310
rect 284 262 374 310
rect 284 126 295 262
rect 363 126 374 262
rect 284 110 374 126
rect 404 110 446 310
rect 476 262 532 310
rect 476 126 487 262
rect 521 126 532 262
rect 476 110 532 126
rect 562 262 615 310
rect 562 126 573 262
rect 607 126 615 262
rect 562 110 615 126
rect 687 262 740 310
rect 687 126 695 262
rect 729 126 740 262
rect 687 110 740 126
rect 770 262 826 310
rect 770 126 781 262
rect 815 126 826 262
rect 770 110 826 126
rect 856 262 909 310
rect 856 126 867 262
rect 901 126 909 262
rect 856 110 909 126
rect 963 262 1016 310
rect 963 126 971 262
rect 1005 126 1016 262
rect 963 110 1016 126
rect 1046 262 1102 310
rect 1046 126 1057 262
rect 1091 126 1102 262
rect 1046 110 1102 126
rect 1132 262 1188 310
rect 1132 126 1143 262
rect 1177 126 1188 262
rect 1132 110 1188 126
rect 1218 262 1271 310
rect 1218 126 1229 262
rect 1263 126 1271 262
rect 1218 110 1271 126
<< pdiff >>
rect -233 1196 -180 1212
rect -233 652 -225 1196
rect -191 652 -180 1196
rect -233 612 -180 652
rect -150 612 -108 1212
rect -78 1196 -25 1212
rect -78 788 -67 1196
rect -33 788 -25 1196
rect -78 612 -25 788
rect 43 1196 96 1212
rect 43 720 51 1196
rect 85 720 96 1196
rect 43 612 96 720
rect 126 1196 182 1212
rect 126 720 137 1196
rect 171 720 182 1196
rect 126 612 182 720
rect 212 612 254 1212
rect 284 1196 374 1212
rect 284 652 295 1196
rect 363 652 374 1196
rect 284 612 374 652
rect 404 612 446 1212
rect 476 1196 532 1212
rect 476 652 487 1196
rect 521 652 532 1196
rect 476 612 532 652
rect 562 1196 615 1212
rect 562 652 573 1196
rect 607 652 615 1196
rect 562 612 615 652
rect 687 1196 740 1212
rect 687 652 695 1196
rect 729 652 740 1196
rect 687 612 740 652
rect 770 1196 826 1212
rect 770 652 781 1196
rect 815 652 826 1196
rect 770 612 826 652
rect 856 1196 909 1212
rect 856 652 867 1196
rect 901 652 909 1196
rect 856 612 909 652
rect 963 1196 1016 1212
rect 963 720 971 1196
rect 1005 720 1016 1196
rect 963 612 1016 720
rect 1046 612 1102 1212
rect 1132 1196 1188 1212
rect 1132 788 1143 1196
rect 1177 788 1188 1196
rect 1132 612 1188 788
rect 1218 1196 1271 1212
rect 1218 652 1229 1196
rect 1263 652 1271 1196
rect 1218 612 1271 652
<< ndiffc >>
rect -225 126 -191 262
rect -139 126 -105 262
rect -53 126 -19 262
rect 51 126 85 262
rect 137 126 171 262
rect 295 126 363 262
rect 487 126 521 262
rect 573 126 607 262
rect 695 126 729 262
rect 781 126 815 262
rect 867 126 901 262
rect 971 126 1005 262
rect 1057 126 1091 262
rect 1143 126 1177 262
rect 1229 126 1263 262
<< pdiffc >>
rect -225 652 -191 1196
rect -67 788 -33 1196
rect 51 720 85 1196
rect 137 720 171 1196
rect 295 652 363 1196
rect 487 652 521 1196
rect 573 652 607 1196
rect 695 652 729 1196
rect 781 652 815 1196
rect 867 652 901 1196
rect 971 720 1005 1196
rect 1143 788 1177 1196
rect 1229 652 1263 1196
<< psubdiff >>
rect -233 22 -209 56
rect -175 22 -151 56
rect -97 22 -73 56
rect -39 22 -15 56
rect 88 22 112 56
rect 146 22 170 56
rect 224 22 248 56
rect 282 22 306 56
rect 360 22 384 56
rect 418 22 442 56
rect 496 22 520 56
rect 554 22 578 56
rect 632 22 656 56
rect 690 22 714 56
rect 768 22 792 56
rect 826 22 850 56
rect 963 22 987 56
rect 1021 22 1045 56
rect 1099 22 1123 56
rect 1157 22 1181 56
<< nsubdiff >>
rect -233 1266 -209 1300
rect -175 1266 -151 1300
rect -97 1266 -73 1300
rect -39 1266 -15 1300
rect 88 1266 112 1300
rect 146 1266 170 1300
rect 224 1266 248 1300
rect 282 1266 306 1300
rect 360 1266 384 1300
rect 418 1266 442 1300
rect 496 1266 520 1300
rect 554 1266 578 1300
rect 632 1266 656 1300
rect 690 1266 714 1300
rect 768 1266 792 1300
rect 826 1266 850 1300
rect 963 1266 987 1300
rect 1021 1266 1045 1300
rect 1099 1266 1123 1300
rect 1157 1266 1181 1300
<< psubdiffcont >>
rect -209 22 -175 56
rect -73 22 -39 56
rect 112 22 146 56
rect 248 22 282 56
rect 384 22 418 56
rect 520 22 554 56
rect 656 22 690 56
rect 792 22 826 56
rect 987 22 1021 56
rect 1123 22 1157 56
<< nsubdiffcont >>
rect -209 1266 -175 1300
rect -73 1266 -39 1300
rect 112 1266 146 1300
rect 248 1266 282 1300
rect 384 1266 418 1300
rect 520 1266 554 1300
rect 656 1266 690 1300
rect 792 1266 826 1300
rect 987 1266 1021 1300
rect 1123 1266 1157 1300
<< poly >>
rect -180 1212 -150 1238
rect -108 1212 -78 1238
rect 96 1212 126 1238
rect 182 1212 212 1238
rect 254 1212 284 1238
rect 374 1212 404 1238
rect 446 1212 476 1238
rect 532 1212 562 1238
rect 740 1212 770 1238
rect 826 1212 856 1238
rect 1016 1212 1046 1238
rect 1102 1212 1132 1238
rect 1188 1212 1218 1238
rect -180 446 -150 612
rect -108 579 -78 612
rect 96 590 126 612
rect -108 563 -35 579
rect -108 529 -79 563
rect -45 529 -35 563
rect -108 513 -35 529
rect 86 556 126 590
rect -204 430 -150 446
rect -204 396 -194 430
rect -160 396 -150 430
rect -204 380 -150 396
rect -180 310 -150 380
rect -94 310 -64 513
rect 86 398 116 556
rect 182 513 212 612
rect 254 581 284 612
rect 374 581 404 612
rect 254 565 308 581
rect 254 531 264 565
rect 298 531 308 565
rect 254 515 308 531
rect 350 565 404 581
rect 350 531 360 565
rect 394 531 404 565
rect 350 515 404 531
rect 158 497 212 513
rect 158 463 168 497
rect 202 463 212 497
rect 350 470 380 515
rect 158 447 212 463
rect 86 382 140 398
rect 86 348 96 382
rect 130 348 140 382
rect 86 332 140 348
rect 96 310 126 332
rect 182 310 212 447
rect 254 440 380 470
rect 446 472 476 612
rect 532 581 562 612
rect 740 596 770 612
rect 532 565 603 581
rect 532 551 559 565
rect 543 531 559 551
rect 593 531 603 565
rect 543 515 603 531
rect 730 566 770 596
rect 446 456 500 472
rect 254 310 284 440
rect 446 422 456 456
rect 490 422 500 456
rect 446 406 500 422
rect 350 382 404 398
rect 350 348 360 382
rect 394 348 404 382
rect 350 332 404 348
rect 374 310 404 332
rect 446 310 476 406
rect 543 358 573 515
rect 730 472 760 566
rect 826 472 856 612
rect 1016 563 1046 612
rect 963 547 1046 563
rect 963 513 973 547
rect 1007 513 1046 547
rect 963 497 1046 513
rect 1102 505 1132 612
rect 1188 587 1218 612
rect 1188 557 1225 587
rect 705 456 760 472
rect 705 422 715 456
rect 749 422 760 456
rect 705 406 760 422
rect 802 456 856 472
rect 802 422 812 456
rect 846 422 856 456
rect 802 406 856 422
rect 532 328 573 358
rect 730 355 760 406
rect 532 310 562 328
rect 730 325 770 355
rect 740 310 770 325
rect 826 310 856 406
rect 1016 310 1046 497
rect 1099 489 1153 505
rect 1099 455 1109 489
rect 1143 455 1153 489
rect 1099 439 1153 455
rect 1102 310 1132 439
rect 1195 415 1225 557
rect 1195 399 1249 415
rect 1195 379 1205 399
rect 1188 365 1205 379
rect 1239 365 1249 399
rect 1188 349 1249 365
rect 1188 310 1218 349
rect -180 84 -150 110
rect -94 84 -64 110
rect 96 84 126 110
rect 182 84 212 110
rect 254 84 284 110
rect 374 84 404 110
rect 446 84 476 110
rect 532 84 562 110
rect 740 84 770 110
rect 826 84 856 110
rect 1016 84 1046 110
rect 1102 84 1132 110
rect 1188 84 1218 110
<< polycont >>
rect -79 529 -45 563
rect -194 396 -160 430
rect 264 531 298 565
rect 360 531 394 565
rect 168 463 202 497
rect 96 348 130 382
rect 559 531 593 565
rect 456 422 490 456
rect 360 348 394 382
rect 973 513 1007 547
rect 715 422 749 456
rect 812 422 846 456
rect 1109 455 1143 489
rect 1205 365 1239 399
<< locali >>
rect -267 1306 1317 1327
rect -267 1266 -209 1306
rect -175 1266 -73 1306
rect -39 1266 112 1306
rect 146 1266 248 1306
rect 282 1266 384 1306
rect 418 1266 520 1306
rect 554 1266 656 1306
rect 690 1266 792 1306
rect 826 1266 987 1306
rect 1021 1266 1123 1306
rect 1157 1266 1317 1306
rect -225 1196 -191 1212
rect -67 1196 -33 1266
rect -67 772 -33 788
rect 51 1196 85 1212
rect 28 720 51 786
rect 28 703 85 720
rect 137 1196 171 1266
rect 137 704 171 720
rect 295 1196 363 1212
rect -225 530 -191 652
rect -147 430 -113 570
rect -79 563 -45 644
rect -79 513 -45 529
rect -210 396 -194 430
rect -160 396 -113 430
rect 28 456 62 703
rect 295 649 363 652
rect -225 262 -191 278
rect -225 56 -191 126
rect 28 291 62 422
rect 96 615 363 649
rect 487 1196 521 1266
rect 487 636 521 652
rect 573 1196 607 1212
rect 573 649 607 652
rect 695 1196 729 1212
rect 573 615 661 649
rect 96 382 130 615
rect 360 565 394 581
rect 248 531 264 565
rect 298 531 314 565
rect 168 447 202 463
rect 280 382 314 531
rect 360 530 394 531
rect 559 565 593 581
rect 559 530 593 531
rect 627 456 661 615
rect 695 604 729 652
rect 781 1196 815 1266
rect 781 636 815 652
rect 867 1196 901 1212
rect 971 1196 1005 1212
rect 1143 1196 1177 1266
rect 1143 772 1177 788
rect 1229 1196 1263 1212
rect 1005 720 1075 738
rect 971 704 1075 720
rect 901 644 914 661
rect 867 627 914 644
rect 695 565 729 570
rect 695 531 846 565
rect 812 456 846 531
rect 440 422 456 456
rect 490 422 506 456
rect 573 422 661 456
rect 699 422 715 456
rect 749 422 765 456
rect 573 382 607 422
rect 812 382 846 422
rect 130 348 239 382
rect 280 348 360 382
rect 394 348 607 382
rect 96 332 130 348
rect 205 298 239 348
rect -139 262 -105 274
rect -139 110 -105 126
rect -53 262 -19 278
rect 28 262 85 291
rect 28 257 51 262
rect -53 56 -19 126
rect 51 110 85 126
rect 137 262 171 278
rect 205 264 363 298
rect 137 56 171 126
rect 295 262 363 264
rect 295 110 363 126
rect 487 262 521 278
rect 487 56 521 126
rect 573 262 607 348
rect 573 110 607 126
rect 695 348 846 382
rect 695 262 729 348
rect 880 314 914 627
rect 973 547 1007 570
rect 973 497 1007 513
rect 1041 399 1075 704
rect 1109 530 1143 644
rect 1229 530 1263 652
rect 1109 489 1143 496
rect 1109 439 1143 455
rect 1041 365 1205 399
rect 1239 365 1255 399
rect 867 280 914 314
rect 695 110 729 126
rect 781 262 815 278
rect 781 56 815 126
rect 867 262 901 280
rect 867 110 901 126
rect 971 262 1005 278
rect 971 56 1005 126
rect 1057 262 1091 365
rect 1057 110 1091 126
rect 1143 262 1177 278
rect 1143 56 1177 126
rect 1229 262 1263 274
rect 1229 110 1263 126
rect -267 16 -209 56
rect -175 16 -73 56
rect -39 16 112 56
rect 146 16 248 56
rect 282 16 384 56
rect 418 16 520 56
rect 554 16 656 56
rect 690 16 792 56
rect 826 16 987 56
rect 1021 16 1123 56
rect 1157 16 1317 56
rect -267 -5 1317 16
<< viali >>
rect -209 1300 -175 1306
rect -209 1272 -175 1300
rect -73 1300 -39 1306
rect -73 1272 -39 1300
rect 112 1300 146 1306
rect 112 1272 146 1300
rect 248 1300 282 1306
rect 248 1272 282 1300
rect 384 1300 418 1306
rect 384 1272 418 1300
rect 520 1300 554 1306
rect 520 1272 554 1300
rect 656 1300 690 1306
rect 656 1272 690 1300
rect 792 1300 826 1306
rect 792 1272 826 1300
rect 987 1300 1021 1306
rect 987 1272 1021 1300
rect 1123 1300 1157 1306
rect 1123 1272 1157 1300
rect -79 644 -45 678
rect -225 496 -191 530
rect -147 570 -113 604
rect 28 422 62 456
rect -139 274 -105 308
rect 168 497 202 531
rect 360 496 394 530
rect 559 496 593 530
rect 867 652 901 678
rect 867 644 901 652
rect 695 570 729 604
rect 456 422 490 456
rect 715 422 749 456
rect 973 570 1007 604
rect 1109 644 1143 678
rect 1109 496 1143 530
rect 1229 496 1263 530
rect 1229 274 1263 308
rect -209 22 -175 50
rect -209 16 -175 22
rect -73 22 -39 50
rect -73 16 -39 22
rect 112 22 146 50
rect 112 16 146 22
rect 248 22 282 50
rect 248 16 282 22
rect 384 22 418 50
rect 384 16 418 22
rect 520 22 554 50
rect 520 16 554 22
rect 656 22 690 50
rect 656 16 690 22
rect 792 22 826 50
rect 792 16 826 22
rect 987 22 1021 50
rect 987 16 1021 22
rect 1123 22 1157 50
rect 1123 16 1157 22
<< metal1 >>
rect -267 1306 1317 1327
rect -267 1272 -209 1306
rect -175 1272 -73 1306
rect -39 1272 112 1306
rect 146 1272 248 1306
rect 282 1272 384 1306
rect 418 1272 520 1306
rect 554 1272 656 1306
rect 690 1272 792 1306
rect 826 1272 987 1306
rect 1021 1272 1123 1306
rect 1157 1272 1317 1306
rect -267 1266 1317 1272
rect -91 678 -33 684
rect 855 678 913 684
rect 1097 678 1155 684
rect -112 644 -79 678
rect -45 644 -33 678
rect 832 644 867 678
rect 901 644 913 678
rect 1076 644 1109 678
rect 1143 644 1155 678
rect -91 638 -33 644
rect 855 638 913 644
rect 1097 638 1155 644
rect -159 604 -101 610
rect 683 604 741 610
rect 961 604 1019 610
rect -181 570 -147 604
rect -113 570 -101 604
rect 676 603 695 604
rect 661 571 695 603
rect 676 570 695 571
rect 729 570 973 604
rect 1007 570 1041 604
rect -159 564 -101 570
rect 683 564 741 570
rect 961 564 1019 570
rect -237 530 -179 536
rect 156 531 215 537
rect 156 530 168 531
rect -237 496 -225 530
rect -191 497 168 530
rect 202 497 235 531
rect 348 530 406 536
rect 547 530 605 536
rect 1097 530 1155 536
rect -191 496 215 497
rect -237 490 -179 496
rect -139 314 -105 496
rect 156 491 215 496
rect 348 496 360 530
rect 394 496 559 530
rect 593 496 1109 530
rect 1143 496 1155 530
rect 348 490 406 496
rect 547 490 605 496
rect 1097 490 1155 496
rect 1217 530 1275 536
rect 1217 496 1229 530
rect 1263 496 1275 530
rect 1217 490 1275 496
rect 15 456 74 462
rect 15 422 28 456
rect 62 449 74 456
rect 444 456 503 462
rect 444 449 456 456
rect 62 422 456 449
rect 490 453 503 456
rect 703 456 761 462
rect 703 453 715 456
rect 490 425 715 453
rect 490 422 503 425
rect 15 421 503 422
rect 15 416 74 421
rect 444 416 503 421
rect 703 422 715 425
rect 749 422 761 456
rect 703 416 761 422
rect 1229 314 1263 490
rect -151 308 -93 314
rect -151 274 -139 308
rect -105 274 -93 308
rect -151 268 -93 274
rect 1217 308 1275 314
rect 1217 274 1229 308
rect 1263 274 1275 308
rect 1217 268 1275 274
rect -267 50 1317 56
rect -267 16 -209 50
rect -175 16 -73 50
rect -39 16 112 50
rect 146 16 248 50
rect 282 16 384 50
rect 418 16 520 50
rect 554 16 656 50
rect 690 16 792 50
rect 826 16 987 50
rect 1021 16 1123 50
rect 1157 16 1317 50
rect -267 -5 1317 16
<< labels >>
rlabel viali -130 587 -130 587 1 SE
rlabel viali -61 660 -61 660 1 E
rlabel viali 576 513 576 513 1 CK
rlabel viali 1246 513 1246 513 1 ECK
rlabel viali -192 36 -192 36 1 gnd
rlabel viali -56 34 -56 34 1 gnd
rlabel viali 129 34 129 34 1 gnd
rlabel viali 265 34 265 34 1 gnd
rlabel viali 400 35 400 35 1 gnd
rlabel viali 536 33 536 33 1 gnd
rlabel viali 673 33 673 33 1 gnd
rlabel viali 810 34 810 34 1 gnd
rlabel viali 1005 34 1005 34 1 gnd
rlabel viali 1139 35 1139 35 1 gnd
rlabel nwell -191 1287 -190 1287 1 vdd
rlabel nwell -56 1288 -55 1288 1 vdd
rlabel nwell 129 1288 130 1288 1 vdd
rlabel viali 264 1287 264 1287 1 vdd
rlabel viali 401 1289 401 1289 1 vdd
rlabel viali 538 1289 538 1289 1 vdd
rlabel nwell 674 1289 674 1290 1 vdd
rlabel nwell 809 1290 809 1291 1 vdd
rlabel nwell 1004 1289 1004 1290 1 vdd
rlabel nwell 1141 1289 1141 1290 1 vdd
<< end >>
