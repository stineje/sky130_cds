magic
tech sky130A
magscale 1 2
timestamp 1606864607
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 286 1341
<< nmos >>
rect 80 115 110 315
rect 166 115 196 315
<< pmos >>
rect 80 617 110 1217
rect 152 617 182 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 166 315
rect 110 131 121 267
rect 155 131 166 267
rect 110 115 166 131
rect 196 267 249 315
rect 196 131 207 267
rect 241 131 249 267
rect 196 115 249 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 657 35 1201
rect 69 657 80 1201
rect 27 617 80 657
rect 110 617 152 1217
rect 182 1201 235 1217
rect 182 793 193 1201
rect 227 793 235 1201
rect 182 617 235 793
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 207 131 241 267
<< pdiffc >>
rect 35 657 69 1201
rect 193 793 227 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 152 1217 182 1243
rect 80 451 110 617
rect 152 584 182 617
rect 152 568 225 584
rect 152 534 181 568
rect 215 534 225 568
rect 152 518 225 534
rect 56 435 110 451
rect 56 401 66 435
rect 100 401 110 435
rect 56 385 110 401
rect 80 315 110 385
rect 166 315 196 518
rect 80 89 110 115
rect 166 89 196 115
<< polycont >>
rect 181 534 215 568
rect 66 401 100 435
<< locali >>
rect 0 1311 286 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 286 1311
rect 35 1201 69 1217
rect 193 1201 227 1271
rect 193 777 227 793
rect 35 535 69 657
rect 113 435 147 575
rect 181 568 215 649
rect 181 518 215 534
rect 50 401 66 435
rect 100 401 147 435
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 279
rect 121 115 155 131
rect 207 267 241 283
rect 207 61 241 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 181 649 215 683
rect 35 501 69 535
rect 113 575 147 609
rect 121 279 155 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 286 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 286 1311
rect 0 1271 286 1277
rect 169 683 227 689
rect 148 649 181 683
rect 215 649 227 683
rect 169 643 227 649
rect 101 609 159 615
rect 79 575 113 609
rect 147 575 159 609
rect 101 569 159 575
rect 23 535 81 541
rect 23 501 35 535
rect 69 501 155 535
rect 23 495 81 501
rect 121 319 155 501
rect 109 313 167 319
rect 109 279 121 313
rect 155 279 167 313
rect 109 273 167 279
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 137 393 137 393 1 Y
port 1 n
rlabel metal1 130 592 130 592 1 B
port 2 n
rlabel metal1 198 666 198 666 1 A
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
