* File: sky130_osu_sc_18T_hs__dffr_1.pex.spice
* Created: Fri Nov 12 13:48:58 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%GND 1 2 3 4 5 6 7 8 9 121 125 127 134
+ 136 143 152 154 164 166 176 178 185 187 194 196 203 230 232
c221 176 0 1.67294e-19 $X=6.09 $Y=0.825
c222 152 0 3.07193e-19 $X=2.59 $Y=0.825
c223 121 0 1.27355e-19 $X=-0.05 $Y=0
r224 230 232 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.175 $Y2=0.152
r225 205 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.152
+ $X2=8.85 $Y2=0.152
r226 201 226 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.152
r227 201 203 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.825
r228 196 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.152
+ $X2=8.85 $Y2=0.152
r229 192 194 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.825
r230 188 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.152
+ $X2=7.04 $Y2=0.152
r231 183 222 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.152
r232 183 185 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.825
r233 179 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.152
+ $X2=6.09 $Y2=0.152
r234 178 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.152
+ $X2=7.04 $Y2=0.152
r235 174 221 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.152
r236 174 176 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.825
r237 166 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.152
+ $X2=6.09 $Y2=0.152
r238 162 164 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.34 $Y=0.305
+ $X2=4.34 $Y2=0.825
r239 155 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.152
+ $X2=2.59 $Y2=0.152
r240 150 217 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.152
r241 150 152 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.825
r242 146 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.152
+ $X2=2.07 $Y2=0.152
r243 145 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.152
+ $X2=2.59 $Y2=0.152
r244 141 216 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.152
r245 141 143 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.825
r246 137 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.152
+ $X2=1.21 $Y2=0.152
r247 136 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.152
+ $X2=2.07 $Y2=0.152
r248 132 215 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.152
r249 132 134 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.825
r250 127 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.152
+ $X2=1.21 $Y2=0.152
r251 123 125 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r252 121 232 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=0.19 $X2=9.175 $Y2=0.19
r253 121 230 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=0.19 $X2=0.335 $Y2=0.19
r254 121 192 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r255 121 187 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r256 121 197 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.985 $Y2=0.152
r257 121 162 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.34 $Y2=0.305
r258 121 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.255 $Y2=0.152
r259 121 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.425 $Y2=0.152
r260 121 123 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r261 121 128 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r262 121 205 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.935 $Y2=0.152
r263 121 196 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.765 $Y2=0.152
r264 121 197 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=7.985 $Y2=0.152
r265 121 187 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r266 121 188 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.125 $Y2=0.152
r267 121 178 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.955 $Y2=0.152
r268 121 179 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.175 $Y2=0.152
r269 121 166 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.005 $Y2=0.152
r270 121 167 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.425 $Y2=0.152
r271 121 154 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=4.255 $Y2=0.152
r272 121 155 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=2.675 $Y2=0.152
r273 121 145 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.505 $Y2=0.152
r274 121 146 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.155 $Y2=0.152
r275 121 136 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.985 $Y2=0.152
r276 121 137 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.295 $Y2=0.152
r277 121 127 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.125 $Y2=0.152
r278 121 128 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r279 9 203 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.575 $X2=8.85 $Y2=0.825
r280 8 194 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.825
r281 7 185 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.575 $X2=7.04 $Y2=0.825
r282 6 176 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.95
+ $Y=0.575 $X2=6.09 $Y2=0.825
r283 5 164 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.575 $X2=4.34 $Y2=0.825
r284 4 152 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=2.465
+ $Y=0.575 $X2=2.59 $Y2=0.825
r285 3 143 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.825
r286 2 134 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.825
r287 1 125 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%VDD 1 2 3 4 5 6 7 85 89 93 101 111 115
+ 123 127 135 139 147 151 157 163 178 182
r117 178 182 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=6.507
+ $X2=9.175 $Y2=6.507
r118 167 178 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=6.47 $X2=0.335 $Y2=6.47
r119 163 182 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=6.47 $X2=9.175 $Y2=6.47
r120 161 176 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=6.507
+ $X2=8.85 $Y2=6.507
r121 161 163 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=8.935 $Y=6.507
+ $X2=9.175 $Y2=6.507
r122 157 160 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=8.85 $Y=4.475
+ $X2=8.85 $Y2=5.835
r123 155 176 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.85 $Y=6.355
+ $X2=8.85 $Y2=6.507
r124 155 160 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.85 $Y=6.355
+ $X2=8.85 $Y2=5.835
r125 152 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=6.507
+ $X2=7.83 $Y2=6.507
r126 152 154 21.9153 $w=3.03e-07 $l=5.8e-07 $layer=LI1_cond $X=7.915 $Y=6.507
+ $X2=8.495 $Y2=6.507
r127 151 176 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=6.507
+ $X2=8.85 $Y2=6.507
r128 151 154 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.765 $Y=6.507
+ $X2=8.495 $Y2=6.507
r129 147 150 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.83 $Y=4.475
+ $X2=7.83 $Y2=5.835
r130 145 175 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.83 $Y=6.355
+ $X2=7.83 $Y2=6.507
r131 145 150 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.83 $Y=6.355
+ $X2=7.83 $Y2=5.835
r132 142 144 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.455 $Y=6.507
+ $X2=7.135 $Y2=6.507
r133 140 173 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.09 $Y2=6.507
r134 140 142 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.455 $Y2=6.507
r135 139 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=6.507
+ $X2=7.83 $Y2=6.507
r136 139 144 23.0489 $w=3.03e-07 $l=6.1e-07 $layer=LI1_cond $X=7.745 $Y=6.507
+ $X2=7.135 $Y2=6.507
r137 135 138 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.09 $Y=3.455
+ $X2=6.09 $Y2=5.835
r138 133 173 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=6.507
r139 133 138 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=5.835
r140 130 132 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=6.507
+ $X2=5.775 $Y2=6.507
r141 128 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=6.507
+ $X2=4.34 $Y2=6.507
r142 128 130 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.425 $Y=6.507
+ $X2=5.095 $Y2=6.507
r143 127 173 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=6.09 $Y2=6.507
r144 127 132 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=5.775 $Y2=6.507
r145 123 126 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.34 $Y=3.795
+ $X2=4.34 $Y2=5.835
r146 121 172 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.34 $Y=6.355
+ $X2=4.34 $Y2=6.507
r147 121 126 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.34 $Y=6.355
+ $X2=4.34 $Y2=5.835
r148 118 120 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=6.507
+ $X2=3.735 $Y2=6.507
r149 116 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=6.507
+ $X2=2.59 $Y2=6.507
r150 116 118 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.675 $Y=6.507
+ $X2=3.055 $Y2=6.507
r151 115 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=6.507
+ $X2=4.34 $Y2=6.507
r152 115 120 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=4.255 $Y=6.507
+ $X2=3.735 $Y2=6.507
r153 111 114 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.59 $Y=3.795
+ $X2=2.59 $Y2=5.835
r154 109 170 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.59 $Y=6.355
+ $X2=2.59 $Y2=6.507
r155 109 114 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.59 $Y=6.355
+ $X2=2.59 $Y2=5.835
r156 106 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=6.507
+ $X2=2 $Y2=6.507
r157 106 108 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=2.085 $Y=6.507
+ $X2=2.375 $Y2=6.507
r158 105 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=6.507
+ $X2=2.59 $Y2=6.507
r159 105 108 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=6.507
+ $X2=2.375 $Y2=6.507
r160 101 104 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2 $Y=4.475 $X2=2
+ $Y2=5.835
r161 99 169 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2 $Y=6.355 $X2=2
+ $Y2=6.507
r162 99 104 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2 $Y=6.355 $X2=2
+ $Y2=5.835
r163 96 98 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=6.507
+ $X2=1.695 $Y2=6.507
r164 94 167 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r165 94 96 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.015 $Y2=6.507
r166 93 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=6.507
+ $X2=2 $Y2=6.507
r167 93 98 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.915 $Y=6.507
+ $X2=1.695 $Y2=6.507
r168 89 92 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r169 87 167 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r170 87 92 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r171 85 163 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=6.355 $X2=9.175 $Y2=6.44
r172 85 154 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=6.355 $X2=8.495 $Y2=6.44
r173 85 175 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=6.355 $X2=7.815 $Y2=6.44
r174 85 144 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=6.355 $X2=7.135 $Y2=6.44
r175 85 142 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=6.355 $X2=6.455 $Y2=6.44
r176 85 132 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=6.355 $X2=5.775 $Y2=6.44
r177 85 130 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=6.355 $X2=5.095 $Y2=6.44
r178 85 172 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=6.355 $X2=4.415 $Y2=6.44
r179 85 120 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=6.355 $X2=3.735 $Y2=6.44
r180 85 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=6.355 $X2=3.055 $Y2=6.44
r181 85 108 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=6.355 $X2=2.375 $Y2=6.44
r182 85 98 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=6.355 $X2=1.695 $Y2=6.44
r183 85 96 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=6.355 $X2=1.015 $Y2=6.44
r184 85 167 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=6.355 $X2=0.335 $Y2=6.44
r185 7 160 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=3.085 $X2=8.85 $Y2=5.835
r186 7 157 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=3.085 $X2=8.85 $Y2=4.475
r187 6 150 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=4.085 $X2=7.83 $Y2=5.835
r188 6 147 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=4.085 $X2=7.83 $Y2=4.475
r189 5 138 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5.95
+ $Y=3.085 $X2=6.09 $Y2=5.835
r190 5 135 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5.95
+ $Y=3.085 $X2=6.09 $Y2=3.455
r191 4 126 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=4.2
+ $Y=3.085 $X2=4.34 $Y2=5.835
r192 4 123 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=4.2
+ $Y=3.085 $X2=4.34 $Y2=3.795
r193 3 114 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=2.465 $Y=3.085 $X2=2.59 $Y2=5.835
r194 3 111 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=2.465 $Y=3.085 $X2=2.59 $Y2=3.795
r195 2 104 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=4.085 $X2=2 $Y2=5.835
r196 2 101 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=4.085 $X2=2 $Y2=4.475
r197 1 92 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r198 1 89 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%RN 3 5 7 13 15 21
c38 21 0 7.48684e-20 $X=0.325 $Y=3.33
c39 3 0 1.0751e-19 $X=0.475 $Y=1.075
r40 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=3.33
+ $X2=0.325 $Y2=3.33
r41 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=2.305
+ $X2=0.53 $Y2=2.305
r42 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r43 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.47
+ $X2=0.32 $Y2=2.305
r44 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=2.47 $X2=0.32
+ $Y2=3.33
r45 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=2.305 $X2=0.53 $Y2=2.305
r46 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.53 $Y2=2.305
r47 5 7 1084.5 $w=1.5e-07 $l=2.115e-06 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=4.585
r48 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.53 $Y2=2.305
r49 1 3 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_110_115# 1 3 9 11 14 18 20 22 26 32 36
+ 40 45 46 47 49 59 62 67 68 73
c173 68 0 1.63751e-20 $X=1.375 $Y=1.48
c174 62 0 9.11346e-20 $X=1.23 $Y=1.48
c175 59 0 7.48684e-20 $X=0.87 $Y=2.74
c176 18 0 1.88625e-19 $X=7.615 $Y=5.085
r177 68 70 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.375 $Y=1.48
+ $X2=1.23 $Y2=1.48
r178 67 73 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.665 $Y=1.48
+ $X2=7.81 $Y2=1.48
r179 67 68 6.05653 $w=1.7e-07 $l=6.29e-06 $layer=MET1_cond $X=7.665 $Y=1.48
+ $X2=1.375 $Y2=1.48
r180 62 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.48
+ $X2=1.23 $Y2=1.48
r181 62 65 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.23 $Y=1.48
+ $X2=1.23 $Y2=1.59
r182 57 59 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.74
+ $X2=0.87 $Y2=2.74
r183 54 56 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.87 $Y2=1.59
r184 49 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.81 $Y=1.48
+ $X2=7.81 $Y2=1.48
r185 49 52 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.81 $Y=1.48
+ $X2=7.81 $Y2=1.59
r186 47 56 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.59
+ $X2=0.87 $Y2=1.59
r187 46 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=1.23 $Y2=1.59
r188 46 47 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=0.955 $Y2=1.59
r189 45 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.655
+ $X2=0.87 $Y2=2.74
r190 44 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=1.59
r191 44 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=2.655
r192 40 42 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r193 38 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=2.74
r194 38 40 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=3.455
r195 34 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=1.59
r196 34 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=0.825
r197 32 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.81
+ $Y=1.59 $X2=7.81 $Y2=1.59
r198 30 32 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.685 $Y=1.59
+ $X2=7.81 $Y2=1.59
r199 28 30 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.615 $Y=1.59
+ $X2=7.685 $Y2=1.59
r200 24 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.59 $X2=1.23 $Y2=1.59
r201 24 26 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.23 $Y=1.59
+ $X2=1.425 $Y2=1.59
r202 20 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.685 $Y=1.425
+ $X2=7.685 $Y2=1.59
r203 20 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.685 $Y=1.425
+ $X2=7.685 $Y2=0.945
r204 16 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.755
+ $X2=7.615 $Y2=1.59
r205 16 18 1707.51 $w=1.5e-07 $l=3.33e-06 $layer=POLY_cond $X=7.615 $Y=1.755
+ $X2=7.615 $Y2=5.085
r206 12 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.755
+ $X2=1.425 $Y2=1.59
r207 12 14 1707.51 $w=1.5e-07 $l=3.33e-06 $layer=POLY_cond $X=1.425 $Y=1.755
+ $X2=1.425 $Y2=5.085
r208 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.425
+ $X2=1.425 $Y2=1.59
r209 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.425
+ $X2=1.425 $Y2=0.945
r210 3 42 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r211 3 40 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r212 1 36 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_342_518# 1 3 11 15 18 22 24 25 26 27
+ 28 30 33 37 44 47
c86 47 0 1.71621e-19 $X=3.457 $Y=1.415
c87 25 0 1.29912e-19 $X=3.28 $Y=1.765
r88 46 47 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.457 $Y=1.245
+ $X2=3.457 $Y2=1.415
r89 42 44 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.94 $Y=2.755
+ $X2=2.11 $Y2=2.755
r90 37 39 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=3.465 $Y=3.455
+ $X2=3.465 $Y2=5.835
r91 35 37 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=3.465 $Y=3.27
+ $X2=3.465 $Y2=3.455
r92 33 46 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=3.465 $Y=0.825
+ $X2=3.465 $Y2=1.245
r93 30 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=1.68
+ $X2=3.365 $Y2=1.415
r94 27 35 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.295 $Y=3.185
+ $X2=3.465 $Y2=3.27
r95 27 28 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.295 $Y=3.185
+ $X2=2.195 $Y2=3.185
r96 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=1.765
+ $X2=3.365 $Y2=1.68
r97 25 26 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.28 $Y=1.765
+ $X2=2.195 $Y2=1.765
r98 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=3.1
+ $X2=2.195 $Y2=3.185
r99 23 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=2.92
+ $X2=2.11 $Y2=2.755
r100 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.11 $Y=2.92
+ $X2=2.11 $Y2=3.1
r101 22 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=2.59
+ $X2=2.11 $Y2=2.755
r102 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=1.85
+ $X2=2.195 $Y2=1.765
r103 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.11 $Y=1.85
+ $X2=2.11 $Y2=2.59
r104 18 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.755 $X2=1.94 $Y2=2.755
r105 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.755
+ $X2=1.892 $Y2=2.92
r106 18 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.755
+ $X2=1.892 $Y2=2.59
r107 15 19 843.5 $w=1.5e-07 $l=1.645e-06 $layer=POLY_cond $X=1.855 $Y=0.945
+ $X2=1.855 $Y2=2.59
r108 11 20 1110.14 $w=1.5e-07 $l=2.165e-06 $layer=POLY_cond $X=1.785 $Y=5.085
+ $X2=1.785 $Y2=2.92
r109 3 39 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=3.24
+ $Y=3.085 $X2=3.465 $Y2=5.835
r110 3 37 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=3.24
+ $Y=3.085 $X2=3.465 $Y2=3.455
r111 1 33 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=3.24
+ $Y=0.575 $X2=3.465 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%D 3 7 10 14 19
c41 19 0 1.41836e-19 $X=2.865 $Y=2.22
c42 10 0 1.12321e-19 $X=2.865 $Y=2.22
r43 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.865 $Y=2.22
+ $X2=2.865 $Y2=2.22
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=2.22 $X2=2.865 $Y2=2.22
r45 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=2.22
+ $X2=2.865 $Y2=2.385
r46 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=2.22
+ $X2=2.865 $Y2=2.055
r47 7 12 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=2.805 $Y=4.585
+ $X2=2.805 $Y2=2.385
r48 3 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.805 $Y=1.075
+ $X2=2.805 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c219 55 0 6.79641e-20 $X=5.06 $Y=2.59
c220 48 0 1.98654e-19 $X=3.705 $Y=1.85
c221 44 0 1.86602e-19 $X=3.62 $Y=2.59
c222 30 0 1.29912e-19 $X=3.705 $Y=1.685
c223 25 0 1.41836e-19 $X=3.225 $Y=2.765
r224 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=2.59
+ $X2=5.455 $Y2=2.59
r225 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.305 $Y=2.59
+ $X2=6.45 $Y2=2.59
r226 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.305 $Y=2.59
+ $X2=5.6 $Y2=2.59
r227 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.37 $Y=2.59
+ $X2=3.225 $Y2=2.59
r228 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.31 $Y=2.59
+ $X2=5.455 $Y2=2.59
r229 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.31 $Y=2.59
+ $X2=3.37 $Y2=2.59
r230 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=2.59
+ $X2=5.455 $Y2=2.59
r231 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.455 $Y=2.59
+ $X2=5.455 $Y2=2.765
r232 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.225 $Y=2.59
+ $X2=3.225 $Y2=2.59
r233 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.225 $Y=2.59
+ $X2=3.225 $Y2=2.765
r234 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.45 $Y=2.59
+ $X2=6.45 $Y2=2.59
r235 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.45 $Y=2.59
+ $X2=6.45 $Y2=2.765
r236 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.59
+ $X2=5.455 $Y2=2.59
r237 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.37 $Y=2.59
+ $X2=5.06 $Y2=2.59
r238 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=2.505
+ $X2=5.06 $Y2=2.59
r239 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.975 $Y=2.505
+ $X2=4.975 $Y2=1.85
r240 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.705 $Y=2.505
+ $X2=3.705 $Y2=1.85
r241 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.59
+ $X2=3.225 $Y2=2.59
r242 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.59
+ $X2=3.705 $Y2=2.505
r243 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.62 $Y=2.59
+ $X2=3.31 $Y2=2.59
r244 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=2.765 $X2=6.45 $Y2=2.765
r245 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.332 $Y=1.685
+ $X2=6.332 $Y2=1.835
r246 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=2.765 $X2=5.455 $Y2=2.765
r247 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=2.765
+ $X2=5.455 $Y2=2.93
r248 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.85 $X2=4.975 $Y2=1.85
r249 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.85
+ $X2=4.975 $Y2=1.685
r250 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.85 $X2=3.705 $Y2=1.85
r251 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.85
+ $X2=3.705 $Y2=1.685
r252 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=2.765 $X2=3.225 $Y2=2.765
r253 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.765
+ $X2=3.225 $Y2=2.93
r254 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.36 $Y=2.6
+ $X2=6.407 $Y2=2.765
r255 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.36 $Y=2.6
+ $X2=6.36 $Y2=1.835
r256 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.305 $Y=2.93
+ $X2=6.407 $Y2=2.765
r257 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=6.305 $Y=2.93
+ $X2=6.305 $Y2=4.585
r258 17 40 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.305 $Y=1.075
+ $X2=6.305 $Y2=1.685
r259 13 39 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.515 $Y=4.585
+ $X2=5.515 $Y2=2.93
r260 10 34 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.915 $Y=1.075
+ $X2=4.915 $Y2=1.685
r261 7 30 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.765 $Y=1.075
+ $X2=3.765 $Y2=1.685
r262 3 27 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.165 $Y=4.585
+ $X2=3.165 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_217_817# 1 3 11 15 17 18 21 22 27 31
+ 35 39 40 43 49 54 55 56 61
c140 55 0 1.35571e-19 $X=4.06 $Y=1.85
c141 49 0 1.5821e-19 $X=4.295 $Y=2.765
c142 31 0 6.36774e-20 $X=4.555 $Y=4.585
c143 22 0 1.86602e-19 $X=4.2 $Y=2.765
c144 21 0 6.79641e-20 $X=4.48 $Y=2.765
c145 15 0 6.36774e-20 $X=4.125 $Y=4.585
r146 56 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.785 $Y=1.85
+ $X2=1.64 $Y2=1.85
r147 55 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.85
+ $X2=4.205 $Y2=1.85
r148 55 56 2.19056 $w=1.7e-07 $l=2.275e-06 $layer=MET1_cond $X=4.06 $Y=1.85
+ $X2=1.785 $Y2=1.85
r149 52 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=1.85
+ $X2=4.205 $Y2=1.85
r150 52 54 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=1.81
+ $X2=4.295 $Y2=1.81
r151 47 54 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.295 $Y=1.935
+ $X2=4.295 $Y2=1.81
r152 47 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.295 $Y=1.935
+ $X2=4.295 $Y2=2.765
r153 46 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.85
+ $X2=1.64 $Y2=1.85
r154 43 46 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=1.64 $Y=0.825
+ $X2=1.64 $Y2=1.85
r155 41 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=1.935
+ $X2=1.64 $Y2=1.85
r156 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=2.02
+ $X2=1.64 $Y2=1.935
r157 39 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.555 $Y=2.02
+ $X2=1.295 $Y2=2.02
r158 35 37 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.21 $Y=4.475
+ $X2=1.21 $Y2=5.835
r159 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.295 $Y2=2.02
r160 33 35 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.21 $Y2=4.475
r161 29 31 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.555 $Y2=4.585
r162 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.555 $Y2=1.075
r163 24 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=2.765 $X2=4.295 $Y2=2.765
r164 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=2.765
+ $X2=4.295 $Y2=2.765
r165 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=2.765
+ $X2=4.555 $Y2=2.9
r166 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=2.765
+ $X2=4.295 $Y2=2.765
r167 20 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.85 $X2=4.295 $Y2=1.85
r168 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=1.85
+ $X2=4.295 $Y2=1.85
r169 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=1.85
+ $X2=4.555 $Y2=1.715
r170 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=1.85
+ $X2=4.295 $Y2=1.85
r171 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=2.9
+ $X2=4.2 $Y2=2.765
r172 13 15 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.125 $Y=2.9
+ $X2=4.125 $Y2=4.585
r173 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=1.715
+ $X2=4.2 $Y2=1.85
r174 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.125 $Y=1.715
+ $X2=4.125 $Y2=1.075
r175 3 37 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=4.085 $X2=1.21 $Y2=5.835
r176 3 35 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=4.085 $X2=1.21 $Y2=4.475
r177 1 43 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_618_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c187 35 0 1.98654e-19 $X=3.285 $Y=1.76
c188 18 0 1.12321e-19 $X=3.765 $Y=4.585
r189 66 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=3.185
+ $X2=6.795 $Y2=3.185
r190 62 64 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=2.19
+ $X2=6.795 $Y2=2.19
r191 60 68 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=3.1
+ $X2=6.795 $Y2=3.185
r192 59 64 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.275
+ $X2=6.795 $Y2=2.19
r193 59 60 50.8333 $w=1.78e-07 $l=8.25e-07 $layer=LI1_cond $X=6.795 $Y=2.275
+ $X2=6.795 $Y2=3.1
r194 55 57 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.52 $Y=3.455
+ $X2=6.52 $Y2=5.835
r195 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=3.27
+ $X2=6.52 $Y2=3.185
r196 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.52 $Y=3.27
+ $X2=6.52 $Y2=3.455
r197 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.105
+ $X2=6.52 $Y2=2.19
r198 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.935
+ $X2=6.52 $Y2=1.85
r199 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=1.935
+ $X2=6.52 $Y2=2.105
r200 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.765
+ $X2=6.52 $Y2=1.85
r201 47 49 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.52 $Y=1.765
+ $X2=6.52 $Y2=0.825
r202 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=1.85
+ $X2=6.52 $Y2=1.85
r203 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.435 $Y=1.85
+ $X2=5.455 $Y2=1.85
r204 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.85 $X2=5.455 $Y2=1.85
r205 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.85
+ $X2=5.455 $Y2=2.015
r206 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.85
+ $X2=5.455 $Y2=1.685
r207 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.165 $Y=1.76
+ $X2=3.285 $Y2=1.76
r208 32 41 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.515 $Y=1.075
+ $X2=5.515 $Y2=1.685
r209 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.395 $Y=2.225
+ $X2=5.395 $Y2=2.015
r210 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.99 $Y=2.3
+ $X2=4.915 $Y2=2.3
r211 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.32 $Y=2.3
+ $X2=5.395 $Y2=2.225
r212 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.32 $Y=2.3
+ $X2=4.99 $Y2=2.3
r213 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.915 $Y=2.375
+ $X2=4.915 $Y2=2.3
r214 22 24 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=4.915 $Y=2.375
+ $X2=4.915 $Y2=4.585
r215 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.3
+ $X2=3.765 $Y2=2.3
r216 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=2.3
+ $X2=4.915 $Y2=2.3
r217 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.84 $Y=2.3 $X2=3.84
+ $Y2=2.3
r218 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=2.375
+ $X2=3.765 $Y2=2.3
r219 16 18 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=3.765 $Y=2.375
+ $X2=3.765 $Y2=4.585
r220 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=2.3
+ $X2=3.765 $Y2=2.3
r221 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.69 $Y=2.3
+ $X2=3.36 $Y2=2.3
r222 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.285 $Y=2.225
+ $X2=3.36 $Y2=2.3
r223 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.835
+ $X2=3.285 $Y2=1.76
r224 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.285 $Y=1.835
+ $X2=3.285 $Y2=2.225
r225 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.685
+ $X2=3.165 $Y2=1.76
r226 9 11 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.165 $Y=1.685
+ $X2=3.165 $Y2=1.075
r227 3 57 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=5.835
r228 3 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=3.455
r229 1 49 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_1160_89# 1 3 11 15 23 26 28 32 33 35
+ 36 37 38 40 46 50 51 54 57 60 63 64 65 70
c160 37 0 8.77106e-20 $X=8.61 $Y=2.855
c161 32 0 2.20654e-19 $X=8.52 $Y=2.19
r162 65 67 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=2.19
+ $X2=5.935 $Y2=2.19
r163 64 70 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.375 $Y=2.19
+ $X2=8.52 $Y2=2.19
r164 64 65 2.20982 $w=1.7e-07 $l=2.295e-06 $layer=MET1_cond $X=8.375 $Y=2.19
+ $X2=6.08 $Y2=2.19
r165 60 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.52 $Y=2.19
+ $X2=8.52 $Y2=2.19
r166 58 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=2.19
+ $X2=7.47 $Y2=2.19
r167 58 60 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.555 $Y=2.19
+ $X2=8.52 $Y2=2.19
r168 56 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=2.275
+ $X2=7.47 $Y2=2.19
r169 56 57 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.47 $Y=2.275
+ $X2=7.47 $Y2=3.695
r170 52 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=2.105
+ $X2=7.47 $Y2=2.19
r171 52 54 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=7.47 $Y=2.105
+ $X2=7.47 $Y2=0.825
r172 50 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=3.78
+ $X2=7.47 $Y2=3.695
r173 50 51 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.385 $Y=3.78
+ $X2=7.125 $Y2=3.78
r174 46 48 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.04 $Y=4.475
+ $X2=7.04 $Y2=5.835
r175 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=3.865
+ $X2=7.125 $Y2=3.78
r176 44 46 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.04 $Y=3.865
+ $X2=7.04 $Y2=4.475
r177 40 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.935 $Y=2.19
+ $X2=5.935 $Y2=2.19
r178 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=2.855
+ $X2=8.61 $Y2=3.005
r179 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=1.65 $X2=8.61
+ $Y2=1.8
r180 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=8.585 $Y=2.355
+ $X2=8.585 $Y2=2.855
r181 33 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.585 $Y=2.025
+ $X2=8.585 $Y2=1.8
r182 32 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.52
+ $Y=2.19 $X2=8.52 $Y2=2.19
r183 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=2.19
+ $X2=8.522 $Y2=2.355
r184 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=2.19
+ $X2=8.522 $Y2=2.025
r185 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.935
+ $Y=2.19 $X2=5.935 $Y2=2.19
r186 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=2.19
+ $X2=5.935 $Y2=2.355
r187 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=2.19
+ $X2=5.935 $Y2=2.025
r188 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=8.635 $Y=4.585
+ $X2=8.635 $Y2=3.005
r189 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.635 $Y=1.075
+ $X2=8.635 $Y2=1.65
r190 15 30 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=5.875 $Y=4.585
+ $X2=5.875 $Y2=2.355
r191 11 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.875 $Y=1.075
+ $X2=5.875 $Y2=2.025
r192 3 48 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=4.085 $X2=7.04 $Y2=5.835
r193 3 46 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=4.085 $X2=7.04 $Y2=4.475
r194 1 54 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.575 $X2=7.47 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_998_115# 1 3 11 13 15 22 23 24 25 26
+ 29 33 38 42 43 48
c131 43 0 1.5821e-19 $X=4.78 $Y=1.85
c132 23 0 1.67294e-19 $X=5.045 $Y=1.43
c133 22 0 1.57671e-19 $X=4.635 $Y=1.85
r134 43 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.78 $Y=1.85
+ $X2=4.635 $Y2=1.85
r135 42 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=1.85
+ $X2=7.13 $Y2=1.85
r136 42 43 2.12316 $w=1.7e-07 $l=2.205e-06 $layer=MET1_cond $X=6.985 $Y=1.85
+ $X2=4.78 $Y2=1.85
r137 38 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=1.85
+ $X2=7.13 $Y2=1.85
r138 33 35 69.1466 $w=3.38e-07 $l=2.04e-06 $layer=LI1_cond $X=5.215 $Y=3.795
+ $X2=5.215 $Y2=5.835
r139 31 33 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=5.215 $Y=3.27
+ $X2=5.215 $Y2=3.795
r140 27 29 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=5.215 $Y=1.345
+ $X2=5.215 $Y2=0.825
r141 25 31 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=3.185
+ $X2=5.215 $Y2=3.27
r142 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=3.185
+ $X2=4.72 $Y2=3.185
r143 23 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=1.43
+ $X2=5.215 $Y2=1.345
r144 23 24 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=1.43
+ $X2=4.72 $Y2=1.43
r145 22 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.85
+ $X2=4.635 $Y2=1.85
r146 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=3.1
+ $X2=4.72 $Y2=3.185
r147 20 22 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.635 $Y=3.1
+ $X2=4.635 $Y2=1.85
r148 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=1.515
+ $X2=4.72 $Y2=1.43
r149 19 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.635 $Y=1.515
+ $X2=4.635 $Y2=1.85
r150 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.85 $X2=7.13 $Y2=1.85
r151 13 18 38.6212 $w=3.33e-07 $l=2.06325e-07 $layer=POLY_cond $X=7.255 $Y=2.015
+ $X2=7.162 $Y2=1.85
r152 13 15 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=7.255 $Y=2.015
+ $X2=7.255 $Y2=5.085
r153 9 18 39.3449 $w=3.33e-07 $l=2.11447e-07 $layer=POLY_cond $X=7.255 $Y=1.68
+ $X2=7.162 $Y2=1.85
r154 9 11 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=7.255 $Y=1.68
+ $X2=7.255 $Y2=0.945
r155 3 35 171.429 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=3 $X=4.99
+ $Y=3.085 $X2=5.215 $Y2=5.835
r156 3 33 171.429 $w=1.7e-07 $l=8.1477e-07 $layer=licon1_PDIFF $count=3 $X=4.99
+ $Y=3.085 $X2=5.215 $Y2=3.795
r157 1 29 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=4.99
+ $Y=0.575 $X2=5.215 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c80 44 0 8.77106e-20 $X=8.425 $Y=2.96
c81 35 0 9.99996e-20 $X=8.92 $Y=2.765
c82 33 0 1.20654e-19 $X=8.92 $Y=1.85
c83 23 0 1.88625e-19 $X=8.42 $Y=0.825
r84 42 44 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=8.42 $Y=2.96
+ $X2=8.425 $Y2=2.96
r85 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.005 $Y=2.68
+ $X2=9.005 $Y2=2.395
r86 37 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.005 $Y=1.935
+ $X2=9.005 $Y2=2.395
r87 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=2.765
+ $X2=9.005 $Y2=2.68
r88 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=2.765
+ $X2=8.505 $Y2=2.765
r89 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=1.85
+ $X2=9.005 $Y2=1.935
r90 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=1.85
+ $X2=8.505 $Y2=1.85
r91 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=8.42 $Y=4.475
+ $X2=8.42 $Y2=5.835
r92 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.42 $Y=2.96
+ $X2=8.42 $Y2=2.96
r93 27 29 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=8.42 $Y=2.96
+ $X2=8.42 $Y2=4.475
r94 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=2.85
+ $X2=8.505 $Y2=2.765
r95 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.42 $Y=2.85
+ $X2=8.42 $Y2=2.96
r96 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=1.765
+ $X2=8.505 $Y2=1.85
r97 21 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=8.42 $Y=1.765
+ $X2=8.42 $Y2=0.825
r98 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=2.395 $X2=9.005 $Y2=2.395
r99 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=2.395
+ $X2=9.005 $Y2=2.56
r100 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=2.395
+ $X2=9.005 $Y2=2.23
r101 15 20 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=9.065 $Y=4.585
+ $X2=9.065 $Y2=2.56
r102 11 19 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.065 $Y=1.075
+ $X2=9.065 $Y2=2.23
r103 3 31 240 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=3.085 $X2=8.42 $Y2=5.835
r104 3 29 240 $w=1.7e-07 $l=1.45115e-06 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=3.085 $X2=8.42 $Y2=4.475
r105 1 23 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.575 $X2=8.42 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%Q 1 3 11 15 20 23 27 30
r21 27 28 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=3.287
+ $X2=9.395 $Y2=3.287
r22 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=3.33
+ $X2=9.275 $Y2=3.33
r23 26 27 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=9.275 $Y=3.287
+ $X2=9.28 $Y2=3.287
r24 21 23 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=1.515
+ $X2=9.395 $Y2=1.515
r25 20 28 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.395 $Y=3.16
+ $X2=9.395 $Y2=3.287
r26 19 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.6
+ $X2=9.395 $Y2=1.515
r27 19 20 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=9.395 $Y=1.6
+ $X2=9.395 $Y2=3.16
r28 15 17 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=9.28 $Y=4.475
+ $X2=9.28 $Y2=5.835
r29 13 27 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.28 $Y=3.415
+ $X2=9.28 $Y2=3.287
r30 13 15 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=9.28 $Y=3.415
+ $X2=9.28 $Y2=4.475
r31 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=1.43 $X2=9.28
+ $Y2=1.515
r32 9 11 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.28 $Y=1.43
+ $X2=9.28 $Y2=0.825
r33 3 17 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=3.085 $X2=9.28 $Y2=5.835
r34 3 15 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=3.085 $X2=9.28 $Y2=4.475
r35 1 11 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.575 $X2=9.28 $Y2=0.825
.ends

