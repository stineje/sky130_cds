* File: sky130_osu_sc_15T_ms__inv_6.spice
* Created: Fri Nov 12 14:44:28 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__inv_6.pex.spice"
.subckt sky130_osu_sc_15T_ms__inv_6  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1003 N_GND_M1003_d N_A_M1003_g N_Y_M1001_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1007 N_GND_M1003_d N_A_M1007_g N_Y_M1007_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_GND_M1009_d N_A_M1009_g N_Y_M1007_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_GND_M1009_d N_A_M1010_g N_Y_M1010_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_GND_M1011_d N_A_M1011_g N_Y_M1010_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75002.3 A=0.3 P=4.3 MULT=1
MM1002 N_VDD_M1002_d N_A_M1002_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75001.9 A=0.3 P=4.3 MULT=1
MM1004 N_VDD_M1002_d N_A_M1004_g N_Y_M1004_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001 SB=75001.5
+ A=0.3 P=4.3 MULT=1
MM1005 N_VDD_M1005_d N_A_M1005_g N_Y_M1004_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001.5 SB=75001
+ A=0.3 P=4.3 MULT=1
MM1006 N_VDD_M1005_d N_A_M1006_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001.9
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1008 N_VDD_M1008_d N_A_M1008_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75002.3
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX12_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=9.558 P=12.38
pX13_noxref noxref_5 A A PROBETYPE=1
pX14_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__inv_6.pxi.spice"
*
.ends
*
*
