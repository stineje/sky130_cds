* File: sky130_osu_sc_18T_hs__ncgate_1.pex.spice
* Created: Thu Mar 10 17:10:01 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%GND 1 2 3 4 5 6 7 89 93 95 102 104 111
+ 113 123 125 135 137 141 143 151 168 170 175 177 179 181 183 185 187 189 191
+ 193
c181 135 0 1.97615e-19 $X=3.99 $Y=0.8
r182 191 193 0.00232861 $w=3.05e-07 $l=5e-09 $layer=MET1_cond $X=5.695 $Y=0.127
+ $X2=5.7 $Y2=0.127
r183 189 191 0.312033 $w=3.05e-07 $l=6.7e-07 $layer=MET1_cond $X=5.025 $Y=0.127
+ $X2=5.695 $Y2=0.127
r184 187 189 0.454078 $w=3.05e-07 $l=9.75e-07 $layer=MET1_cond $X=4.05 $Y=0.127
+ $X2=5.025 $Y2=0.127
r185 185 187 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=3.365 $Y=0.127
+ $X2=4.05 $Y2=0.127
r186 183 185 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=2.68 $Y=0.127
+ $X2=3.365 $Y2=0.127
r187 181 183 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=2 $Y=0.127
+ $X2=2.68 $Y2=0.127
r188 179 181 0.314362 $w=3.05e-07 $l=6.75e-07 $layer=MET1_cond $X=1.325 $Y=0.127
+ $X2=2 $Y2=0.127
r189 177 179 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.645 $Y=0.127
+ $X2=1.325 $Y2=0.127
r190 175 177 0.430792 $w=3.05e-07 $l=9.25e-07 $layer=MET1_cond $X=-0.28 $Y=0.127
+ $X2=0.645 $Y2=0.127
r191 173 175 0.316225 $w=3.05e-07 $l=6.79e-07 $layer=MET1_cond $X=-0.959
+ $Y=0.127 $X2=-0.28 $Y2=0.127
r192 170 173 0.000465721 $w=3.05e-07 $l=1e-09 $layer=MET1_cond $X=-0.96 $Y=0.127
+ $X2=-0.959 $Y2=0.127
r193 149 168 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.8 $Y=0.28
+ $X2=5.8 $Y2=0.127
r194 149 151 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.8 $Y=0.28
+ $X2=5.8 $Y2=0.8
r195 143 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=0.127
+ $X2=5.8 $Y2=0.127
r196 139 141 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.94 $Y=0.28
+ $X2=4.94 $Y2=0.8
r197 137 138 29.4723 $w=3.03e-07 $l=7.8e-07 $layer=LI1_cond $X=4.855 $Y=0.127
+ $X2=4.075 $Y2=0.127
r198 133 135 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.99 $Y=0.28
+ $X2=3.99 $Y2=0.8
r199 126 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.127
+ $X2=2.52 $Y2=0.127
r200 121 161 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.52 $Y=0.28
+ $X2=2.52 $Y2=0.127
r201 121 123 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.52 $Y=0.28
+ $X2=2.52 $Y2=0.8
r202 114 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.127
+ $X2=0.77 $Y2=0.127
r203 113 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.127
+ $X2=2.52 $Y2=0.127
r204 109 160 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.77 $Y=0.28
+ $X2=0.77 $Y2=0.127
r205 109 111 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.77 $Y=0.28
+ $X2=0.77 $Y2=0.8
r206 105 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.095 $Y=0.127
+ $X2=-0.18 $Y2=0.127
r207 104 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.127
+ $X2=0.77 $Y2=0.127
r208 100 159 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=-0.18 $Y=0.28
+ $X2=-0.18 $Y2=0.127
r209 100 102 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=-0.18 $Y=0.28
+ $X2=-0.18 $Y2=0.8
r210 95 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.265 $Y=0.127
+ $X2=-0.18 $Y2=0.127
r211 91 93 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=-1.04 $Y=0.28
+ $X2=-1.04 $Y2=0.8
r212 89 193 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.7 $Y=0.165
+ $X2=5.7 $Y2=0.165
r213 89 173 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=-0.959 $Y=0.165
+ $X2=-0.959 $Y2=0.165
r214 89 139 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.94 $Y=0.127
+ $X2=4.94 $Y2=0.28
r215 89 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=0.127
+ $X2=4.855 $Y2=0.127
r216 89 144 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=0.127
+ $X2=5.025 $Y2=0.127
r217 89 133 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.99 $Y=0.127
+ $X2=3.99 $Y2=0.28
r218 89 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=0.127
+ $X2=3.905 $Y2=0.127
r219 89 138 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=0.127
+ $X2=4.075 $Y2=0.127
r220 89 91 4.35274 $w=1.7e-07 $l=1.98681e-07 $layer=LI1_cond $X=-1.145 $Y=0.127
+ $X2=-1.04 $Y2=0.28
r221 89 96 3.2055 $w=3.05e-07 $l=1.9e-07 $layer=LI1_cond $X=-1.145 $Y=0.127
+ $X2=-0.955 $Y2=0.127
r222 89 143 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=5.7 $Y=0.127
+ $X2=5.715 $Y2=0.127
r223 89 144 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=5.7 $Y=0.127
+ $X2=5.025 $Y2=0.127
r224 89 125 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.365 $Y=0.127
+ $X2=3.905 $Y2=0.127
r225 89 126 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=2.685 $Y=0.127
+ $X2=2.605 $Y2=0.127
r226 89 113 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.005 $Y=0.127
+ $X2=2.435 $Y2=0.127
r227 89 114 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.325 $Y=0.127
+ $X2=0.855 $Y2=0.127
r228 89 104 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=0.645 $Y=0.127
+ $X2=0.685 $Y2=0.127
r229 89 105 27.9609 $w=3.03e-07 $l=7.4e-07 $layer=LI1_cond $X=0.645 $Y=0.127
+ $X2=-0.095 $Y2=0.127
r230 89 95 0.52899 $w=3.03e-07 $l=1.4e-08 $layer=LI1_cond $X=-0.279 $Y=0.127
+ $X2=-0.265 $Y2=0.127
r231 89 96 25.5427 $w=3.03e-07 $l=6.76e-07 $layer=LI1_cond $X=-0.279 $Y=0.127
+ $X2=-0.955 $Y2=0.127
r232 7 151 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.66
+ $Y=0.55 $X2=5.8 $Y2=0.8
r233 6 141 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=4.815
+ $Y=0.55 $X2=4.94 $Y2=0.8
r234 5 135 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.85
+ $Y=0.55 $X2=3.99 $Y2=0.8
r235 4 123 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.38
+ $Y=0.55 $X2=2.52 $Y2=0.8
r236 3 111 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.55 $X2=0.77 $Y2=0.8
r237 2 102 91 $w=1.7e-07 $l=3.1265e-07 $layer=licon1_NDIFF $count=2 $X=-0.32
+ $Y=0.55 $X2=-0.179 $Y2=0.8
r238 1 93 91 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=2 $X=-1.165
+ $Y=0.55 $X2=-1.039 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%VDD 1 2 3 4 5 61 63 70 74 80 84 92 96
+ 104 108 117 129 134 136 138 140
r108 138 140 1.40182 $w=3.05e-07 $l=3.01e-06 $layer=MET1_cond $X=2.69 $Y=6.482
+ $X2=5.7 $Y2=6.482
r109 136 138 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=2.005 $Y=6.482
+ $X2=2.69 $Y2=6.482
r110 134 136 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=1.32 $Y=6.482
+ $X2=2.005 $Y2=6.482
r111 131 134 1.06138 $w=3.05e-07 $l=2.279e-06 $layer=MET1_cond $X=-0.959
+ $Y=6.482 $X2=1.32 $Y2=6.482
r112 117 120 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=5.8 $Y=4.11
+ $X2=5.8 $Y2=5.81
r113 115 129 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.8 $Y=6.33
+ $X2=5.8 $Y2=6.482
r114 115 120 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.8 $Y=6.33
+ $X2=5.8 $Y2=5.81
r115 113 140 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.7 $Y=6.445
+ $X2=5.7 $Y2=6.445
r116 111 113 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.02 $Y=6.482
+ $X2=5.7 $Y2=6.482
r117 109 128 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=6.482
+ $X2=3.99 $Y2=6.482
r118 109 111 35.7068 $w=3.03e-07 $l=9.45e-07 $layer=LI1_cond $X=4.075 $Y=6.482
+ $X2=5.02 $Y2=6.482
r119 108 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=6.482
+ $X2=5.8 $Y2=6.482
r120 108 113 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=5.715 $Y=6.482
+ $X2=5.7 $Y2=6.482
r121 104 107 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.99 $Y=3.43
+ $X2=3.99 $Y2=5.81
r122 102 128 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.99 $Y=6.33
+ $X2=3.99 $Y2=6.482
r123 102 107 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.99 $Y=6.33
+ $X2=3.99 $Y2=5.81
r124 99 101 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.685 $Y=6.482
+ $X2=3.365 $Y2=6.482
r125 97 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=6.482
+ $X2=2.52 $Y2=6.482
r126 97 99 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=2.605 $Y=6.482
+ $X2=2.685 $Y2=6.482
r127 96 128 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=6.482
+ $X2=3.99 $Y2=6.482
r128 96 101 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.905 $Y=6.482
+ $X2=3.365 $Y2=6.482
r129 92 95 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.52 $Y=3.43
+ $X2=2.52 $Y2=5.81
r130 90 126 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.52 $Y=6.33
+ $X2=2.52 $Y2=6.482
r131 90 95 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.52 $Y=6.33
+ $X2=2.52 $Y2=5.81
r132 87 89 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.325 $Y=6.482
+ $X2=2.005 $Y2=6.482
r133 85 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=6.482
+ $X2=0.77 $Y2=6.482
r134 85 87 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=0.855 $Y=6.482
+ $X2=1.325 $Y2=6.482
r135 84 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=6.482
+ $X2=2.52 $Y2=6.482
r136 84 89 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.435 $Y=6.482
+ $X2=2.005 $Y2=6.482
r137 80 83 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.77 $Y=3.77
+ $X2=0.77 $Y2=5.81
r138 78 125 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.77 $Y=6.33
+ $X2=0.77 $Y2=6.482
r139 78 83 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.77 $Y=6.33
+ $X2=0.77 $Y2=5.81
r140 75 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.165 $Y=6.482
+ $X2=-0.25 $Y2=6.482
r141 75 77 30.6059 $w=3.03e-07 $l=8.1e-07 $layer=LI1_cond $X=-0.165 $Y=6.482
+ $X2=0.645 $Y2=6.482
r142 74 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=6.482
+ $X2=0.77 $Y2=6.482
r143 74 77 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=0.685 $Y=6.482
+ $X2=0.645 $Y2=6.482
r144 70 73 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=-0.25 $Y=4.11
+ $X2=-0.25 $Y2=5.81
r145 68 124 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=-0.25 $Y=6.33
+ $X2=-0.25 $Y2=6.482
r146 68 73 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=-0.25 $Y=6.33
+ $X2=-0.25 $Y2=5.81
r147 65 131 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=-0.959 $Y=6.445
+ $X2=-0.959 $Y2=6.445
r148 63 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.335 $Y=6.482
+ $X2=-0.25 $Y2=6.482
r149 63 65 23.5779 $w=3.03e-07 $l=6.24e-07 $layer=LI1_cond $X=-0.335 $Y=6.482
+ $X2=-0.959 $Y2=6.482
r150 61 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.495 $Y=6.33 $X2=5.7 $Y2=6.415
r151 61 111 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.815 $Y=6.33 $X2=5.02 $Y2=6.415
r152 61 128 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.84 $Y=6.33 $X2=4.045 $Y2=6.415
r153 61 101 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.16 $Y=6.33 $X2=3.365 $Y2=6.415
r154 61 99 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.48 $Y=6.33 $X2=2.685 $Y2=6.415
r155 61 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.8 $Y=6.33 $X2=2.005 $Y2=6.415
r156 61 87 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.12 $Y=6.33 $X2=1.325 $Y2=6.415
r157 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.44 $Y=6.33 $X2=0.645 $Y2=6.415
r158 61 124 182 $w=1.7e-07 $l=2.44839e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=-0.485 $Y=6.33 $X2=-0.279 $Y2=6.415
r159 61 65 182 $w=1.7e-07 $l=2.44839e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=-1.165 $Y=6.33 $X2=-0.959 $Y2=6.415
r160 5 120 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=5.66
+ $Y=3.06 $X2=5.8 $Y2=5.81
r161 5 117 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=5.66
+ $Y=3.06 $X2=5.8 $Y2=4.11
r162 4 107 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.85
+ $Y=3.06 $X2=3.99 $Y2=5.81
r163 4 104 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.85
+ $Y=3.06 $X2=3.99 $Y2=3.43
r164 3 95 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.38
+ $Y=3.06 $X2=2.52 $Y2=5.81
r165 3 92 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.38
+ $Y=3.06 $X2=2.52 $Y2=3.43
r166 2 83 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.63
+ $Y=3.06 $X2=0.77 $Y2=5.81
r167 2 80 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.63
+ $Y=3.06 $X2=0.77 $Y2=3.77
r168 1 73 200 $w=1.7e-07 $l=2.81962e-06 $layer=licon1_PDIFF $count=3 $X=-0.39
+ $Y=3.06 $X2=-0.249 $Y2=5.81
r169 1 70 200 $w=1.7e-07 $l=1.11828e-06 $layer=licon1_PDIFF $count=3 $X=-0.39
+ $Y=3.06 $X2=-0.249 $Y2=4.11
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%SE 3 7 10 13 19 22 25
r50 22 25 0.000586854 $w=2.13e-07 $l=1e-09 $layer=MET1_cond $X=-0.65 $Y=2.935
+ $X2=-0.649 $Y2=2.935
r51 19 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-0.649 $Y=2.935
+ $X2=-0.649 $Y2=2.935
r52 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=-0.65 $Y=2.15
+ $X2=-0.65 $Y2=2.935
r53 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=-0.735 $Y=2.065
+ $X2=-0.65 $Y2=2.15
r54 13 15 9.72086 $w=1.68e-07 $l=1.49e-07 $layer=LI1_cond $X=-0.735 $Y=2.065
+ $X2=-0.884 $Y2=2.065
r55 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=-0.884
+ $Y=2.065 $X2=-0.884 $Y2=2.065
r56 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.885 $Y=2.065
+ $X2=-0.885 $Y2=2.23
r57 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.885 $Y=2.065
+ $X2=-0.885 $Y2=1.9
r58 7 12 1194.74 $w=1.5e-07 $l=2.33e-06 $layer=POLY_cond $X=-0.825 $Y=4.56
+ $X2=-0.825 $Y2=2.23
r59 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=-0.825 $Y=1.05
+ $X2=-0.825 $Y2=1.9
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%E 3 7 10 14 22 24
r47 22 24 0.000584112 $w=2.14e-07 $l=1e-09 $layer=MET1_cond $X=-0.305 $Y=3.305
+ $X2=-0.304 $Y2=3.305
r48 20 22 0.00233645 $w=2.14e-07 $l=4e-09 $layer=MET1_cond $X=-0.309 $Y=3.305
+ $X2=-0.305 $Y2=3.305
r49 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-0.309 $Y=3.305
+ $X2=-0.309 $Y2=3.305
r50 14 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=-0.31 $Y=2.73
+ $X2=-0.31 $Y2=3.305
r51 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=-0.309
+ $Y=2.73 $X2=-0.309 $Y2=2.73
r52 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.357 $Y=2.73
+ $X2=-0.357 $Y2=2.895
r53 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.357 $Y=2.73
+ $X2=-0.357 $Y2=2.565
r54 7 11 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=-0.395 $Y=1.05
+ $X2=-0.395 $Y2=2.565
r55 3 12 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=-0.465 $Y=4.56
+ $X2=-0.465 $Y2=2.895
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_86_332# 1 3 13 16 18 19 21 22 23 24
+ 25 27 28 30 31 32 35 39
r83 39 41 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.645 $Y=3.43
+ $X2=1.645 $Y2=5.81
r84 37 39 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=3.43
r85 33 35 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=1.645 $Y=1.32
+ $X2=1.645 $Y2=0.8
r86 31 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.475 $Y=1.405
+ $X2=1.645 $Y2=1.32
r87 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.475 $Y=1.405
+ $X2=1.195 $Y2=1.405
r88 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.11 $Y=1.49
+ $X2=1.195 $Y2=1.405
r89 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.11 $Y=1.49
+ $X2=1.11 $Y2=1.74
r90 27 37 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.475 $Y=3.16
+ $X2=1.645 $Y2=3.245
r91 27 28 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.475 $Y=3.16
+ $X2=0.65 $Y2=3.16
r92 26 44 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.65 $Y=1.825
+ $X2=0.565 $Y2=1.785
r93 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.025 $Y=1.825
+ $X2=1.11 $Y2=1.74
r94 25 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.025 $Y=1.825
+ $X2=0.65 $Y2=1.825
r95 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=3.075
+ $X2=0.65 $Y2=3.16
r96 23 44 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=1.91
+ $X2=0.565 $Y2=1.785
r97 23 24 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=0.565 $Y=1.91
+ $X2=0.565 $Y2=3.075
r98 21 22 56.3681 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=0.53 $Y=2.78 $X2=0.53
+ $Y2=2.95
r99 20 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.505 $Y=1.99
+ $X2=0.505 $Y2=2.78
r100 18 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.825 $X2=0.565 $Y2=1.825
r101 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.825
+ $X2=0.565 $Y2=1.99
r102 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.825
+ $X2=0.565 $Y2=1.66
r103 16 22 517.347 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=0.555 $Y=4.56
+ $X2=0.555 $Y2=2.95
r104 13 19 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.555 $Y=1.05
+ $X2=0.555 $Y2=1.66
r105 3 41 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.42
+ $Y=3.06 $X2=1.645 $Y2=5.81
r106 3 39 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.42
+ $Y=3.06 $X2=1.645 $Y2=3.43
r107 1 35 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.55 $X2=1.645 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_N233_612# 1 3 11 15 18 22 30 36 41
+ 42 44 45 51 53
c104 15 0 1.64001e-19 $X=0.985 $Y=4.56
c105 11 0 1.38221e-19 $X=0.985 $Y=1.05
r106 46 53 0.0529306 $w=1.7e-07 $l=8.5e-08 $layer=MET1_cond $X=-0.525 $Y=2.565
+ $X2=-0.61 $Y2=2.565
r107 45 55 0.0903352 $w=2.14e-07 $l=1.47479e-07 $layer=MET1_cond $X=0.78
+ $Y=2.565 $X2=0.925 $Y2=2.57
r108 45 46 1.25656 $w=1.7e-07 $l=1.305e-06 $layer=MET1_cond $X=0.78 $Y=2.565
+ $X2=-0.525 $Y2=2.565
r109 44 53 0.0137558 $w=1.7e-07 $l=8.5e-08 $layer=MET1_cond $X=-0.61 $Y=2.48
+ $X2=-0.61 $Y2=2.565
r110 43 51 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=-0.61 $Y=1.57
+ $X2=-0.61 $Y2=1.455
r111 43 44 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=-0.61 $Y=1.57
+ $X2=-0.61 $Y2=2.48
r112 42 48 0.102734 $w=2.3e-07 $l=1.44e-07 $layer=MET1_cond $X=-0.895 $Y=2.565
+ $X2=-1.039 $Y2=2.565
r113 41 53 0.0529306 $w=1.7e-07 $l=8.5e-08 $layer=MET1_cond $X=-0.695 $Y=2.565
+ $X2=-0.61 $Y2=2.565
r114 41 42 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=-0.695 $Y=2.565
+ $X2=-0.895 $Y2=2.565
r115 39 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.925 $Y=2.57
+ $X2=0.925 $Y2=2.57
r116 36 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.925 $Y=2.4
+ $X2=0.925 $Y2=2.57
r117 33 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-0.609 $Y=1.455
+ $X2=-0.609 $Y2=1.455
r118 30 33 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=-0.61 $Y=0.8
+ $X2=-0.61 $Y2=1.455
r119 25 27 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=-1.04 $Y=3.43
+ $X2=-1.04 $Y2=5.81
r120 22 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-1.039 $Y=2.565
+ $X2=-1.039 $Y2=2.565
r121 22 25 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=-1.04 $Y=2.565
+ $X2=-1.04 $Y2=3.43
r122 18 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.4 $X2=0.925 $Y2=2.4
r123 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.4
+ $X2=0.925 $Y2=2.565
r124 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.4
+ $X2=0.925 $Y2=2.235
r125 15 20 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=0.985 $Y=4.56
+ $X2=0.985 $Y2=2.565
r126 11 19 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.985 $Y=1.05
+ $X2=0.985 $Y2=2.235
r127 3 27 150 $w=1.7e-07 $l=2.81229e-06 $layer=licon1_PDIFF $count=4 $X=-1.165
+ $Y=3.06 $X2=-1.039 $Y2=5.81
r128 3 25 150 $w=1.7e-07 $l=4.28392e-07 $layer=licon1_PDIFF $count=4 $X=-1.165
+ $Y=3.06 $X2=-1.039 $Y2=3.43
r129 1 30 91 $w=1.7e-07 $l=3.1265e-07 $layer=licon1_NDIFF $count=2 $X=-0.75
+ $Y=0.55 $X2=-0.609 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_254_515# 1 3 11 15 17 21 22 25 26 27
+ 32 35 38 43 47 49 52 56
c126 52 0 1.86741e-19 $X=3.22 $Y=2.195
c127 47 0 9.95038e-20 $X=1.485 $Y=2.74
c128 27 0 1.38221e-19 $X=1.57 $Y=1.825
c129 25 0 1.64001e-19 $X=1.485 $Y=2.655
c130 17 0 1.47633e-20 $X=1.405 $Y=2.74
r131 54 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.95 $Y=3.16
+ $X2=3.22 $Y2=3.16
r132 50 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.95 $Y=2.195
+ $X2=3.22 $Y2=2.195
r133 45 47 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.405 $Y=2.74
+ $X2=1.485 $Y2=2.74
r134 43 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=3.075
+ $X2=3.22 $Y2=3.16
r135 42 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.28
+ $X2=3.22 $Y2=2.195
r136 42 43 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.22 $Y=2.28
+ $X2=3.22 $Y2=3.075
r137 38 40 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.95 $Y=3.43
+ $X2=2.95 $Y2=5.81
r138 36 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=3.245
+ $X2=2.95 $Y2=3.16
r139 36 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.95 $Y=3.245
+ $X2=2.95 $Y2=3.43
r140 35 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=2.11
+ $X2=2.95 $Y2=2.195
r141 34 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=1.91
+ $X2=2.95 $Y2=1.825
r142 34 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.95 $Y=1.91 $X2=2.95
+ $Y2=2.11
r143 30 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=1.74
+ $X2=2.95 $Y2=1.825
r144 30 32 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.95 $Y=1.74
+ $X2=2.95 $Y2=0.8
r145 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.57 $Y=1.825
+ $X2=1.885 $Y2=1.825
r146 26 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.825
+ $X2=2.95 $Y2=1.825
r147 26 29 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.865 $Y=1.825
+ $X2=1.885 $Y2=1.825
r148 25 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=2.655
+ $X2=1.485 $Y2=2.74
r149 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=1.91
+ $X2=1.57 $Y2=1.825
r150 24 25 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.485 $Y=1.91
+ $X2=1.485 $Y2=2.655
r151 21 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=1.825 $X2=1.885 $Y2=1.825
r152 21 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.825
+ $X2=1.885 $Y2=1.66
r153 17 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=2.74 $X2=1.405 $Y2=2.74
r154 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=2.74
+ $X2=1.405 $Y2=2.905
r155 15 22 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.945 $Y=1.05
+ $X2=1.945 $Y2=1.66
r156 11 19 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.345 $Y=4.56
+ $X2=1.345 $Y2=2.905
r157 3 40 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.81
+ $Y=3.06 $X2=2.95 $Y2=5.81
r158 3 38 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.81
+ $Y=3.06 $X2=2.95 $Y2=3.43
r159 1 32 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.81
+ $Y=0.55 $X2=2.95 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%CK 3 5 6 11 15 16 18 21 24 28 31 32 34
+ 35 39 43 49 55 58 62 63 64 65 70 74
c192 63 0 1.47633e-20 $X=2.03 $Y=2.565
c193 39 0 8.03558e-20 $X=5.63 $Y=2.36
c194 31 0 1.2087e-19 $X=1.885 $Y=2.74
c195 5 0 9.95038e-20 $X=1.75 $Y=2.275
r196 65 70 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.025 $Y=2.565
+ $X2=2.88 $Y2=2.565
r197 64 74 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.485 $Y=2.565
+ $X2=5.63 $Y2=2.565
r198 64 65 2.36869 $w=1.7e-07 $l=2.46e-06 $layer=MET1_cond $X=5.485 $Y=2.565
+ $X2=3.025 $Y2=2.565
r199 63 67 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.03 $Y=2.565
+ $X2=1.885 $Y2=2.565
r200 62 70 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.735 $Y=2.565
+ $X2=2.88 $Y2=2.565
r201 62 63 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=2.735 $Y=2.565
+ $X2=2.03 $Y2=2.565
r202 58 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.63 $Y=2.565
+ $X2=5.63 $Y2=2.565
r203 55 58 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.63 $Y=2.36
+ $X2=5.63 $Y2=2.565
r204 49 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.88 $Y=2.565
+ $X2=2.88 $Y2=2.565
r205 49 52 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.88 $Y=2.565
+ $X2=2.88 $Y2=2.74
r206 43 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.885 $Y=2.565
+ $X2=1.885 $Y2=2.565
r207 43 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.885 $Y=2.565
+ $X2=1.885 $Y2=2.74
r208 39 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=2.36 $X2=5.63 $Y2=2.36
r209 39 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=2.36
+ $X2=5.63 $Y2=2.525
r210 39 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=2.36
+ $X2=5.63 $Y2=2.195
r211 37 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=2.74 $X2=2.88 $Y2=2.74
r212 34 35 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.762 $Y=1.64
+ $X2=2.762 $Y2=1.79
r213 31 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=2.74 $X2=1.885 $Y2=2.74
r214 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=2.74
+ $X2=1.885 $Y2=2.905
r215 31 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=2.74
+ $X2=1.885 $Y2=2.575
r216 28 41 1043.48 $w=1.5e-07 $l=2.035e-06 $layer=POLY_cond $X=5.585 $Y=4.56
+ $X2=5.585 $Y2=2.525
r217 24 40 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=5.585 $Y=1.05
+ $X2=5.585 $Y2=2.195
r218 21 37 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=2.79 $Y=2.575
+ $X2=2.837 $Y2=2.74
r219 21 35 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.79 $Y=2.575
+ $X2=2.79 $Y2=1.79
r220 16 37 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=2.735 $Y=2.905
+ $X2=2.837 $Y2=2.74
r221 16 18 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.735 $Y=2.905
+ $X2=2.735 $Y2=4.56
r222 15 34 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.735 $Y=1.05
+ $X2=2.735 $Y2=1.64
r223 11 33 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.945 $Y=4.56
+ $X2=1.945 $Y2=2.905
r224 7 32 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.825 $Y=2.35
+ $X2=1.825 $Y2=2.575
r225 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.75 $Y=2.275
+ $X2=1.825 $Y2=2.35
r226 5 6 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.75 $Y=2.275
+ $X2=1.42 $Y2=2.275
r227 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=2.2
+ $X2=1.42 $Y2=2.275
r228 1 3 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=1.345 $Y=2.2
+ $X2=1.345 $Y2=1.05
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_43_110# 1 3 11 15 23 26 28 32 33 35
+ 36 37 38 42 45 49 54 59 65 68 73 74 78 81 83
c173 81 0 1.2087e-19 $X=2.22 $Y=2.195
c174 74 0 1.86741e-19 $X=2.515 $Y=2.195
c175 37 0 8.77106e-20 $X=3.75 $Y=2.83
c176 32 0 2.20611e-19 $X=3.66 $Y=2.195
r177 80 81 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.365 $Y=2.195
+ $X2=2.22 $Y2=2.195
r178 78 81 2.2896 $w=1.4e-07 $l=1.85e-06 $layer=MET1_cond $X=0.37 $Y=2.175
+ $X2=2.22 $Y2=2.175
r179 76 78 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.225 $Y=2.195
+ $X2=0.37 $Y2=2.195
r180 74 80 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=2.515 $Y=2.195
+ $X2=2.365 $Y2=2.195
r181 73 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.515 $Y=2.195
+ $X2=3.66 $Y2=2.195
r182 73 74 1.23762 $w=1.4e-07 $l=1e-06 $layer=MET1_cond $X=3.515 $Y=2.195
+ $X2=2.515 $Y2=2.195
r183 68 70 8.33135 $w=2.83e-07 $l=1.6e-07 $layer=LI1_cond $X=0.282 $Y=3.77
+ $X2=0.282 $Y2=3.93
r184 68 69 12.1728 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.282 $Y=3.77
+ $X2=0.282 $Y2=3.515
r185 63 65 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.225 $Y=1.37
+ $X2=0.34 $Y2=1.37
r186 59 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.66 $Y=2.195
+ $X2=3.66 $Y2=2.195
r187 54 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.365 $Y=2.195
+ $X2=2.365 $Y2=2.195
r188 49 51 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.34 $Y=4.11
+ $X2=0.34 $Y2=5.81
r189 49 70 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.34 $Y=4.11
+ $X2=0.34 $Y2=3.93
r190 43 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=1.285
+ $X2=0.34 $Y2=1.37
r191 43 45 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.34 $Y=1.285
+ $X2=0.34 $Y2=0.8
r192 42 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.225 $Y=2.195
+ $X2=0.225 $Y2=2.195
r193 42 69 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.225 $Y=2.195
+ $X2=0.225 $Y2=3.515
r194 39 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=1.455
+ $X2=0.225 $Y2=1.37
r195 39 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.225 $Y=1.455
+ $X2=0.225 $Y2=2.195
r196 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.75 $Y=2.83 $X2=3.75
+ $Y2=2.98
r197 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.75 $Y=1.625
+ $X2=3.75 $Y2=1.775
r198 34 37 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.725 $Y=2.36 $X2=3.725
+ $Y2=2.83
r199 33 36 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.725 $Y=2.03
+ $X2=3.725 $Y2=1.775
r200 32 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=2.195 $X2=3.66 $Y2=2.195
r201 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.662 $Y=2.195
+ $X2=3.662 $Y2=2.36
r202 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.662 $Y=2.195
+ $X2=3.662 $Y2=2.03
r203 28 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=2.195 $X2=2.365 $Y2=2.195
r204 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=2.195
+ $X2=2.365 $Y2=2.36
r205 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=2.195
+ $X2=2.365 $Y2=2.03
r206 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=3.775 $Y=4.56
+ $X2=3.775 $Y2=2.98
r207 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.775 $Y=1.05
+ $X2=3.775 $Y2=1.625
r208 15 30 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=2.305 $Y=4.56
+ $X2=2.305 $Y2=2.36
r209 11 29 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.305 $Y=1.05
+ $X2=2.305 $Y2=2.03
r210 3 51 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.215
+ $Y=3.06 $X2=0.34 $Y2=5.81
r211 3 49 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.215
+ $Y=3.06 $X2=0.34 $Y2=4.11
r212 3 68 600 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=3.06 $X2=0.34 $Y2=3.77
r213 1 45 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.55 $X2=0.34 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_687_110# 1 3 11 15 19 23 26 32 36 40
+ 46 47 48 49 53 55 60 61
c122 61 0 8.77106e-20 $X=3.705 $Y=2.935
c123 48 0 1.02575e-19 $X=4.06 $Y=2.74
c124 46 0 1.18035e-19 $X=4.06 $Y=1.825
c125 26 0 1.97615e-19 $X=4.145 $Y=2.195
r126 61 63 0.0909841 $w=2.11e-07 $l=1.45e-07 $layer=MET1_cond $X=3.705 $Y=2.935
+ $X2=3.56 $Y2=2.935
r127 60 65 0.0905464 $w=2.13e-07 $l=1.45e-07 $layer=MET1_cond $X=4.805 $Y=2.935
+ $X2=4.95 $Y2=2.935
r128 60 61 1.05917 $w=1.7e-07 $l=1.1e-06 $layer=MET1_cond $X=4.805 $Y=2.935
+ $X2=3.705 $Y2=2.935
r129 58 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.95 $Y=2.935
+ $X2=4.95 $Y2=2.935
r130 55 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.95 $Y=2.65
+ $X2=4.95 $Y2=2.935
r131 51 53 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.145 $Y=2.655
+ $X2=4.145 $Y2=2.195
r132 50 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.145 $Y=1.91
+ $X2=4.145 $Y2=2.195
r133 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=2.74
+ $X2=4.145 $Y2=2.655
r134 48 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.06 $Y=2.74
+ $X2=3.645 $Y2=2.74
r135 46 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=1.825
+ $X2=4.145 $Y2=1.91
r136 46 47 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.06 $Y=1.825
+ $X2=3.645 $Y2=1.825
r137 42 44 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.56 $Y=3.43
+ $X2=3.56 $Y2=5.81
r138 40 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.56 $Y=2.935
+ $X2=3.56 $Y2=2.935
r139 40 42 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.56 $Y=2.935
+ $X2=3.56 $Y2=3.43
r140 38 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=2.825
+ $X2=3.645 $Y2=2.74
r141 38 40 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.56 $Y=2.825
+ $X2=3.56 $Y2=2.935
r142 34 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=1.74
+ $X2=3.645 $Y2=1.825
r143 34 36 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.56 $Y=1.74
+ $X2=3.56 $Y2=0.8
r144 30 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.95
+ $Y=2.65 $X2=4.95 $Y2=2.65
r145 30 32 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.95 $Y=2.65
+ $X2=5.155 $Y2=2.65
r146 26 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=2.195 $X2=4.145 $Y2=2.195
r147 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.145 $Y=2.195
+ $X2=4.145 $Y2=2.36
r148 26 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.145 $Y=2.195
+ $X2=4.145 $Y2=2.03
r149 21 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=2.815
+ $X2=5.155 $Y2=2.65
r150 21 23 894.777 $w=1.5e-07 $l=1.745e-06 $layer=POLY_cond $X=5.155 $Y=2.815
+ $X2=5.155 $Y2=4.56
r151 17 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=2.485
+ $X2=5.155 $Y2=2.65
r152 17 19 735.819 $w=1.5e-07 $l=1.435e-06 $layer=POLY_cond $X=5.155 $Y=2.485
+ $X2=5.155 $Y2=1.05
r153 15 28 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=4.205 $Y=4.56
+ $X2=4.205 $Y2=2.36
r154 11 27 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.205 $Y=1.05
+ $X2=4.205 $Y2=2.03
r155 3 44 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=3.435
+ $Y=3.06 $X2=3.56 $Y2=5.81
r156 3 42 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=3.435
+ $Y=3.06 $X2=3.56 $Y2=3.43
r157 1 36 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.55 $X2=3.56 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_963_612# 1 3 11 15 16 18 19 24 28 29
+ 31 34 38 40
r80 36 40 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.455 $Y=1.91
+ $X2=5.33 $Y2=1.91
r81 36 38 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.455 $Y=1.91
+ $X2=6.11 $Y2=1.91
r82 32 40 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.37 $Y=1.825
+ $X2=5.33 $Y2=1.91
r83 32 34 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=5.37 $Y=1.825
+ $X2=5.37 $Y2=0.8
r84 30 40 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.29 $Y=1.995
+ $X2=5.33 $Y2=1.91
r85 30 31 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=5.29 $Y=1.995
+ $X2=5.29 $Y2=3.52
r86 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.205 $Y=3.605
+ $X2=5.29 $Y2=3.52
r87 28 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.205 $Y=3.605
+ $X2=5.025 $Y2=3.605
r88 24 26 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.94 $Y=3.77
+ $X2=4.94 $Y2=5.81
r89 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.94 $Y=3.69
+ $X2=5.025 $Y2=3.605
r90 22 24 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.94 $Y=3.69 $X2=4.94
+ $Y2=3.77
r91 21 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.91 $X2=6.11 $Y2=1.91
r92 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=6.032 $Y=2.785
+ $X2=6.032 $Y2=2.935
r93 16 21 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=6.05 $Y=2.075
+ $X2=6.092 $Y2=1.91
r94 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.05 $Y=2.075
+ $X2=6.05 $Y2=2.785
r95 15 19 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=6.015 $Y=4.56
+ $X2=6.015 $Y2=2.935
r96 9 21 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=6.015 $Y=1.745
+ $X2=6.092 $Y2=1.91
r97 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.015 $Y=1.745
+ $X2=6.015 $Y2=1.05
r98 3 26 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=4.815
+ $Y=3.06 $X2=4.94 $Y2=5.81
r99 3 24 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=4.815
+ $Y=3.06 $X2=4.94 $Y2=3.77
r100 1 34 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.55 $X2=5.37 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_856_110# 1 3 11 15 17 24 25
r32 24 25 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=4.485 $Y=1.57
+ $X2=4.485 $Y2=3.135
r33 23 24 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.452 $Y=1.4
+ $X2=4.452 $Y2=1.57
r34 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.42 $Y=3.43
+ $X2=4.42 $Y2=5.81
r35 15 25 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.452 $Y=3.305
+ $X2=4.452 $Y2=3.135
r36 15 17 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.42 $Y=3.305
+ $X2=4.42 $Y2=3.43
r37 11 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.42 $Y=0.8 $X2=4.42
+ $Y2=1.4
r38 3 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.28
+ $Y=3.06 $X2=4.42 $Y2=5.81
r39 3 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.28
+ $Y=3.06 $X2=4.42 $Y2=3.43
r40 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.28
+ $Y=0.55 $X2=4.42 $Y2=0.8
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NCGATE_1%ECK 1 3 10 16 24 26 29
c36 29 0 8.03558e-20 $X=6.23 $Y=2.565
r37 24 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=6.23 $Y=2.45
+ $X2=6.23 $Y2=2.565
r38 23 26 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=6.23 $Y=1.57
+ $X2=6.23 $Y2=1.455
r39 23 24 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=6.23 $Y=1.57
+ $X2=6.23 $Y2=2.45
r40 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.23 $Y=3.43
+ $X2=6.23 $Y2=5.81
r41 16 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.23 $Y=2.565
+ $X2=6.23 $Y2=2.565
r42 16 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.23 $Y=2.565
+ $X2=6.23 $Y2=3.43
r43 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.23 $Y=1.455
+ $X2=6.23 $Y2=1.455
r44 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.23 $Y=0.8
+ $X2=6.23 $Y2=1.455
r45 3 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.09
+ $Y=3.06 $X2=6.23 $Y2=5.81
r46 3 19 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.09
+ $Y=3.06 $X2=6.23 $Y2=3.43
r47 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.09
+ $Y=0.55 $X2=6.23 $Y2=0.8
.ends

