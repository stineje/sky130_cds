* File: sky130_osu_sc_18T_ms__tnbufi_l.pxi.spice
* Created: Thu Oct 29 17:32:02 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_5_p
+ N_GND_c_2_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%GND
x_PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%VDD N_VDD_M1005_d N_VDD_M1005_b N_VDD_c_33_p
+ N_VDD_c_38_p VDD N_VDD_c_34_p N_VDD_c_43_p
+ PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%VDD
x_PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1005_s N_A_27_115#_M1000_g N_A_27_115#_c_57_n N_A_27_115#_c_60_n
+ N_A_27_115#_c_61_n N_A_27_115#_c_62_n N_A_27_115#_c_63_n N_A_27_115#_c_64_n
+ PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%A_27_115#
x_PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%OE N_OE_M1002_g N_OE_c_101_n N_OE_M1005_g
+ N_OE_M1003_g N_OE_c_102_n OE N_OE_c_104_n PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%OE
x_PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%A N_A_M1004_g N_A_M1001_g N_A_c_146_n
+ N_A_c_147_n A N_A_c_148_n PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%A
x_PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%Y N_Y_M1004_d N_Y_M1001_d Y N_Y_c_191_n
+ N_Y_c_192_n N_Y_c_193_n N_Y_c_194_n PM_SKY130_OSU_SC_18T_MS__TNBUFI_L%Y
cc_1 N_GND_M1002_b N_A_27_115#_M1000_g 0.053782f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.945
cc_2 N_GND_c_2_p N_A_27_115#_M1000_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=0.945
cc_3 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.905
+ $Y2=0.945
cc_4 N_GND_M1002_b N_A_27_115#_c_57_n 0.0321466f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_5 N_GND_c_5_p N_A_27_115#_c_57_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_6 N_GND_c_3_p N_A_27_115#_c_57_n 0.00476261f $X=1.02 $Y=0.17 $X2=0.26
+ $Y2=0.825
cc_7 N_GND_M1002_b N_A_27_115#_c_60_n 0.0221237f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=4.475
cc_8 N_GND_M1002_b N_A_27_115#_c_61_n 0.00872418f $X=-0.045 $Y=0 $X2=0.605
+ $Y2=2.175
cc_9 N_GND_M1002_b N_A_27_115#_c_62_n 0.00647094f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.175
cc_10 N_GND_M1002_b N_A_27_115#_c_63_n 0.00739462f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=2.175
cc_11 N_GND_M1002_b N_A_27_115#_c_64_n 0.0434193f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=2.175
cc_12 N_GND_M1002_b N_OE_M1002_g 0.0333262f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_13 N_GND_c_5_p N_OE_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.945
cc_14 N_GND_c_2_p N_OE_M1002_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=0.945
cc_15 N_GND_c_3_p N_OE_M1002_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=0.945
cc_16 N_GND_M1002_b N_OE_c_101_n 0.102331f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.01
cc_17 N_GND_M1002_b N_OE_c_102_n 0.0253119f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.725
cc_18 N_GND_M1002_b OE 5.10551e-19 $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_19 N_GND_M1002_b N_OE_c_104_n 0.00123196f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.765
cc_20 N_GND_M1002_b N_A_M1004_g 0.0596037f $X=-0.045 $Y=0 $X2=1.265 $Y2=0.945
cc_21 N_GND_c_3_p N_A_M1004_g 0.00468827f $X=1.02 $Y=0.17 $X2=1.265 $Y2=0.945
cc_22 N_GND_M1002_b N_A_M1001_g 0.0426097f $X=-0.045 $Y=0 $X2=1.265 $Y2=5.085
cc_23 N_GND_M1002_b N_A_c_146_n 0.00872469f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.09
cc_24 N_GND_M1002_b N_A_c_147_n 0.031953f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.09
cc_25 N_GND_M1002_b N_A_c_148_n 0.0125638f $X=-0.045 $Y=0 $X2=1.14 $Y2=3.33
cc_26 N_GND_M1002_b Y 0.0395158f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.82
cc_27 N_GND_M1002_b N_Y_c_191_n 0.0157993f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.48
cc_28 N_GND_M1002_b N_Y_c_192_n 0.0157299f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.59
cc_29 N_GND_M1002_b N_Y_c_193_n 0.0151339f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.59
cc_30 N_GND_M1002_b N_Y_c_194_n 0.0196224f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.825
cc_31 N_GND_c_3_p N_Y_c_194_n 0.00476261f $X=1.02 $Y=0.17 $X2=1.48 $Y2=0.825
cc_32 N_VDD_M1005_b N_A_27_115#_c_60_n 0.0562932f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.475
cc_33 N_VDD_c_33_p N_A_27_115#_c_60_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=4.475
cc_34 N_VDD_c_34_p N_A_27_115#_c_60_n 0.00476261f $X=1.02 $Y=6.49 $X2=0.26
+ $Y2=4.475
cc_35 N_VDD_M1005_b N_OE_c_101_n 0.0237235f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=3.01
cc_36 N_VDD_M1005_b N_OE_M1005_g 0.0727196f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_37 N_VDD_c_33_p N_OE_M1005_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=5.085
cc_38 N_VDD_c_38_p N_OE_M1005_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.475 $Y2=5.085
cc_39 N_VDD_c_34_p N_OE_M1005_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=5.085
cc_40 N_VDD_M1005_b N_OE_M1003_g 0.0624108f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=5.085
cc_41 N_VDD_c_38_p N_OE_M1003_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.905 $Y2=5.085
cc_42 N_VDD_c_34_p N_OE_M1003_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.905 $Y2=5.085
cc_43 N_VDD_c_43_p N_OE_M1003_g 0.00606474f $X=1.02 $Y=6.44 $X2=0.905 $Y2=5.085
cc_44 N_VDD_M1005_b OE 0.0104205f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_45 N_VDD_M1005_b N_OE_c_104_n 0.00252354f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.765
cc_46 N_VDD_M1005_b N_A_M1001_g 0.0740659f $X=-0.045 $Y=2.905 $X2=1.265
+ $Y2=5.085
cc_47 N_VDD_c_34_p N_A_M1001_g 0.00468827f $X=1.02 $Y=6.49 $X2=1.265 $Y2=5.085
cc_48 N_VDD_c_43_p N_A_M1001_g 0.00606474f $X=1.02 $Y=6.44 $X2=1.265 $Y2=5.085
cc_49 N_VDD_M1005_b A 0.011498f $X=-0.045 $Y=2.905 $X2=1.14 $Y2=3.33
cc_50 N_VDD_M1005_b N_A_c_148_n 0.00640673f $X=-0.045 $Y=2.905 $X2=1.14 $Y2=3.33
cc_51 N_VDD_M1005_b N_Y_c_193_n 0.0577449f $X=-0.045 $Y=2.905 $X2=1.48 $Y2=2.59
cc_52 N_VDD_c_34_p N_Y_c_193_n 0.00476261f $X=1.02 $Y=6.49 $X2=1.48 $Y2=2.59
cc_53 N_VDD_c_43_p N_Y_c_193_n 0.00757793f $X=1.02 $Y=6.44 $X2=1.48 $Y2=2.59
cc_54 N_A_27_115#_M1000_g N_OE_M1002_g 0.0425033f $X=0.905 $Y=0.945 $X2=0.475
+ $Y2=0.945
cc_55 N_A_27_115#_c_57_n N_OE_M1002_g 0.0196674f $X=0.26 $Y=0.825 $X2=0.475
+ $Y2=0.945
cc_56 N_A_27_115#_M1000_g N_OE_c_101_n 0.00301188f $X=0.905 $Y=0.945 $X2=0.475
+ $Y2=3.01
cc_57 N_A_27_115#_c_57_n N_OE_c_101_n 0.0121188f $X=0.26 $Y=0.825 $X2=0.475
+ $Y2=3.01
cc_58 N_A_27_115#_c_60_n N_OE_c_101_n 0.04195f $X=0.26 $Y=4.475 $X2=0.475
+ $Y2=3.01
cc_59 N_A_27_115#_c_61_n N_OE_c_101_n 0.00111679f $X=0.605 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_60 N_A_27_115#_c_62_n N_OE_c_101_n 0.00632922f $X=0.26 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_61 N_A_27_115#_c_63_n N_OE_c_101_n 7.56328e-19 $X=0.69 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_62 N_A_27_115#_c_64_n N_OE_c_101_n 0.0400875f $X=0.905 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_63 N_A_27_115#_c_60_n N_OE_M1005_g 0.0459271f $X=0.26 $Y=4.475 $X2=0.475
+ $Y2=5.085
cc_64 N_A_27_115#_c_57_n N_OE_c_102_n 0.0104429f $X=0.26 $Y=0.825 $X2=0.475
+ $Y2=1.725
cc_65 N_A_27_115#_c_61_n N_OE_c_102_n 0.00711711f $X=0.605 $Y=2.175 $X2=0.475
+ $Y2=1.725
cc_66 N_A_27_115#_c_60_n OE 0.00651113f $X=0.26 $Y=4.475 $X2=0.69 $Y2=2.96
cc_67 N_A_27_115#_c_61_n OE 0.00158904f $X=0.605 $Y=2.175 $X2=0.69 $Y2=2.96
cc_68 N_A_27_115#_c_63_n OE 7.36678e-19 $X=0.69 $Y=2.175 $X2=0.69 $Y2=2.96
cc_69 N_A_27_115#_c_64_n OE 0.00125736f $X=0.905 $Y=2.175 $X2=0.69 $Y2=2.96
cc_70 N_A_27_115#_c_60_n N_OE_c_104_n 0.0193056f $X=0.26 $Y=4.475 $X2=0.69
+ $Y2=2.765
cc_71 N_A_27_115#_c_63_n N_OE_c_104_n 0.00847614f $X=0.69 $Y=2.175 $X2=0.69
+ $Y2=2.765
cc_72 N_A_27_115#_c_64_n N_OE_c_104_n 2.15234e-19 $X=0.905 $Y=2.175 $X2=0.69
+ $Y2=2.765
cc_73 N_A_27_115#_M1000_g N_A_M1004_g 0.0586829f $X=0.905 $Y=0.945 $X2=1.265
+ $Y2=0.945
cc_74 N_A_27_115#_M1000_g N_A_c_146_n 0.00160395f $X=0.905 $Y=0.945 $X2=1.325
+ $Y2=2.09
cc_75 N_A_27_115#_c_63_n N_A_c_146_n 0.00878007f $X=0.69 $Y=2.175 $X2=1.325
+ $Y2=2.09
cc_76 N_A_27_115#_c_63_n N_A_c_147_n 2.55709e-19 $X=0.69 $Y=2.175 $X2=1.325
+ $Y2=2.09
cc_77 N_A_27_115#_c_64_n N_A_c_147_n 0.0586829f $X=0.905 $Y=2.175 $X2=1.325
+ $Y2=2.09
cc_78 N_A_27_115#_c_60_n A 0.00539687f $X=0.26 $Y=4.475 $X2=1.14 $Y2=3.33
cc_79 N_A_27_115#_c_63_n N_A_c_148_n 0.00813625f $X=0.69 $Y=2.175 $X2=1.14
+ $Y2=3.33
cc_80 N_A_27_115#_c_64_n N_A_c_148_n 0.00134082f $X=0.905 $Y=2.175 $X2=1.14
+ $Y2=3.33
cc_81 N_A_27_115#_M1000_g Y 3.32545e-19 $X=0.905 $Y=0.945 $X2=1.525 $Y2=1.82
cc_82 N_A_27_115#_M1000_g N_Y_c_191_n 0.00101819f $X=0.905 $Y=0.945 $X2=1.48
+ $Y2=1.48
cc_83 N_OE_c_101_n N_A_M1001_g 0.20929f $X=0.475 $Y=3.01 $X2=1.265 $Y2=5.085
cc_84 N_OE_c_104_n N_A_M1001_g 4.61952e-19 $X=0.69 $Y=2.765 $X2=1.265 $Y2=5.085
cc_85 N_OE_M1005_g A 8.46663e-19 $X=0.475 $Y=5.085 $X2=1.14 $Y2=3.33
cc_86 N_OE_M1003_g A 0.0104662f $X=0.905 $Y=5.085 $X2=1.14 $Y2=3.33
cc_87 OE A 0.004991f $X=0.69 $Y=2.96 $X2=1.14 $Y2=3.33
cc_88 N_OE_c_101_n N_A_c_148_n 0.0110152f $X=0.475 $Y=3.01 $X2=1.14 $Y2=3.33
cc_89 OE N_A_c_148_n 0.007197f $X=0.69 $Y=2.96 $X2=1.14 $Y2=3.33
cc_90 N_OE_c_104_n N_A_c_148_n 0.0187675f $X=0.69 $Y=2.765 $X2=1.14 $Y2=3.33
cc_91 N_A_M1004_g Y 0.00768908f $X=1.265 $Y=0.945 $X2=1.525 $Y2=1.82
cc_92 N_A_M1001_g Y 0.00511826f $X=1.265 $Y=5.085 $X2=1.525 $Y2=1.82
cc_93 N_A_c_146_n Y 0.0130872f $X=1.325 $Y=2.09 $X2=1.525 $Y2=1.82
cc_94 N_A_c_147_n Y 0.00539093f $X=1.325 $Y=2.09 $X2=1.525 $Y2=1.82
cc_95 N_A_c_148_n Y 0.012418f $X=1.14 $Y=3.33 $X2=1.525 $Y2=1.82
cc_96 N_A_M1004_g N_Y_c_191_n 0.00707709f $X=1.265 $Y=0.945 $X2=1.48 $Y2=1.48
cc_97 N_A_c_146_n N_Y_c_191_n 0.00203451f $X=1.325 $Y=2.09 $X2=1.48 $Y2=1.48
cc_98 N_A_c_147_n N_Y_c_191_n 0.00129509f $X=1.325 $Y=2.09 $X2=1.48 $Y2=1.48
cc_99 N_A_M1001_g N_Y_c_192_n 0.00489736f $X=1.265 $Y=5.085 $X2=1.48 $Y2=2.59
cc_100 N_A_c_146_n N_Y_c_192_n 0.00227834f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_101 N_A_c_147_n N_Y_c_192_n 0.00138163f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_102 N_A_c_148_n N_Y_c_192_n 0.00656407f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_103 N_A_M1001_g N_Y_c_193_n 0.0501139f $X=1.265 $Y=5.085 $X2=1.48 $Y2=2.59
cc_104 N_A_c_146_n N_Y_c_193_n 0.00330615f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_105 N_A_c_147_n N_Y_c_193_n 0.00102058f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_106 A N_Y_c_193_n 0.00706656f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_107 N_A_c_148_n N_Y_c_193_n 0.0606572f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_108 N_A_M1004_g N_Y_c_194_n 0.0152627f $X=1.265 $Y=0.945 $X2=1.48 $Y2=0.825
cc_109 N_A_c_146_n N_Y_c_194_n 0.00231567f $X=1.325 $Y=2.09 $X2=1.48 $Y2=0.825
cc_110 N_A_c_147_n N_Y_c_194_n 8.70049e-19 $X=1.325 $Y=2.09 $X2=1.48 $Y2=0.825
