* File: sky130_osu_sc_18T_hs__ant.pxi.spice
* Created: Thu Oct 29 17:06:22 2020
* 
x_PM_SKY130_OSU_SC_18T_HS__ANT%GND N_GND_M1001_b GND
+ PM_SKY130_OSU_SC_18T_HS__ANT%GND
x_PM_SKY130_OSU_SC_18T_HS__ANT%VDD N_VDD_M1000_d N_VDD_M1000_b N_VDD_c_15_p
+ N_VDD_c_16_p VDD PM_SKY130_OSU_SC_18T_HS__ANT%VDD
x_PM_SKY130_OSU_SC_18T_HS__ANT%A N_A_M1001_s N_A_M1000_s N_A_M1001_g N_A_M1000_g
+ N_A_c_23_n N_A_c_25_n N_A_c_26_n N_A_c_27_n N_A_c_28_n N_A_c_30_n A N_A_c_32_n
+ N_A_c_33_n PM_SKY130_OSU_SC_18T_HS__ANT%A
cc_1 N_GND_M1001_b N_A_M1001_g 0.0850747f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_M1001_b N_A_M1000_g 0.0125577f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_3 N_GND_M1001_b N_A_c_23_n 0.0236328f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.825
cc_4 GND N_A_c_23_n 0.00138205f $X=0.34 $Y=0.22 $X2=0.26 $Y2=0.825
cc_5 N_GND_M1001_b N_A_c_25_n 0.0149833f $X=-0.045 $Y=0 $X2=0.26 $Y2=2.505
cc_6 N_GND_M1001_b N_A_c_26_n 0.00651531f $X=-0.045 $Y=0 $X2=0.26 $Y2=3.455
cc_7 N_GND_M1001_b N_A_c_27_n 0.0199494f $X=-0.045 $Y=0 $X2=0.605 $Y2=2
cc_8 N_GND_M1001_b N_A_c_28_n 0.0238485f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_9 GND N_A_c_28_n 0.00138205f $X=0.34 $Y=0.22 $X2=0.69 $Y2=0.825
cc_10 N_GND_M1001_b N_A_c_30_n 0.00710193f $X=-0.045 $Y=0 $X2=0.26 $Y2=2
cc_11 N_GND_M1001_b A 0.00241298f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.59
cc_12 N_GND_M1001_b N_A_c_32_n 0.0076399f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.59
cc_13 N_GND_M1001_b N_A_c_33_n 0.0562319f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.59
cc_14 N_VDD_M1000_b N_A_M1000_g 0.0299903f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_15 N_VDD_c_15_p N_A_M1000_g 0.00713292f $X=0.69 $Y=3.455 $X2=0.475 $Y2=4.585
cc_16 N_VDD_c_16_p N_A_M1000_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475 $Y2=4.585
cc_17 VDD N_A_M1000_g 0.00468827f $X=0.34 $Y=6.44 $X2=0.475 $Y2=4.585
cc_18 N_VDD_M1000_b N_A_c_26_n 0.0103018f $X=-0.045 $Y=2.905 $X2=0.26 $Y2=3.455
cc_19 N_VDD_c_16_p N_A_c_26_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26 $Y2=3.455
cc_20 VDD N_A_c_26_n 0.00476261f $X=0.34 $Y=6.44 $X2=0.26 $Y2=3.455
