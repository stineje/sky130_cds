* File: sky130_osu_sc_12T_hs__oai21_l.spice
* Created: Fri Nov 12 15:12:17 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__oai21_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__oai21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A0_M1004_g N_A_27_114#_M1004_s N_GND_M1004_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_A_27_114#_M1001_d N_A1_M1001_g N_GND_M1004_d N_GND_M1004_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_114#_M1001_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_A0_M1000_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.9 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A1_M1005_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.23814 AS=0.1323 PD=1.92 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_B0_M1003_g N_VDD_M1005_d N_VDD_M1000_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.15876 PD=2.21 PS=1.28 NRD=0 NRS=14.0658 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=3.9449 P=7.95
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__oai21_l.pxi.spice"
*
.ends
*
*
