* File: sky130_osu_sc_18T_hs__tbufi_l.pxi.spice
* Created: Thu Oct 29 17:10:09 2020
* 
x_PM_SKY130_OSU_SC_18T_HS__TBUFI_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_3_p
+ N_GND_c_4_p GND N_GND_c_5_p PM_SKY130_OSU_SC_18T_HS__TBUFI_L%GND
x_PM_SKY130_OSU_SC_18T_HS__TBUFI_L%VDD N_VDD_M1005_d N_VDD_M1005_b N_VDD_c_37_p
+ N_VDD_c_38_p VDD N_VDD_c_39_p N_VDD_c_45_p
+ PM_SKY130_OSU_SC_18T_HS__TBUFI_L%VDD
x_PM_SKY130_OSU_SC_18T_HS__TBUFI_L%OE N_OE_c_57_n N_OE_M1002_g N_OE_M1005_g
+ N_OE_M1000_g N_OE_c_65_n N_OE_c_66_n N_OE_c_67_n OE N_OE_c_69_n
+ PM_SKY130_OSU_SC_18T_HS__TBUFI_L%OE
x_PM_SKY130_OSU_SC_18T_HS__TBUFI_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1005_s N_A_27_115#_M1003_g N_A_27_115#_c_120_n
+ N_A_27_115#_c_123_n N_A_27_115#_c_124_n N_A_27_115#_c_125_n
+ N_A_27_115#_c_126_n N_A_27_115#_c_127_n
+ PM_SKY130_OSU_SC_18T_HS__TBUFI_L%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__TBUFI_L%A N_A_M1004_g N_A_M1001_g N_A_c_172_n
+ N_A_c_173_n A N_A_c_174_n PM_SKY130_OSU_SC_18T_HS__TBUFI_L%A
x_PM_SKY130_OSU_SC_18T_HS__TBUFI_L%Y N_Y_M1004_d N_Y_M1001_d Y N_Y_c_216_n
+ N_Y_c_217_n N_Y_c_218_n N_Y_c_219_n PM_SKY130_OSU_SC_18T_HS__TBUFI_L%Y
cc_1 N_GND_M1002_b N_OE_c_57_n 0.0680245f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.86
cc_2 N_GND_M1002_b N_OE_M1002_g 0.0325412f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_OE_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.945
cc_4 N_GND_c_4_p N_OE_M1002_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=0.945
cc_5 N_GND_c_5_p N_OE_M1002_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=0.945
cc_6 N_GND_M1002_b N_OE_M1000_g 0.0329486f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.945
cc_7 N_GND_c_4_p N_OE_M1000_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905 $Y2=0.945
cc_8 N_GND_c_5_p N_OE_M1000_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.905 $Y2=0.945
cc_9 N_GND_M1002_b N_OE_c_65_n 0.00923524f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.935
cc_10 N_GND_M1002_b N_OE_c_66_n 7.18349e-19 $X=-0.045 $Y=0 $X2=0.69 $Y2=1.85
cc_11 N_GND_M1002_b N_OE_c_67_n 0.00260472f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.85
cc_12 N_GND_M1002_b OE 0.0107998f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_13 N_GND_M1002_b N_OE_c_69_n 0.0553909f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.85
cc_14 N_GND_c_4_p N_OE_c_69_n 0.00294633f $X=0.69 $Y=0.825 $X2=0.69 $Y2=1.85
cc_15 N_GND_M1002_b N_A_27_115#_M1003_g 0.014739f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=5.085
cc_16 N_GND_M1002_b N_A_27_115#_c_120_n 0.0426244f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_17 N_GND_c_3_p N_A_27_115#_c_120_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_18 N_GND_c_5_p N_A_27_115#_c_120_n 0.00476261f $X=1.02 $Y=0.17 $X2=0.26
+ $Y2=0.825
cc_19 N_GND_M1002_b N_A_27_115#_c_123_n 0.0116459f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=4.475
cc_20 N_GND_M1002_b N_A_27_115#_c_124_n 0.0101855f $X=-0.045 $Y=0 $X2=0.715
+ $Y2=2.48
cc_21 N_GND_M1002_b N_A_27_115#_c_125_n 0.00665288f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.48
cc_22 N_GND_M1002_b N_A_27_115#_c_126_n 0.00288071f $X=-0.045 $Y=0 $X2=0.8
+ $Y2=2.48
cc_23 N_GND_M1002_b N_A_27_115#_c_127_n 0.0326306f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=2.48
cc_24 N_GND_M1002_b N_A_M1004_g 0.0603023f $X=-0.045 $Y=0 $X2=1.265 $Y2=0.945
cc_25 N_GND_c_5_p N_A_M1004_g 0.00468827f $X=1.02 $Y=0.17 $X2=1.265 $Y2=0.945
cc_26 N_GND_M1002_b N_A_M1001_g 0.0372976f $X=-0.045 $Y=0 $X2=1.265 $Y2=5.085
cc_27 N_GND_M1002_b N_A_c_172_n 0.00983127f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.09
cc_28 N_GND_M1002_b N_A_c_173_n 0.0369358f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.09
cc_29 N_GND_M1002_b N_A_c_174_n 0.00459479f $X=-0.045 $Y=0 $X2=1.14 $Y2=3.33
cc_30 N_GND_M1002_b Y 0.0383474f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.82
cc_31 N_GND_M1002_b N_Y_c_216_n 0.0157993f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.48
cc_32 N_GND_M1002_b N_Y_c_217_n 0.0157299f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.59
cc_33 N_GND_M1002_b N_Y_c_218_n 0.0151339f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.59
cc_34 N_GND_M1002_b N_Y_c_219_n 0.0196224f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.825
cc_35 N_GND_c_5_p N_Y_c_219_n 0.00476261f $X=1.02 $Y=0.17 $X2=1.48 $Y2=0.825
cc_36 N_VDD_M1005_b N_OE_M1005_g 0.0746788f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_37 N_VDD_c_37_p N_OE_M1005_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=5.085
cc_38 N_VDD_c_38_p N_OE_M1005_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.475 $Y2=5.085
cc_39 N_VDD_c_39_p N_OE_M1005_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=5.085
cc_40 N_VDD_M1005_b N_OE_c_65_n 0.0152497f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.935
cc_41 N_VDD_M1005_b OE 0.0109902f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_42 N_VDD_M1005_b N_A_27_115#_M1003_g 0.0692342f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=5.085
cc_43 N_VDD_c_38_p N_A_27_115#_M1003_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.905
+ $Y2=5.085
cc_44 N_VDD_c_39_p N_A_27_115#_M1003_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.905
+ $Y2=5.085
cc_45 N_VDD_c_45_p N_A_27_115#_M1003_g 0.00606474f $X=1.02 $Y=6.44 $X2=0.905
+ $Y2=5.085
cc_46 N_VDD_M1005_b N_A_27_115#_c_123_n 0.0562104f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.475
cc_47 N_VDD_c_37_p N_A_27_115#_c_123_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=4.475
cc_48 N_VDD_c_39_p N_A_27_115#_c_123_n 0.00476261f $X=1.02 $Y=6.49 $X2=0.26
+ $Y2=4.475
cc_49 N_VDD_M1005_b N_A_M1001_g 0.0740659f $X=-0.045 $Y=2.905 $X2=1.265
+ $Y2=5.085
cc_50 N_VDD_c_39_p N_A_M1001_g 0.00468827f $X=1.02 $Y=6.49 $X2=1.265 $Y2=5.085
cc_51 N_VDD_c_45_p N_A_M1001_g 0.00606474f $X=1.02 $Y=6.44 $X2=1.265 $Y2=5.085
cc_52 N_VDD_M1005_b A 0.011498f $X=-0.045 $Y=2.905 $X2=1.14 $Y2=3.33
cc_53 N_VDD_M1005_b N_A_c_174_n 0.00605669f $X=-0.045 $Y=2.905 $X2=1.14 $Y2=3.33
cc_54 N_VDD_M1005_b N_Y_c_218_n 0.0577449f $X=-0.045 $Y=2.905 $X2=1.48 $Y2=2.59
cc_55 N_VDD_c_39_p N_Y_c_218_n 0.00476261f $X=1.02 $Y=6.49 $X2=1.48 $Y2=2.59
cc_56 N_VDD_c_45_p N_Y_c_218_n 0.00757793f $X=1.02 $Y=6.44 $X2=1.48 $Y2=2.59
cc_57 N_OE_c_57_n N_A_27_115#_M1003_g 0.00266681f $X=0.27 $Y=2.86 $X2=0.905
+ $Y2=5.085
cc_58 N_OE_c_65_n N_A_27_115#_M1003_g 0.0710901f $X=0.475 $Y=2.935 $X2=0.905
+ $Y2=5.085
cc_59 OE N_A_27_115#_M1003_g 0.0135769f $X=0.69 $Y=2.96 $X2=0.905 $Y2=5.085
cc_60 N_OE_c_57_n N_A_27_115#_c_120_n 0.0232517f $X=0.27 $Y=2.86 $X2=0.26
+ $Y2=0.825
cc_61 N_OE_M1002_g N_A_27_115#_c_120_n 0.0196674f $X=0.475 $Y=0.945 $X2=0.26
+ $Y2=0.825
cc_62 N_OE_c_66_n N_A_27_115#_c_120_n 0.00367353f $X=0.69 $Y=1.85 $X2=0.26
+ $Y2=0.825
cc_63 N_OE_c_67_n N_A_27_115#_c_120_n 0.0116068f $X=0.69 $Y=1.85 $X2=0.26
+ $Y2=0.825
cc_64 OE N_A_27_115#_c_120_n 0.015341f $X=0.69 $Y=2.96 $X2=0.26 $Y2=0.825
cc_65 N_OE_c_69_n N_A_27_115#_c_120_n 0.0135784f $X=0.69 $Y=1.85 $X2=0.26
+ $Y2=0.825
cc_66 N_OE_c_57_n N_A_27_115#_c_123_n 0.0103172f $X=0.27 $Y=2.86 $X2=0.26
+ $Y2=4.475
cc_67 N_OE_M1005_g N_A_27_115#_c_123_n 0.0464726f $X=0.475 $Y=5.085 $X2=0.26
+ $Y2=4.475
cc_68 N_OE_c_65_n N_A_27_115#_c_123_n 0.00887831f $X=0.475 $Y=2.935 $X2=0.26
+ $Y2=4.475
cc_69 OE N_A_27_115#_c_123_n 0.0193905f $X=0.69 $Y=2.96 $X2=0.26 $Y2=4.475
cc_70 N_OE_c_65_n N_A_27_115#_c_124_n 0.00703932f $X=0.475 $Y=2.935 $X2=0.715
+ $Y2=2.48
cc_71 N_OE_c_66_n N_A_27_115#_c_124_n 0.00123496f $X=0.69 $Y=1.85 $X2=0.715
+ $Y2=2.48
cc_72 N_OE_c_67_n N_A_27_115#_c_124_n 0.00456286f $X=0.69 $Y=1.85 $X2=0.715
+ $Y2=2.48
cc_73 OE N_A_27_115#_c_124_n 0.0142208f $X=0.69 $Y=2.96 $X2=0.715 $Y2=2.48
cc_74 N_OE_c_69_n N_A_27_115#_c_124_n 0.00292172f $X=0.69 $Y=1.85 $X2=0.715
+ $Y2=2.48
cc_75 N_OE_c_57_n N_A_27_115#_c_125_n 0.00700951f $X=0.27 $Y=2.86 $X2=0.26
+ $Y2=2.48
cc_76 N_OE_c_57_n N_A_27_115#_c_126_n 7.28524e-19 $X=0.27 $Y=2.86 $X2=0.8
+ $Y2=2.48
cc_77 N_OE_c_66_n N_A_27_115#_c_126_n 0.00129814f $X=0.69 $Y=1.85 $X2=0.8
+ $Y2=2.48
cc_78 N_OE_c_67_n N_A_27_115#_c_126_n 0.00377605f $X=0.69 $Y=1.85 $X2=0.8
+ $Y2=2.48
cc_79 OE N_A_27_115#_c_126_n 0.0157069f $X=0.69 $Y=2.96 $X2=0.8 $Y2=2.48
cc_80 N_OE_c_69_n N_A_27_115#_c_126_n 7.06691e-19 $X=0.69 $Y=1.85 $X2=0.8
+ $Y2=2.48
cc_81 N_OE_c_57_n N_A_27_115#_c_127_n 0.0126749f $X=0.27 $Y=2.86 $X2=0.905
+ $Y2=2.48
cc_82 N_OE_c_67_n N_A_27_115#_c_127_n 4.88301e-19 $X=0.69 $Y=1.85 $X2=0.905
+ $Y2=2.48
cc_83 OE N_A_27_115#_c_127_n 0.00242154f $X=0.69 $Y=2.96 $X2=0.905 $Y2=2.48
cc_84 N_OE_c_69_n N_A_27_115#_c_127_n 0.0119465f $X=0.69 $Y=1.85 $X2=0.905
+ $Y2=2.48
cc_85 N_OE_M1000_g N_A_M1004_g 0.0839097f $X=0.905 $Y=0.945 $X2=1.265 $Y2=0.945
cc_86 N_OE_c_67_n N_A_M1004_g 0.00287993f $X=0.69 $Y=1.85 $X2=1.265 $Y2=0.945
cc_87 N_OE_c_69_n N_A_M1004_g 0.00693622f $X=0.69 $Y=1.85 $X2=1.265 $Y2=0.945
cc_88 OE N_A_c_172_n 0.00765298f $X=0.69 $Y=2.96 $X2=1.325 $Y2=2.09
cc_89 N_OE_c_69_n N_A_c_172_n 2.20759e-19 $X=0.69 $Y=1.85 $X2=1.325 $Y2=2.09
cc_90 OE N_A_c_173_n 2.30744e-19 $X=0.69 $Y=2.96 $X2=1.325 $Y2=2.09
cc_91 N_OE_M1005_g A 8.46663e-19 $X=0.475 $Y=5.085 $X2=1.14 $Y2=3.33
cc_92 OE A 0.004991f $X=0.69 $Y=2.96 $X2=1.14 $Y2=3.33
cc_93 OE N_A_c_174_n 0.0257797f $X=0.69 $Y=2.96 $X2=1.14 $Y2=3.33
cc_94 N_OE_c_66_n Y 0.0105247f $X=0.69 $Y=1.85 $X2=1.525 $Y2=1.82
cc_95 N_OE_c_67_n Y 0.00375884f $X=0.69 $Y=1.85 $X2=1.525 $Y2=1.82
cc_96 N_OE_c_69_n Y 2.15427e-19 $X=0.69 $Y=1.85 $X2=1.525 $Y2=1.82
cc_97 N_OE_M1000_g N_Y_c_216_n 0.00101819f $X=0.905 $Y=0.945 $X2=1.48 $Y2=1.48
cc_98 OE N_Y_c_217_n 0.0100845f $X=0.69 $Y=2.96 $X2=1.48 $Y2=2.59
cc_99 N_A_27_115#_c_126_n N_A_M1001_g 2.80054e-19 $X=0.8 $Y=2.48 $X2=1.265
+ $Y2=5.085
cc_100 N_A_27_115#_c_127_n N_A_M1001_g 0.233224f $X=0.905 $Y=2.48 $X2=1.265
+ $Y2=5.085
cc_101 N_A_27_115#_M1003_g A 0.01062f $X=0.905 $Y=5.085 $X2=1.14 $Y2=3.33
cc_102 N_A_27_115#_c_123_n A 0.00539687f $X=0.26 $Y=4.475 $X2=1.14 $Y2=3.33
cc_103 N_A_27_115#_c_126_n N_A_c_174_n 0.0209392f $X=0.8 $Y=2.48 $X2=1.14
+ $Y2=3.33
cc_104 N_A_27_115#_c_127_n N_A_c_174_n 0.0186036f $X=0.905 $Y=2.48 $X2=1.14
+ $Y2=3.33
cc_105 N_A_M1004_g Y 0.00631192f $X=1.265 $Y=0.945 $X2=1.525 $Y2=1.82
cc_106 N_A_M1001_g Y 0.00511826f $X=1.265 $Y=5.085 $X2=1.525 $Y2=1.82
cc_107 N_A_c_172_n Y 0.0167787f $X=1.325 $Y=2.09 $X2=1.525 $Y2=1.82
cc_108 N_A_c_173_n Y 0.0051471f $X=1.325 $Y=2.09 $X2=1.525 $Y2=1.82
cc_109 N_A_c_174_n Y 0.012418f $X=1.14 $Y=3.33 $X2=1.525 $Y2=1.82
cc_110 N_A_M1004_g N_Y_c_216_n 0.00707709f $X=1.265 $Y=0.945 $X2=1.48 $Y2=1.48
cc_111 N_A_c_172_n N_Y_c_216_n 0.00203451f $X=1.325 $Y=2.09 $X2=1.48 $Y2=1.48
cc_112 N_A_c_173_n N_Y_c_216_n 0.00129509f $X=1.325 $Y=2.09 $X2=1.48 $Y2=1.48
cc_113 N_A_M1001_g N_Y_c_217_n 0.00445157f $X=1.265 $Y=5.085 $X2=1.48 $Y2=2.59
cc_114 N_A_c_172_n N_Y_c_217_n 0.00227834f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_115 N_A_c_173_n N_Y_c_217_n 0.00138163f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_116 N_A_c_174_n N_Y_c_217_n 0.0031919f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_117 N_A_M1001_g N_Y_c_218_n 0.0501139f $X=1.265 $Y=5.085 $X2=1.48 $Y2=2.59
cc_118 N_A_c_172_n N_Y_c_218_n 0.00330615f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_119 N_A_c_173_n N_Y_c_218_n 0.00102058f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_120 A N_Y_c_218_n 0.00706656f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_121 N_A_c_174_n N_Y_c_218_n 0.0606572f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_122 N_A_M1004_g N_Y_c_219_n 0.0152627f $X=1.265 $Y=0.945 $X2=1.48 $Y2=0.825
cc_123 N_A_c_172_n N_Y_c_219_n 0.00231567f $X=1.325 $Y=2.09 $X2=1.48 $Y2=0.825
cc_124 N_A_c_173_n N_Y_c_219_n 8.70049e-19 $X=1.325 $Y=2.09 $X2=1.48 $Y2=0.825
