magic
tech sky130A
magscale 1 2
timestamp 1612373489
<< nwell >>
rect -9 529 553 1119
<< nmoslvt >>
rect 80 115 110 243
rect 270 115 300 243
rect 356 115 386 243
<< pmos >>
rect 80 565 110 965
rect 270 565 300 965
rect 356 565 386 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 163 243
rect 110 131 121 215
rect 155 131 163 215
rect 110 115 163 131
rect 217 215 270 243
rect 217 131 225 215
rect 259 131 270 215
rect 217 115 270 131
rect 300 215 356 243
rect 300 131 311 215
rect 345 131 356 215
rect 300 115 356 131
rect 386 215 439 243
rect 386 131 397 215
rect 431 131 439 215
rect 386 115 439 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 949 163 965
rect 110 605 121 949
rect 155 605 163 949
rect 110 565 163 605
rect 217 949 270 965
rect 217 605 225 949
rect 259 605 270 949
rect 217 565 270 605
rect 300 949 356 965
rect 300 605 311 949
rect 345 605 356 949
rect 300 565 356 605
rect 386 949 439 965
rect 386 605 397 949
rect 431 605 439 949
rect 386 565 439 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 225 131 259 215
rect 311 131 345 215
rect 397 131 431 215
<< pdiffc >>
rect 35 741 69 949
rect 121 605 155 949
rect 225 605 259 949
rect 311 605 345 949
rect 397 605 431 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 435 1049 459 1083
rect 493 1049 517 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 459 1049 493 1083
<< poly >>
rect 80 980 300 1010
rect 80 965 110 980
rect 270 965 300 980
rect 356 965 386 991
rect 80 442 110 565
rect 270 539 300 565
rect 152 503 218 513
rect 152 469 168 503
rect 202 489 218 503
rect 356 489 386 565
rect 202 469 386 489
rect 152 459 386 469
rect 27 426 110 442
rect 27 392 37 426
rect 71 417 110 426
rect 71 392 386 417
rect 27 387 386 392
rect 27 376 110 387
rect 80 243 110 376
rect 152 335 218 345
rect 152 301 168 335
rect 202 321 218 335
rect 202 301 300 321
rect 152 291 300 301
rect 270 243 300 291
rect 356 243 386 387
rect 80 89 110 115
rect 270 89 300 115
rect 356 89 386 115
<< polycont >>
rect 168 469 202 503
rect 37 392 71 426
rect 168 301 202 335
<< locali >>
rect 0 1089 550 1110
rect 0 1049 459 1089
rect 493 1049 550 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 121 949 155 965
rect 37 426 71 597
rect 37 376 71 392
rect 121 519 155 605
rect 225 949 259 965
rect 311 949 345 965
rect 225 571 270 605
rect 236 557 270 571
rect 121 503 202 519
rect 121 469 168 503
rect 121 453 202 469
rect 121 351 155 453
rect 121 335 202 351
rect 121 301 168 335
rect 121 285 202 301
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 285
rect 236 249 270 523
rect 311 409 345 605
rect 397 949 431 965
rect 397 483 431 605
rect 121 115 155 131
rect 225 215 270 249
rect 311 215 345 227
rect 225 115 259 131
rect 311 115 345 131
rect 397 215 431 449
rect 397 115 431 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 550 61
rect 0 0 550 21
<< viali >>
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 37 597 71 631
rect 236 523 270 557
rect 311 375 345 409
rect 397 449 431 483
rect 311 227 345 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1089 550 1110
rect 0 1055 459 1089
rect 493 1055 550 1089
rect 0 1049 550 1055
rect 25 631 83 637
rect 25 597 37 631
rect 71 597 117 631
rect 25 591 83 597
rect 224 557 282 563
rect 190 523 236 557
rect 270 523 282 557
rect 224 517 282 523
rect 385 483 443 489
rect 351 449 397 483
rect 431 449 443 483
rect 385 443 443 449
rect 299 409 357 415
rect 299 375 311 409
rect 345 375 357 409
rect 299 369 357 375
rect 311 267 345 369
rect 299 261 357 267
rect 299 227 311 261
rect 345 227 357 261
rect 299 221 357 227
rect 0 55 550 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 550 55
rect 0 0 550 21
<< labels >>
rlabel viali 54 614 54 614 1 S0
port 1 n
rlabel viali 328 392 328 392 1 Y
port 2 n
rlabel viali 253 540 253 540 1 A0
port 3 n
rlabel viali 414 466 414 466 1 A1
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 476 1062 476 1062 1 vdd
<< end >>
