* File: sky130_osu_sc_15T_hs__tiehi.spice
* Created: Fri Nov 12 14:33:30 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__tiehi.pex.spice"
.subckt sky130_osu_sc_15T_hs__tiehi  GND VDD Y
* 
* Y	Y
* VDD	VDD
* GND	GND
MM1000 N_A_80_89#_M1000_d N_A_80_89#_M1000_g N_GND_M1000_s N_GND_M1000_b NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_Y_M1001_d N_A_80_89#_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX2_noxref N_GND_M1000_b N_VDD_M1001_b NWDIODE A=3.068 P=7.98
pX3_noxref noxref_5 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__tiehi.pxi.spice"
*
.ends
*
*
