* File: sky130_osu_sc_15T_ms__oai22_l.pex.spice
* Created: Fri Nov 12 14:45:43 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%GND 1 23 25 33 48 50
r46 48 50 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r47 35 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r48 31 44 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r49 31 33 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r50 25 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r51 23 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r52 23 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r53 23 35 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r54 23 25 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r55 1 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%VDD 1 2 21 25 29 38 49 53
r26 49 53 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.7 $Y2=5.397
r27 45 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r28 38 41 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.91 $Y=3.885
+ $X2=1.91 $Y2=4.565
r29 36 47 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.91 $Y=5.245
+ $X2=1.91 $Y2=5.397
r30 36 41 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.91 $Y=5.245
+ $X2=1.91 $Y2=4.565
r31 34 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=5.36 $X2=1.7
+ $Y2=5.36
r32 32 34 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=5.397
+ $X2=1.7 $Y2=5.397
r33 30 45 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r34 30 32 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r35 29 47 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=5.397
+ $X2=1.91 $Y2=5.397
r36 29 34 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=5.397
+ $X2=1.7 $Y2=5.397
r37 25 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r38 23 45 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r39 23 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r40 21 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r41 21 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r42 21 45 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r43 2 41 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=2.825 $X2=1.91 $Y2=4.565
r44 2 38 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=2.825 $X2=1.91 $Y2=3.885
r45 1 28 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r46 1 25 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%A0 3 5 8 12 15 16 19 25
r36 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.415 $Y=3.07
+ $X2=0.415 $Y2=3.07
r37 19 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.415 $Y=2.5
+ $X2=0.415 $Y2=3.07
r38 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=2.5 $X2=0.415 $Y2=2.5
r39 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.5
+ $X2=0.415 $Y2=2.665
r40 15 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.5
+ $X2=0.415 $Y2=2.335
r41 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=0.355 $Y=1.515
+ $X2=0.475 $Y2=1.515
r42 8 17 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.665
r43 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=1.515
r44 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=0.945
r45 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.355 $Y=1.59
+ $X2=0.355 $Y2=1.515
r46 1 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.355 $Y=1.59
+ $X2=0.355 $Y2=2.335
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%A1 3 7 10 15 18 22
c52 22 0 1.46798e-19 $X=0.895 $Y=2.7
c53 15 0 8.80277e-21 $X=0.815 $Y=1.96
r54 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.895 $Y=2.7
+ $X2=0.895 $Y2=2.7
r55 18 19 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=2.7
+ $X2=0.855 $Y2=2.615
r56 15 19 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.815 $Y=1.96
+ $X2=0.815 $Y2=2.615
r57 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=1.96 $X2=0.815 $Y2=1.96
r58 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.815 $Y=1.96
+ $X2=0.815 $Y2=2.095
r59 10 11 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.815 $Y=1.96
+ $X2=0.815 $Y2=1.825
r60 7 11 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=1.825
r61 3 12 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=0.835 $Y=3.825
+ $X2=0.835 $Y2=2.095
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%B0 3 7 10 15 20 23
c49 15 0 1.46798e-19 $X=1.2 $Y=2.33
c50 10 0 8.80277e-21 $X=1.325 $Y=1.64
r51 17 20 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.64
+ $X2=1.325 $Y2=1.64
r52 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.33 $X2=1.2
+ $Y2=2.33
r53 13 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=1.805 $X2=1.2
+ $Y2=1.64
r54 13 15 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.2 $Y=1.805
+ $X2=1.2 $Y2=2.33
r55 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.64 $X2=1.325 $Y2=1.64
r56 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.64
+ $X2=1.325 $Y2=1.805
r57 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.64
+ $X2=1.325 $Y2=1.475
r58 7 12 1035.79 $w=1.5e-07 $l=2.02e-06 $layer=POLY_cond $X=1.335 $Y=3.825
+ $X2=1.335 $Y2=1.805
r59 3 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=0.945
+ $X2=1.335 $Y2=1.475
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%B1 3 6 10 11 15 18 23
r31 18 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.005 $Y=1.965
+ $X2=2.005 $Y2=1.965
r32 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=1.965 $X2=2.005 $Y2=1.965
r33 12 15 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.765 $Y=1.965
+ $X2=2.005 $Y2=1.965
r34 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.73 $Y=2.55
+ $X2=1.73 $Y2=2.7
r35 8 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.13
+ $X2=1.765 $Y2=1.965
r36 8 10 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.765 $Y=2.13
+ $X2=1.765 $Y2=2.55
r37 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.8
+ $X2=1.765 $Y2=1.965
r38 4 6 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.765 $Y=1.8
+ $X2=1.765 $Y2=0.945
r39 3 11 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.695 $Y=3.825
+ $X2=1.695 $Y2=2.7
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%Y 1 3 11 15 16 19 23 28 31 33 36
r46 31 36 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.665 $Y=1.475
+ $X2=1.665 $Y2=1.59
r47 30 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.665 $Y=1.335
+ $X2=1.665 $Y2=1.22
r48 30 31 0.134804 $w=1.7e-07 $l=1.4e-07 $layer=MET1_cond $X=1.665 $Y=1.335
+ $X2=1.665 $Y2=1.475
r49 28 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.665 $Y=1.22
+ $X2=1.665 $Y2=1.22
r50 25 28 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=1.22
+ $X2=1.665 $Y2=1.22
r51 23 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.665 $Y=1.59
+ $X2=1.665 $Y2=1.59
r52 21 23 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=1.665 $Y=3.07
+ $X2=1.665 $Y2=1.59
r53 17 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.135
+ $X2=1.55 $Y2=1.22
r54 17 19 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.55 $Y=1.135
+ $X2=1.55 $Y2=0.99
r55 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=3.155
+ $X2=1.665 $Y2=3.07
r56 15 16 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.58 $Y=3.155
+ $X2=1.17 $Y2=3.155
r57 11 13 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.085 $Y=3.545
+ $X2=1.085 $Y2=4.565
r58 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.085 $Y=3.24
+ $X2=1.17 $Y2=3.155
r59 9 11 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.085 $Y=3.24
+ $X2=1.085 $Y2=3.545
r60 3 13 300 $w=1.7e-07 $l=1.8254e-06 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.825 $X2=1.085 $Y2=4.565
r61 3 11 300 $w=1.7e-07 $l=8.02745e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.825 $X2=1.085 $Y2=3.545
r62 1 19 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.99
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OAI22_L%A_27_115# 1 2 3 15 17 18 23 24 25
r28 25 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.98 $Y=0.56
+ $X2=1.98 $Y2=0.74
r29 23 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.56
+ $X2=1.98 $Y2=0.56
r30 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=0.56
+ $X2=1.205 $Y2=0.56
r31 20 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.12 $Y=1.075
+ $X2=1.12 $Y2=0.865
r32 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.645
+ $X2=1.205 $Y2=0.56
r33 19 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.12 $Y=0.645
+ $X2=1.12 $Y2=0.865
r34 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=1.12 $Y2=1.075
r35 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.345 $Y2=1.16
r36 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.345 $Y2=1.16
r37 13 15 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.26 $Y2=0.865
r38 3 28 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.74
r39 2 22 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r40 1 15 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

