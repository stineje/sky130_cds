* File: sky130_osu_sc_15T_ms__tbufi_l.spice
* Created: Fri Nov 12 14:46:42 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__tbufi_l.pex.spice"
.subckt sky130_osu_sc_15T_ms__tbufi_l  GND VDD OE A Y
* 
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_OE_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1000 A_196_115# N_OE_M1000_g N_GND_M1002_d N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.5 A=0.078 P=1.34 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_196_115# N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0546 PD=1.57 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75001
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1001 N_VDD_M1001_d N_OE_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001 A=0.189 P=2.82 MULT=1
MM1005 A_196_713# N_A_27_115#_M1005_g N_VDD_M1001_d N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g A_196_713# N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=5.664 P=9.74
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__tbufi_l.pxi.spice"
*
.ends
*
*
