* File: sky130_osu_sc_15T_ls__inv_l.pex.spice
* Created: Fri Nov 12 14:58:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__INV_L%GND 1 11 15 24 27
r14 24 27 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=0.19
+ $X2=0.495 $Y2=0.24
r15 13 15 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r16 11 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r17 11 13 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r18 1 15 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__INV_L%VDD 1 9 13 18 21
r10 21 24 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=5.31
+ $X2=0.495 $Y2=5.36
r11 18 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r12 11 18 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r13 11 13 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r14 9 18 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r15 1 13 600 $w=1.7e-07 $l=1.06066e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.565
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__INV_L%A 3 7 10 15 17 19 22
r34 17 19 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.045
+ $X2=0.535 $Y2=2.045
r35 15 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r36 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.405 $Y2=2.045
r37 13 15 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.32 $Y2=3.07
r38 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.045 $X2=0.535 $Y2=2.045
r39 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=2.21
r40 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=1.88
r41 7 12 1017.84 $w=1.5e-07 $l=1.985e-06 $layer=POLY_cond $X=0.475 $Y=4.195
+ $X2=0.475 $Y2=2.21
r42 3 11 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.88
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__INV_L%Y 1 3 10 16 24 27 30
r30 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=2.7
r31 22 24 0.616245 $w=1.7e-07 $l=6.4e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=1.945
r32 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.22
r33 21 24 0.587358 $w=1.7e-07 $l=6.1e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.945
r34 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.7 $X2=0.69
+ $Y2=2.7
r35 16 19 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=4.565
r36 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.22
+ $X2=0.69 $Y2=1.22
r37 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.69 $Y=0.74
+ $X2=0.69 $Y2=1.22
r38 3 19 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.565 $X2=0.69 $Y2=4.565
r39 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

