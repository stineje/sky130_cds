* File: sky130_osu_sc_12T_ls__inv_3.pex.spice
* Created: Fri Nov 12 15:37:48 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__INV_3%GND 1 2 21 25 27 35 42 44 47
r49 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r50 33 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r51 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r52 27 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r53 23 25 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r54 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r55 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r56 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r57 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r58 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r59 2 35 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
r60 1 25 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_3%VDD 1 2 17 21 23 30 38 40 43
r33 40 43 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r34 30 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r35 28 38 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r36 28 33 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135 $X2=1.12
+ $Y2=3.635
r37 26 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r38 24 37 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r39 24 26 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r40 23 38 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r41 23 26 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r42 19 37 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r43 19 21 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135 $X2=0.26
+ $Y2=3.635
r44 17 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r45 17 37 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r46 2 33 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r47 2 30 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r48 1 21 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_3%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 34 36 37 38 41 43 45 48
c96 33 0 1.50926e-19 $X=0.535 $Y=1.825
c97 28 0 1.33323e-19 $X=1.335 $Y=2.48
c98 25 0 1.33323e-19 $X=1.335 $Y=1.22
c99 18 0 1.33323e-19 $X=0.905 $Y=2.48
c100 15 0 1.33323e-19 $X=0.905 $Y=1.22
r101 48 51 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=2.845
+ $X2=0.405 $Y2=2.85
r102 43 45 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=1.825
+ $X2=0.535 $Y2=1.825
r103 41 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r104 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.405 $Y2=1.825
r105 39 41 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.32 $Y2=2.85
r106 33 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.825 $X2=0.535 $Y2=1.825
r107 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.99
r108 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.66
r109 28 30 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r110 25 27 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=0.835
r111 24 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.405
+ $X2=0.905 $Y2=2.405
r112 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=1.335 $Y2=2.48
r113 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=0.98 $Y2=2.405
r114 22 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.295
+ $X2=0.905 $Y2=1.295
r115 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=1.335 $Y2=1.22
r116 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=0.98 $Y2=1.295
r117 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=2.405
r118 18 20 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=3.235
r119 15 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=1.295
r120 15 17 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=0.835
r121 14 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.405
+ $X2=0.475 $Y2=2.405
r122 13 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.905 $Y2=2.405
r123 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.55 $Y2=2.405
r124 12 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.475 $Y2=1.295
r125 11 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.905 $Y2=1.295
r126 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.55 $Y2=1.295
r127 8 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=2.405
r128 8 10 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=3.235
r129 7 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=2.405
r130 7 35 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=1.99
r131 4 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.295
r132 4 34 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.66
r133 1 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=1.295
r134 1 3 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_3%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c78 55 0 1.33323e-19 $X=1.55 $Y=2.365
c79 54 0 1.33323e-19 $X=1.55 $Y=1.115
c80 46 0 1.33323e-19 $X=0.69 $Y=2.365
c81 45 0 1.33323e-19 $X=0.69 $Y=1.115
c82 18 0 1.50926e-19 $X=0.69 $Y=0.755
r83 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.48
r84 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r85 54 55 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=2.365
r86 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.48
+ $X2=0.69 $Y2=2.48
r87 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=1.55 $Y2=2.48
r88 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=0.835 $Y2=2.48
r89 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1
+ $X2=0.69 $Y2=1
r90 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=1.55 $Y2=1
r91 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=0.835 $Y2=1
r92 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.48
r93 46 48 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=1.72
r94 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1
r95 45 48 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1.72
r96 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r97 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.48
r98 38 41 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.955
r99 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r100 32 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r101 27 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r102 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r103 24 27 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.955
r104 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1 $X2=0.69
+ $Y2=1
r105 18 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0.755
+ $X2=0.69 $Y2=1
r106 6 43 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r107 6 41 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r108 5 29 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r109 5 27 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r110 2 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
r111 1 18 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

