* File: sky130_osu_sc_18T_ms__tbufi_l.pex.spice
* Created: Thu Oct 29 17:31:39 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%GND 1 12 14 21 26 29
r35 26 29 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r36 23 24 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r37 19 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r38 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r39 14 24 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r40 12 23 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r41 12 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r42 12 14 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r43 1 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%VDD 1 10 12 18 25 28 32
r21 28 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r22 25 28 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r23 22 32 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507 $X2=1.02
+ $Y2=6.507
r24 22 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r25 18 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=4.475
+ $X2=0.69 $Y2=5.835
r26 16 23 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r27 16 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r28 12 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r29 12 14 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r30 10 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r31 10 14 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r32 1 21 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=5.835
r33 1 18 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%OE 2 5 9 13 17 22 23 26 32
c62 22 0 2.60266e-19 $X=0.69 $Y=1.85
r63 23 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.85 $X2=0.69 $Y2=1.85
r64 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=1.85
r65 19 22 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.965
+ $X2=0.69 $Y2=1.85
r66 19 26 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=0.69 $Y=1.965
+ $X2=0.69 $Y2=2.845
r67 15 17 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.935
+ $X2=0.475 $Y2=2.935
r68 11 32 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.905 $Y=1.65
+ $X2=0.69 $Y2=1.832
r69 11 13 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=1.65
+ $X2=0.905 $Y2=0.945
r70 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.475 $Y2=2.935
r71 7 9 1063.99 $w=1.5e-07 $l=2.075e-06 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.475 $Y2=5.085
r72 3 32 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.69 $Y2=1.832
r73 3 5 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=1.65 $X2=0.475
+ $Y2=0.945
r74 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.86 $X2=0.27
+ $Y2=2.935
r75 1 3 44.3094 $w=2.23e-07 $l=2.69768e-07 $layer=POLY_cond $X=0.27 $Y=1.8
+ $X2=0.475 $Y2=1.65
r76 1 2 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.8 $X2=0.27
+ $Y2=2.86
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%A_27_115# 1 2 9 13 17 21 23 26 31
r50 27 31 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.8 $Y=2.48
+ $X2=0.905 $Y2=2.48
r51 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=2.48 $X2=0.8 $Y2=2.48
r52 22 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.48
+ $X2=0.26 $Y2=2.48
r53 21 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.48
+ $X2=0.8 $Y2=2.48
r54 21 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=2.48
+ $X2=0.345 $Y2=2.48
r55 17 19 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=4.475
+ $X2=0.26 $Y2=5.835
r56 15 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.565
+ $X2=0.26 $Y2=2.48
r57 15 17 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=0.26 $Y=2.565
+ $X2=0.26 $Y2=4.475
r58 11 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.395
+ $X2=0.26 $Y2=2.48
r59 11 13 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=0.26 $Y=2.395
+ $X2=0.26 $Y2=0.825
r60 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.645
+ $X2=0.905 $Y2=2.48
r61 7 9 1251.15 $w=1.5e-07 $l=2.44e-06 $layer=POLY_cond $X=0.905 $Y=2.645
+ $X2=0.905 $Y2=5.085
r62 2 19 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=5.835
r63 2 17 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=4.475
r64 1 13 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%A 3 7 13 14 17 19
c46 14 0 1.90743e-19 $X=1.325 $Y=2.09
c47 3 0 6.95226e-20 $X=1.265 $Y=0.945
r48 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=3.33
+ $X2=1.14 $Y2=3.33
r49 14 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.09
+ $X2=1.325 $Y2=2.255
r50 14 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.09
+ $X2=1.325 $Y2=1.925
r51 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.09 $X2=1.325 $Y2=2.09
r52 10 19 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=2.175
+ $X2=1.14 $Y2=3.33
r53 9 13 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=2.09
+ $X2=1.325 $Y2=2.09
r54 9 10 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.09 $X2=1.14
+ $Y2=2.175
r55 7 23 1451.13 $w=1.5e-07 $l=2.83e-06 $layer=POLY_cond $X=1.265 $Y=5.085
+ $X2=1.265 $Y2=2.255
r56 3 22 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.265 $Y=0.945
+ $X2=1.265 $Y2=1.925
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%Y 1 2 10 13 17 18 21
r34 28 30 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.48 $Y=4.475
+ $X2=1.48 $Y2=5.835
r35 18 28 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=1.48 $Y=2.59
+ $X2=1.48 $Y2=4.475
r36 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.59
+ $X2=1.48 $Y2=2.59
r37 14 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.48 $Y=1.48
+ $X2=1.48 $Y2=0.825
r38 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.48
+ $X2=1.48 $Y2=1.48
r39 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.475
+ $X2=1.48 $Y2=2.59
r40 8 10 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.475
+ $X2=1.48 $Y2=1.82
r41 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.595
+ $X2=1.48 $Y2=1.48
r42 7 10 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.595
+ $X2=1.48 $Y2=1.82
r43 2 30 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=4.085 $X2=1.48 $Y2=5.835
r44 2 28 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=4.085 $X2=1.48 $Y2=4.475
r45 1 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.825
.ends

