* File: sky130_osu_sc_12T_ms__dlat_1.spice
* Created: Fri Nov 12 15:23:29 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ms__dlat_1.pex.spice"
.subckt sky130_osu_sc_12T_ms__dlat_1  GND VDD D CK ON Q
* 
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1002 A_115_115# N_D_M1002_g N_GND_M1002_s N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1015 N_D_M1015_d N_CK_M1015_g A_115_115# N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1013 A_307_115# N_A_157_349#_M1013_g N_D_M1015_d N_GND_M1002_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.1 SB=75001 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_A_349_89#_M1007_g A_307_115# N_GND_M1002_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.5 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1008 N_A_157_349#_M1008_d N_CK_M1008_g N_GND_M1007_d N_GND_M1002_b NSHORT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.9 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1009 N_A_349_89#_M1009_d N_D_M1009_g N_GND_M1009_s N_GND_M1002_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.1378 PD=1.57 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1011 N_GND_M1011_d N_A_349_89#_M1011_g N_ON_M1011_s N_GND_M1002_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1012 N_Q_M1012_d N_ON_M1012_g N_GND_M1011_d N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1014 A_115_521# N_D_M1014_g N_VDD_M1014_s N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1010 N_D_M1010_d N_A_157_349#_M1010_g A_115_521# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1006 A_307_521# N_CK_M1006_g N_D_M1010_d N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.1 SB=75001 A=0.189 P=2.82 MULT=1
MM1000 N_VDD_M1000_d N_A_349_89#_M1000_g A_307_521# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_157_349#_M1001_d N_CK_M1001_g N_VDD_M1000_d N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_349_89#_M1003_d N_D_M1003_g N_VDD_M1003_s N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_349_89#_M1004_g N_ON_M1004_s N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Q_M1005_d N_ON_M1005_g N_VDD_M1004_d N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref N_GND_M1002_b N_VDD_M1014_b NWDIODE A=10.5987 P=14.41
pX17_noxref noxref_13 D D PROBETYPE=1
pX18_noxref noxref_14 CK CK PROBETYPE=1
pX19_noxref noxref_15 ON ON PROBETYPE=1
pX20_noxref noxref_16 Q Q PROBETYPE=1
c_836 A_115_521# 0 1.57671e-19 $X=0.575 $Y=2.605
*
.include "sky130_osu_sc_12T_ms__dlat_1.pxi.spice"
*
.ends
*
*
