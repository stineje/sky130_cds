* File: sky130_osu_sc_15T_ms__or2_2.pxi.spice
* Created: Fri Nov 12 14:46:00 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__OR2_2%GND N_GND_M1005_s N_GND_M1001_d N_GND_M1007_s
+ N_GND_M1005_b N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p N_GND_c_24_p
+ GND N_GND_c_4_p PM_SKY130_OSU_SC_15T_MS__OR2_2%GND
x_PM_SKY130_OSU_SC_15T_MS__OR2_2%VDD N_VDD_M1003_d N_VDD_M1004_d N_VDD_M1006_b
+ N_VDD_c_45_p N_VDD_c_51_p N_VDD_c_58_p N_VDD_c_64_p VDD N_VDD_c_46_p
+ PM_SKY130_OSU_SC_15T_MS__OR2_2%VDD
x_PM_SKY130_OSU_SC_15T_MS__OR2_2%B N_B_M1005_g N_B_M1006_g N_B_c_79_n N_B_c_80_n
+ B PM_SKY130_OSU_SC_15T_MS__OR2_2%B
x_PM_SKY130_OSU_SC_15T_MS__OR2_2%A N_A_M1001_g N_A_M1003_g N_A_c_107_n
+ N_A_c_108_n A PM_SKY130_OSU_SC_15T_MS__OR2_2%A
x_PM_SKY130_OSU_SC_15T_MS__OR2_2%A_27_565# N_A_27_565#_M1005_d
+ N_A_27_565#_M1006_s N_A_27_565#_M1002_g N_A_27_565#_c_165_n
+ N_A_27_565#_M1000_g N_A_27_565#_c_150_n N_A_27_565#_c_151_n
+ N_A_27_565#_M1007_g N_A_27_565#_c_170_n N_A_27_565#_M1004_g
+ N_A_27_565#_c_156_n N_A_27_565#_c_157_n N_A_27_565#_c_176_n
+ N_A_27_565#_c_180_n N_A_27_565#_c_182_n N_A_27_565#_c_158_n
+ N_A_27_565#_c_159_n N_A_27_565#_c_162_n N_A_27_565#_c_164_n
+ PM_SKY130_OSU_SC_15T_MS__OR2_2%A_27_565#
x_PM_SKY130_OSU_SC_15T_MS__OR2_2%Y N_Y_M1002_d N_Y_M1000_s N_Y_c_236_n
+ N_Y_c_239_n Y N_Y_c_241_n N_Y_c_244_n PM_SKY130_OSU_SC_15T_MS__OR2_2%Y
cc_1 N_GND_M1005_b N_B_M1005_g 0.083817f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_B_M1005_g 0.00866533f $X=0.26 $Y=0.865 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_B_M1005_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.945
cc_4 N_GND_c_4_p N_B_M1005_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=0.945
cc_5 N_GND_M1005_b N_B_M1006_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_6 N_GND_M1005_b N_B_c_79_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.415
cc_7 N_GND_M1005_b N_B_c_80_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.415
cc_8 N_GND_M1005_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.7
cc_9 N_GND_M1005_b N_A_M1001_g 0.0440597f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.945
cc_10 N_GND_c_3_p N_A_M1001_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.945
cc_11 N_GND_c_11_p N_A_M1001_g 0.00388248f $X=1.12 $Y=0.865 $X2=0.905 $Y2=0.945
cc_12 N_GND_c_4_p N_A_M1001_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.905 $Y2=0.945
cc_13 N_GND_M1005_b N_A_M1003_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_14 N_GND_M1005_b N_A_c_107_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.125
cc_15 N_GND_M1005_b N_A_c_108_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.125
cc_16 N_GND_M1005_b N_A_27_565#_M1002_g 0.0207501f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.945
cc_17 N_GND_c_11_p N_A_27_565#_M1002_g 0.00388248f $X=1.12 $Y=0.865 $X2=1.335
+ $Y2=0.945
cc_18 N_GND_c_18_p N_A_27_565#_M1002_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.945
cc_19 N_GND_c_4_p N_A_27_565#_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335
+ $Y2=0.945
cc_20 N_GND_M1005_b N_A_27_565#_c_150_n 0.0466273f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.55
cc_21 N_GND_M1005_b N_A_27_565#_c_151_n 0.0244031f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.625
cc_22 N_GND_M1005_b N_A_27_565#_M1007_g 0.0264941f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.945
cc_23 N_GND_c_18_p N_A_27_565#_M1007_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.945
cc_24 N_GND_c_24_p N_A_27_565#_M1007_g 0.00866533f $X=1.98 $Y=0.865 $X2=1.765
+ $Y2=0.945
cc_25 N_GND_c_4_p N_A_27_565#_M1007_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765
+ $Y2=0.945
cc_26 N_GND_M1005_b N_A_27_565#_c_156_n 0.00567173f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.625
cc_27 N_GND_M1005_b N_A_27_565#_c_157_n 0.0539419f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_28 N_GND_M1005_b N_A_27_565#_c_158_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.285
cc_29 N_GND_M1005_b N_A_27_565#_c_159_n 0.00710171f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.865
cc_30 N_GND_c_3_p N_A_27_565#_c_159_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.865
cc_31 N_GND_c_4_p N_A_27_565#_c_159_n 0.00475776f $X=1.7 $Y=0.19 $X2=0.69
+ $Y2=0.865
cc_32 N_GND_M1005_b N_A_27_565#_c_162_n 0.0190355f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_33 N_GND_c_11_p N_A_27_565#_c_162_n 0.00702738f $X=1.12 $Y=0.865 $X2=1.43
+ $Y2=1.675
cc_34 N_GND_M1005_b N_A_27_565#_c_164_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.675
cc_35 N_GND_M1005_b N_Y_c_236_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.865
cc_36 N_GND_c_18_p N_Y_c_236_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.865
cc_37 N_GND_c_4_p N_Y_c_236_n 0.00475776f $X=1.7 $Y=0.19 $X2=1.55 $Y2=0.865
cc_38 N_GND_M1005_b N_Y_c_239_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_39 N_GND_M1005_b Y 0.0306725f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.96
cc_40 N_GND_M1005_b N_Y_c_241_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.22
cc_41 N_GND_c_11_p N_Y_c_241_n 0.00125659f $X=1.12 $Y=0.865 $X2=1.55 $Y2=1.22
cc_42 N_GND_c_24_p N_Y_c_241_n 0.00125659f $X=1.98 $Y=0.865 $X2=1.55 $Y2=1.22
cc_43 N_GND_M1005_b N_Y_c_244_n 0.0111067f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_44 N_VDD_M1006_b N_B_M1006_g 0.0264002f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_45 N_VDD_c_45_p N_B_M1006_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475 $Y2=3.825
cc_46 N_VDD_c_46_p N_B_M1006_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.475 $Y2=3.825
cc_47 N_VDD_M1006_b N_B_c_80_n 0.00375034f $X=-0.045 $Y=2.645 $X2=0.27 $Y2=2.415
cc_48 N_VDD_M1006_b B 0.0108395f $X=-0.045 $Y=2.645 $X2=0.27 $Y2=2.7
cc_49 N_VDD_M1006_b N_A_M1003_g 0.0199048f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_50 N_VDD_c_45_p N_A_M1003_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905 $Y2=3.825
cc_51 N_VDD_c_51_p N_A_M1003_g 0.00362996f $X=1.12 $Y=3.885 $X2=0.905 $Y2=3.825
cc_52 N_VDD_c_46_p N_A_M1003_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.905 $Y2=3.825
cc_53 N_VDD_M1006_b N_A_c_108_n 0.00153494f $X=-0.045 $Y=2.645 $X2=0.95
+ $Y2=2.125
cc_54 N_VDD_M1003_d A 0.0077995f $X=0.98 $Y=2.825 $X2=0.95 $Y2=3.07
cc_55 N_VDD_c_51_p A 0.00247404f $X=1.12 $Y=3.885 $X2=0.95 $Y2=3.07
cc_56 N_VDD_M1006_b N_A_27_565#_c_165_n 0.0174876f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.7
cc_57 N_VDD_c_51_p N_A_27_565#_c_165_n 0.00362996f $X=1.12 $Y=3.885 $X2=1.335
+ $Y2=2.7
cc_58 N_VDD_c_58_p N_A_27_565#_c_165_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335
+ $Y2=2.7
cc_59 N_VDD_c_46_p N_A_27_565#_c_165_n 0.00429146f $X=1.7 $Y=5.36 $X2=1.335
+ $Y2=2.7
cc_60 N_VDD_M1006_b N_A_27_565#_c_151_n 0.00813142f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_61 N_VDD_M1006_b N_A_27_565#_c_170_n 0.0216047f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.7
cc_62 N_VDD_c_51_p N_A_27_565#_c_170_n 3.67508e-19 $X=1.12 $Y=3.885 $X2=1.765
+ $Y2=2.7
cc_63 N_VDD_c_58_p N_A_27_565#_c_170_n 0.00500229f $X=1.895 $Y=5.397 $X2=1.765
+ $Y2=2.7
cc_64 N_VDD_c_64_p N_A_27_565#_c_170_n 0.00771008f $X=1.98 $Y=3.205 $X2=1.765
+ $Y2=2.7
cc_65 N_VDD_c_46_p N_A_27_565#_c_170_n 0.00430409f $X=1.7 $Y=5.36 $X2=1.765
+ $Y2=2.7
cc_66 N_VDD_M1006_b N_A_27_565#_c_156_n 0.00216365f $X=-0.045 $Y=2.645 $X2=1.352
+ $Y2=2.625
cc_67 N_VDD_M1006_b N_A_27_565#_c_176_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.545
cc_68 N_VDD_c_45_p N_A_27_565#_c_176_n 0.00452684f $X=1.035 $Y=5.397 $X2=0.26
+ $Y2=3.545
cc_69 N_VDD_c_46_p N_A_27_565#_c_176_n 0.00435496f $X=1.7 $Y=5.36 $X2=0.26
+ $Y2=3.545
cc_70 N_VDD_M1006_b N_A_27_565#_c_158_n 0.00106577f $X=-0.045 $Y=2.645 $X2=0.61
+ $Y2=3.285
cc_71 N_VDD_M1006_b N_Y_c_239_n 0.00410619f $X=-0.045 $Y=2.645 $X2=1.55 $Y2=2.33
cc_72 N_VDD_c_58_p N_Y_c_239_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.33
cc_73 N_VDD_c_46_p N_Y_c_239_n 0.00434939f $X=1.7 $Y=5.36 $X2=1.55 $Y2=2.33
cc_74 N_B_M1005_g N_A_M1001_g 0.0430073f $X=0.475 $Y=0.945 $X2=0.905 $Y2=0.945
cc_75 N_B_c_79_n N_A_M1003_g 0.112923f $X=0.475 $Y=2.415 $X2=0.905 $Y2=3.825
cc_76 N_B_M1005_g N_A_c_107_n 0.0148656f $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.125
cc_77 N_B_M1005_g N_A_c_108_n 0.00121111f $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.125
cc_78 N_B_M1006_g N_A_27_565#_c_180_n 0.0142177f $X=0.475 $Y=3.825 $X2=0.525
+ $Y2=3.37
cc_79 B N_A_27_565#_c_180_n 0.00520961f $X=0.27 $Y=2.7 $X2=0.525 $Y2=3.37
cc_80 N_B_c_80_n N_A_27_565#_c_182_n 0.00369517f $X=0.27 $Y=2.415 $X2=0.345
+ $Y2=3.37
cc_81 B N_A_27_565#_c_182_n 0.00431991f $X=0.27 $Y=2.7 $X2=0.345 $Y2=3.37
cc_82 N_B_M1005_g N_A_27_565#_c_158_n 0.0231435f $X=0.475 $Y=0.945 $X2=0.61
+ $Y2=3.285
cc_83 N_B_M1006_g N_A_27_565#_c_158_n 0.026563f $X=0.475 $Y=3.825 $X2=0.61
+ $Y2=3.285
cc_84 N_B_c_79_n N_A_27_565#_c_158_n 0.00764878f $X=0.475 $Y=2.415 $X2=0.61
+ $Y2=3.285
cc_85 N_B_c_80_n N_A_27_565#_c_158_n 0.0350086f $X=0.27 $Y=2.415 $X2=0.61
+ $Y2=3.285
cc_86 B N_A_27_565#_c_158_n 0.00758489f $X=0.27 $Y=2.7 $X2=0.61 $Y2=3.285
cc_87 N_B_M1005_g N_A_27_565#_c_159_n 0.00799668f $X=0.475 $Y=0.945 $X2=0.69
+ $Y2=0.865
cc_88 N_B_M1005_g N_A_27_565#_c_164_n 0.0113001f $X=0.475 $Y=0.945 $X2=0.65
+ $Y2=1.675
cc_89 N_A_M1001_g N_A_27_565#_M1002_g 0.033724f $X=0.905 $Y=0.945 $X2=1.335
+ $Y2=0.945
cc_90 A N_A_27_565#_c_165_n 0.00374181f $X=0.95 $Y=3.07 $X2=1.335 $Y2=2.7
cc_91 N_A_M1003_g N_A_27_565#_c_150_n 0.00914307f $X=0.905 $Y=3.825 $X2=1.37
+ $Y2=2.55
cc_92 N_A_c_107_n N_A_27_565#_c_150_n 0.0204279f $X=0.95 $Y=2.125 $X2=1.37
+ $Y2=2.55
cc_93 N_A_c_108_n N_A_27_565#_c_150_n 0.00375034f $X=0.95 $Y=2.125 $X2=1.37
+ $Y2=2.55
cc_94 N_A_M1003_g N_A_27_565#_c_156_n 0.0553014f $X=0.905 $Y=3.825 $X2=1.352
+ $Y2=2.625
cc_95 N_A_c_108_n N_A_27_565#_c_156_n 0.00355256f $X=0.95 $Y=2.125 $X2=1.352
+ $Y2=2.625
cc_96 N_A_M1001_g N_A_27_565#_c_157_n 0.0119161f $X=0.905 $Y=0.945 $X2=1.43
+ $Y2=1.675
cc_97 N_A_M1003_g N_A_27_565#_c_180_n 0.00457566f $X=0.905 $Y=3.825 $X2=0.525
+ $Y2=3.37
cc_98 N_A_M1001_g N_A_27_565#_c_158_n 0.00429604f $X=0.905 $Y=0.945 $X2=0.61
+ $Y2=3.285
cc_99 N_A_M1003_g N_A_27_565#_c_158_n 0.00776428f $X=0.905 $Y=3.825 $X2=0.61
+ $Y2=3.285
cc_100 N_A_c_107_n N_A_27_565#_c_158_n 0.0021255f $X=0.95 $Y=2.125 $X2=0.61
+ $Y2=3.285
cc_101 N_A_c_108_n N_A_27_565#_c_158_n 0.0822139f $X=0.95 $Y=2.125 $X2=0.61
+ $Y2=3.285
cc_102 A N_A_27_565#_c_158_n 0.00866797f $X=0.95 $Y=3.07 $X2=0.61 $Y2=3.285
cc_103 N_A_M1001_g N_A_27_565#_c_159_n 0.00799668f $X=0.905 $Y=0.945 $X2=0.69
+ $Y2=0.865
cc_104 N_A_M1001_g N_A_27_565#_c_162_n 0.0163305f $X=0.905 $Y=0.945 $X2=1.43
+ $Y2=1.675
cc_105 N_A_c_107_n N_A_27_565#_c_162_n 0.00276813f $X=0.95 $Y=2.125 $X2=1.43
+ $Y2=1.675
cc_106 N_A_c_108_n N_A_27_565#_c_162_n 0.0114342f $X=0.95 $Y=2.125 $X2=1.43
+ $Y2=1.675
cc_107 A A_110_565# 0.0123256f $X=0.95 $Y=3.07 $X2=0.55 $Y2=2.825
cc_108 N_A_c_108_n N_Y_c_239_n 0.0206732f $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.33
cc_109 A N_Y_c_239_n 0.00659455f $X=0.95 $Y=3.07 $X2=1.55 $Y2=2.33
cc_110 N_A_M1001_g Y 6.73508e-19 $X=0.905 $Y=0.945 $X2=1.555 $Y2=1.96
cc_111 N_A_c_108_n Y 0.00825539f $X=0.95 $Y=2.125 $X2=1.555 $Y2=1.96
cc_112 N_A_M1001_g N_Y_c_241_n 7.99941e-19 $X=0.905 $Y=0.945 $X2=1.55 $Y2=1.22
cc_113 N_A_c_107_n N_Y_c_244_n 3.65268e-19 $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.33
cc_114 N_A_c_108_n N_Y_c_244_n 0.00535705f $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.33
cc_115 N_A_27_565#_c_180_n A_110_565# 0.00613297f $X=0.525 $Y=3.37 $X2=0.55
+ $Y2=2.825
cc_116 N_A_27_565#_c_158_n A_110_565# 0.00377193f $X=0.61 $Y=3.285 $X2=0.55
+ $Y2=2.825
cc_117 N_A_27_565#_M1002_g N_Y_c_236_n 0.00265306f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=0.865
cc_118 N_A_27_565#_M1007_g N_Y_c_236_n 0.00265306f $X=1.765 $Y=0.945 $X2=1.55
+ $Y2=0.865
cc_119 N_A_27_565#_c_157_n N_Y_c_236_n 0.00171364f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.865
cc_120 N_A_27_565#_c_162_n N_Y_c_236_n 0.00500271f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.865
cc_121 N_A_27_565#_c_165_n N_Y_c_239_n 0.00234922f $X=1.335 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_122 N_A_27_565#_c_150_n N_Y_c_239_n 0.00744772f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_123 N_A_27_565#_c_151_n N_Y_c_239_n 0.0160452f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_124 N_A_27_565#_c_170_n N_Y_c_239_n 0.00401146f $X=1.765 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_125 N_A_27_565#_c_157_n N_Y_c_239_n 0.0013767f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_126 N_A_27_565#_c_162_n N_Y_c_239_n 0.00273485f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_127 N_A_27_565#_M1002_g Y 0.00251111f $X=1.335 $Y=0.945 $X2=1.555 $Y2=1.96
cc_128 N_A_27_565#_c_150_n Y 0.00892438f $X=1.37 $Y=2.55 $X2=1.555 $Y2=1.96
cc_129 N_A_27_565#_M1007_g Y 0.00251111f $X=1.765 $Y=0.945 $X2=1.555 $Y2=1.96
cc_130 N_A_27_565#_c_157_n Y 0.0120226f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_131 N_A_27_565#_c_162_n Y 0.0147088f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_132 N_A_27_565#_M1002_g N_Y_c_241_n 0.00527857f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=1.22
cc_133 N_A_27_565#_M1007_g N_Y_c_241_n 0.00908199f $X=1.765 $Y=0.945 $X2=1.55
+ $Y2=1.22
cc_134 N_A_27_565#_c_162_n N_Y_c_241_n 0.00238892f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=1.22
cc_135 N_A_27_565#_c_150_n N_Y_c_244_n 0.00740115f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_136 N_A_27_565#_c_151_n N_Y_c_244_n 0.00229755f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_137 N_A_27_565#_c_157_n N_Y_c_244_n 0.00174847f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_138 N_A_27_565#_c_162_n N_Y_c_244_n 0.00181779f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
