* File: sky130_osu_sc_15T_ms__aoi21_l.pex.spice
* Created: Fri Nov 12 14:41:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%GND 1 2 21 25 27 35 41 44
c41 21 0 6.36774e-20 $X=-0.045 $Y=0
r42 41 44 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r43 33 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.54 $Y=0.305
+ $X2=1.54 $Y2=0.74
r44 27 33 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.455 $Y=0.152
+ $X2=1.54 $Y2=0.305
r45 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r46 21 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r47 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r48 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r49 21 27 16.4365 $w=3.03e-07 $l=4.35e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.455 $Y2=0.152
r50 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r51 2 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.74
r52 1 25 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%VDD 1 13 15 21 25 29 32
r26 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r27 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r28 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r29 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397 $X2=1.02
+ $Y2=5.397
r30 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r31 19 21 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.235
r32 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r33 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r34 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r35 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r36 1 21 300 $w=1.7e-07 $l=1.47834e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.235
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%A0 2 3 5 8 12 18 21 27
c37 8 0 6.36774e-20 $X=0.475 $Y=3.825
r38 24 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=3.07
+ $X2=0.385 $Y2=3.07
r39 21 24 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.385 $Y=2.505
+ $X2=0.385 $Y2=3.07
r40 17 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.505 $X2=0.385 $Y2=2.505
r41 17 18 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.505
+ $X2=0.475 $Y2=2.505
r42 14 17 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.505
+ $X2=0.385 $Y2=2.505
r43 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.51
+ $X2=0.475 $Y2=1.51
r44 6 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.64
+ $X2=0.475 $Y2=2.505
r45 6 8 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.475 $Y=2.64
+ $X2=0.475 $Y2=3.825
r46 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.43 $X2=0.475
+ $Y2=1.51
r47 3 5 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.475 $Y=1.43
+ $X2=0.475 $Y2=0.945
r48 2 14 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.37
+ $X2=0.295 $Y2=2.505
r49 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.59 $X2=0.295
+ $Y2=1.51
r50 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.59
+ $X2=0.295 $Y2=2.37
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%A1 3 7 10 15 20 23
c50 23 0 1.38614e-19 $X=0.725 $Y=2.7
r51 17 20 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.725 $Y=1.995
+ $X2=0.815 $Y2=1.995
r52 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.7
+ $X2=0.725 $Y2=2.7
r53 13 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=2.16
+ $X2=0.725 $Y2=1.995
r54 13 15 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.725 $Y=2.16
+ $X2=0.725 $Y2=2.7
r55 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=1.995 $X2=0.815 $Y2=1.995
r56 10 12 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.995
+ $X2=0.825 $Y2=2.16
r57 10 11 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.995
+ $X2=0.825 $Y2=1.83
r58 7 12 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.16
r59 3 11 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=1.83
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%B0 3 7 10 13 16 21 23 25 28
c54 7 0 1.38614e-19 $X=1.335 $Y=3.825
r55 23 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.25 $Y=1.6 $X2=1.53
+ $Y2=1.6
r56 21 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.33
+ $X2=1.165 $Y2=2.33
r57 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.165 $Y=1.685
+ $X2=1.25 $Y2=1.6
r58 19 21 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.165 $Y=1.685
+ $X2=1.165 $Y2=2.33
r59 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.53
+ $Y=1.6 $X2=1.53 $Y2=1.6
r60 16 18 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.47 $Y=1.6 $X2=1.53
+ $Y2=1.6
r61 11 13 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.335 $Y=2.56
+ $X2=1.47 $Y2=2.56
r62 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=2.485
+ $X2=1.47 $Y2=2.56
r63 9 16 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=1.765
+ $X2=1.47 $Y2=1.6
r64 9 10 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.47 $Y=1.765
+ $X2=1.47 $Y2=2.485
r65 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.635
+ $X2=1.335 $Y2=2.56
r66 5 7 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=1.335 $Y=2.635
+ $X2=1.335 $Y2=3.825
r67 1 16 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.325 $Y=1.435
+ $X2=1.47 $Y2=1.6
r68 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.325 $Y=1.435 $X2=1.325
+ $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%A_27_565# 1 2 11 15 16 19
r16 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=3.895
+ $X2=1.12 $Y2=4.575
r17 17 19 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=3.815 $X2=1.12
+ $Y2=3.895
r18 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.73
+ $X2=1.12 $Y2=3.815
r19 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.73
+ $X2=0.345 $Y2=3.73
r20 11 13 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.895
+ $X2=0.26 $Y2=4.575
r21 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.815
+ $X2=0.345 $Y2=3.73
r22 9 11 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=3.815 $X2=0.26
+ $Y2=3.895
r23 2 21 400 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r24 2 19 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.895
r25 1 13 400 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r26 1 11 400 $w=1.7e-07 $l=1.13077e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI21_L%Y 1 3 10 16 23 24 28 34
r46 26 34 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.845
+ $X2=1.55 $Y2=1.96
r47 26 28 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.55 $Y=1.845
+ $X2=1.55 $Y2=1.81
r48 25 28 0.486256 $w=1.7e-07 $l=5.05e-07 $layer=MET1_cond $X=1.55 $Y=1.305
+ $X2=1.55 $Y2=1.81
r49 24 31 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.195 $Y=1.22
+ $X2=1.05 $Y2=1.22
r50 23 25 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.465 $Y=1.22
+ $X2=1.55 $Y2=1.305
r51 23 24 0.259978 $w=1.7e-07 $l=2.7e-07 $layer=MET1_cond $X=1.465 $Y=1.22
+ $X2=1.195 $Y2=1.22
r52 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.55 $Y=3.555
+ $X2=1.55 $Y2=4.575
r53 16 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.96
+ $X2=1.55 $Y2=1.96
r54 16 19 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=1.55 $Y=1.96
+ $X2=1.55 $Y2=3.555
r55 13 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.05 $Y=1.22
+ $X2=1.05 $Y2=1.22
r56 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.05 $Y=0.74
+ $X2=1.05 $Y2=1.22
r57 3 21 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.575
r58 3 19 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.555
r59 1 10 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

