* File: sky130_osu_sc_18T_ls__and2_1.pex.spice
* Created: Fri Nov 12 14:13:20 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__AND2_1%GND 1 17 19 26 35 38
r36 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r37 24 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r38 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r39 17 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r40 17 19 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r41 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r42 1 26 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_1%VDD 1 2 17 21 25 32 40 42 45
r29 42 45 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r30 32 35 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r31 30 40 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r32 30 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r33 28 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r34 26 39 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r35 26 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r36 25 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r37 25 28 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r38 21 24 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r39 19 39 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r40 19 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r41 17 28 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r42 17 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r43 2 35 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r44 2 32 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r45 1 24 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r46 1 21 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_1%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=3.33
+ $X2=0.275 $Y2=3.33
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.765
+ $X2=0.27 $Y2=3.33
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.765 $X2=0.27 $Y2=2.765
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.765
+ $X2=0.475 $Y2=2.765
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=2.765
r38 5 7 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=4.585
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=2.765
r40 1 3 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_1%B 3 7 10 14 22
r41 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.96
+ $X2=0.955 $Y2=2.96
r42 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.96
r43 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.425
+ $X2=0.95 $Y2=2.96
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.425 $X2=0.95 $Y2=2.425
r45 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.59
r46 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.26
r47 7 12 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.59
r48 3 11 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_1%A_27_115# 1 3 11 15 16 18 19 24 26 27 32
+ 38 40 41 42
r69 41 42 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.545
+ $X2=0.65 $Y2=3.715
r70 36 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=0.61 $Y2=1.935
r71 36 38 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=1.43 $Y2=1.935
r72 32 34 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.69 $Y=3.795
+ $X2=0.69 $Y2=5.835
r73 32 42 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.795 $X2=0.69
+ $Y2=3.715
r74 28 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=2.02 $X2=0.61
+ $Y2=1.935
r75 28 41 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r76 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.61 $Y2=1.935
r77 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.345 $Y2=1.935
r78 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.345 $Y2=1.935
r79 22 24 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r80 21 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r81 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.81
+ $X2=1.352 $Y2=2.96
r82 16 21 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.412 $Y2=1.935
r83 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1 $X2=1.37
+ $Y2=2.81
r84 15 19 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.96
r85 9 21 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.412 $Y2=1.935
r86 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r87 3 34 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r88 3 32 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.795
r89 1 24 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_1%Y 1 3 10 16 26 29 32
r35 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r36 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r37 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r38 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r39 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r40 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r41 16 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r42 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r43 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r44 3 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r45 3 19 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r46 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

