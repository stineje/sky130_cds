* File: sky130_osu_sc_18T_ls__mux2_1.pxi.spice
* Created: Fri Nov 12 14:18:10 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%GND N_GND_M1004_s N_GND_M1004_b N_GND_c_15_p
+ GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_LS__MUX2_1%GND
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%VDD N_VDD_M1002_s N_VDD_M1002_b N_VDD_c_43_p
+ N_VDD_c_37_p VDD PM_SKY130_OSU_SC_18T_LS__MUX2_1%VDD
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%A_110_115# N_A_110_115#_M1004_d
+ N_A_110_115#_M1002_d N_A_110_115#_c_66_n N_A_110_115#_c_67_n
+ N_A_110_115#_M1003_g N_A_110_115#_M1001_g N_A_110_115#_c_71_n
+ N_A_110_115#_c_72_n N_A_110_115#_c_73_n N_A_110_115#_c_75_n
+ N_A_110_115#_c_76_n N_A_110_115#_c_77_n N_A_110_115#_c_78_n
+ PM_SKY130_OSU_SC_18T_LS__MUX2_1%A_110_115#
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%S0 N_S0_M1004_g N_S0_M1002_g N_S0_c_139_n
+ N_S0_c_146_n N_S0_c_147_n N_S0_c_150_n N_S0_M1005_g N_S0_M1000_g N_S0_c_142_n
+ N_S0_c_143_n S0 PM_SKY130_OSU_SC_18T_LS__MUX2_1%S0
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%A0 N_A0_M1003_s N_A0_M1005_s N_A0_c_200_n
+ N_A0_c_204_n N_A0_c_202_n N_A0_c_220_n N_A0_c_221_n A0
+ PM_SKY130_OSU_SC_18T_LS__MUX2_1%A0
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%Y N_Y_M1003_d N_Y_M1005_d N_Y_c_241_n
+ N_Y_c_243_n N_Y_c_244_n N_Y_c_245_n Y PM_SKY130_OSU_SC_18T_LS__MUX2_1%Y
x_PM_SKY130_OSU_SC_18T_LS__MUX2_1%A1 N_A1_M1000_d N_A1_M1001_d N_A1_c_278_n A1
+ PM_SKY130_OSU_SC_18T_LS__MUX2_1%A1
cc_1 N_GND_M1004_b N_A_110_115#_c_66_n 0.0249482f $X=-0.045 $Y=0 $X2=1.35
+ $Y2=1.79
cc_2 N_GND_M1004_b N_A_110_115#_c_67_n 0.0492602f $X=-0.045 $Y=0 $X2=1.78
+ $Y2=2.63
cc_3 N_GND_M1004_b N_A_110_115#_M1003_g 0.0282724f $X=-0.045 $Y=0 $X2=1.425
+ $Y2=1.075
cc_4 N_GND_c_4_p N_A_110_115#_M1003_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.425
+ $Y2=1.075
cc_5 N_GND_M1004_b N_A_110_115#_M1001_g 0.0124911f $X=-0.045 $Y=0 $X2=1.855
+ $Y2=4.585
cc_6 N_GND_M1004_b N_A_110_115#_c_71_n 0.0308275f $X=-0.045 $Y=0 $X2=1.09
+ $Y2=1.85
cc_7 N_GND_M1004_b N_A_110_115#_c_72_n 0.0294566f $X=-0.045 $Y=0 $X2=1.09
+ $Y2=2.69
cc_8 N_GND_M1004_b N_A_110_115#_c_73_n 0.0116497f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.825
cc_9 N_GND_c_4_p N_A_110_115#_c_73_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.69
+ $Y2=0.825
cc_10 N_GND_M1004_b N_A_110_115#_c_75_n 0.00868012f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=2.525
cc_11 N_GND_M1004_b N_A_110_115#_c_76_n 0.00123275f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=3.455
cc_12 N_GND_M1004_b N_A_110_115#_c_77_n 0.0152259f $X=-0.045 $Y=0 $X2=0.925
+ $Y2=1.85
cc_13 N_GND_M1004_b N_A_110_115#_c_78_n 0.0125647f $X=-0.045 $Y=0 $X2=0.925
+ $Y2=2.69
cc_14 N_GND_M1004_b N_S0_M1004_g 0.0669951f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_15 N_GND_c_15_p N_S0_M1004_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.075
cc_16 N_GND_c_4_p N_S0_M1004_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=1.075
cc_17 N_GND_M1004_b N_S0_M1002_g 0.0239334f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_18 N_GND_M1004_b N_S0_c_139_n 0.0722202f $X=-0.045 $Y=0 $X2=1.78 $Y2=2.27
cc_19 N_GND_M1004_b N_S0_M1000_g 0.0589672f $X=-0.045 $Y=0 $X2=1.855 $Y2=1.075
cc_20 N_GND_c_4_p N_S0_M1000_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.855 $Y2=1.075
cc_21 N_GND_M1004_b N_S0_c_142_n 0.0541332f $X=-0.045 $Y=0 $X2=0.55 $Y2=2.305
cc_22 N_GND_M1004_b N_S0_c_143_n 0.0261885f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.305
cc_23 N_GND_M1004_b N_A0_c_200_n 0.00901144f $X=-0.045 $Y=0 $X2=1.21 $Y2=0.825
cc_24 N_GND_c_4_p N_A0_c_200_n 0.00476261f $X=2.38 $Y=0.19 $X2=1.21 $Y2=0.825
cc_25 N_GND_M1004_b N_A0_c_202_n 0.0147072f $X=-0.045 $Y=0 $X2=1.265 $Y2=2.96
cc_26 N_GND_M1004_b A0 0.00472861f $X=-0.045 $Y=0 $X2=1.265 $Y2=2.96
cc_27 N_GND_M1004_b N_Y_c_241_n 0.00889125f $X=-0.045 $Y=0 $X2=1.64 $Y2=0.825
cc_28 N_GND_c_4_p N_Y_c_241_n 0.00475776f $X=2.38 $Y=0.19 $X2=1.64 $Y2=0.825
cc_29 N_GND_M1004_b N_Y_c_243_n 0.00910312f $X=-0.045 $Y=0 $X2=1.64 $Y2=2.22
cc_30 N_GND_M1004_b N_Y_c_244_n 0.00926001f $X=-0.045 $Y=0 $X2=1.64 $Y2=2.105
cc_31 N_GND_M1004_b N_Y_c_245_n 9.50189e-19 $X=-0.045 $Y=0 $X2=1.64 $Y2=1.48
cc_32 N_GND_M1004_b Y 0.00174495f $X=-0.045 $Y=0 $X2=1.64 $Y2=2.22
cc_33 N_GND_M1004_b N_A1_c_278_n 0.0671272f $X=-0.045 $Y=0 $X2=2.07 $Y2=0.825
cc_34 N_GND_c_4_p N_A1_c_278_n 0.00476261f $X=2.38 $Y=0.19 $X2=2.07 $Y2=0.825
cc_35 N_GND_M1004_b A1 0.0205786f $X=-0.045 $Y=0 $X2=2.07 $Y2=2.59
cc_36 N_VDD_M1002_b N_A_110_115#_M1001_g 0.0247516f $X=-0.045 $Y=2.905 $X2=1.855
+ $Y2=4.585
cc_37 N_VDD_c_37_p N_A_110_115#_M1001_g 0.00606474f $X=2.38 $Y=6.44 $X2=1.855
+ $Y2=4.585
cc_38 VDD N_A_110_115#_M1001_g 0.00468827f $X=2.38 $Y=6.42 $X2=1.855 $Y2=4.585
cc_39 N_VDD_M1002_b N_A_110_115#_c_76_n 0.00432876f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=3.455
cc_40 N_VDD_c_37_p N_A_110_115#_c_76_n 0.00757661f $X=2.38 $Y=6.44 $X2=0.69
+ $Y2=3.455
cc_41 VDD N_A_110_115#_c_76_n 0.00476261f $X=2.38 $Y=6.42 $X2=0.69 $Y2=3.455
cc_42 N_VDD_M1002_b N_S0_M1002_g 0.0135427f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_43 N_VDD_c_43_p N_S0_M1002_g 0.0127705f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_44 N_VDD_M1002_b N_S0_c_146_n 0.0650873f $X=-0.045 $Y=2.905 $X2=1.35
+ $Y2=6.235
cc_45 N_VDD_M1002_b N_S0_c_147_n 0.00987228f $X=-0.045 $Y=2.905 $X2=0.55
+ $Y2=6.235
cc_46 N_VDD_c_37_p N_S0_c_147_n 0.0405421f $X=2.38 $Y=6.44 $X2=0.55 $Y2=6.235
cc_47 VDD N_S0_c_147_n 0.0318799f $X=2.38 $Y=6.42 $X2=0.55 $Y2=6.235
cc_48 N_VDD_M1002_b N_S0_c_150_n 0.01729f $X=-0.045 $Y=2.905 $X2=1.425 $Y2=6.16
cc_49 N_VDD_M1002_s N_S0_c_143_n 0.0129471f $X=0.135 $Y=3.085 $X2=0.27 $Y2=2.305
cc_50 N_VDD_M1002_b N_S0_c_143_n 0.00842093f $X=-0.045 $Y=2.905 $X2=0.27
+ $Y2=2.305
cc_51 N_VDD_c_43_p N_S0_c_143_n 0.00370742f $X=0.26 $Y=4.135 $X2=0.27 $Y2=2.305
cc_52 N_VDD_M1002_s S0 0.00958477f $X=0.135 $Y=3.085 $X2=0.27 $Y2=3.33
cc_53 N_VDD_M1002_b S0 0.0097942f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=3.33
cc_54 N_VDD_c_43_p S0 0.00434783f $X=0.26 $Y=4.135 $X2=0.27 $Y2=3.33
cc_55 N_VDD_M1002_b N_A0_c_204_n 0.00108316f $X=-0.045 $Y=2.905 $X2=1.21
+ $Y2=3.455
cc_56 N_VDD_c_37_p N_A0_c_204_n 0.00757661f $X=2.38 $Y=6.44 $X2=1.21 $Y2=3.455
cc_57 VDD N_A0_c_204_n 0.00476261f $X=2.38 $Y=6.42 $X2=1.21 $Y2=3.455
cc_58 N_VDD_M1002_b N_A0_c_202_n 0.00309888f $X=-0.045 $Y=2.905 $X2=1.265
+ $Y2=2.96
cc_59 N_VDD_M1002_b A0 0.00892563f $X=-0.045 $Y=2.905 $X2=1.265 $Y2=2.96
cc_60 N_VDD_M1002_b N_Y_c_243_n 0.00488986f $X=-0.045 $Y=2.905 $X2=1.64 $Y2=2.22
cc_61 N_VDD_c_37_p N_Y_c_243_n 0.0075556f $X=2.38 $Y=6.44 $X2=1.64 $Y2=2.22
cc_62 VDD N_Y_c_243_n 0.00475776f $X=2.38 $Y=6.42 $X2=1.64 $Y2=2.22
cc_63 N_VDD_M1002_b N_A1_c_278_n 0.00998204f $X=-0.045 $Y=2.905 $X2=2.07
+ $Y2=0.825
cc_64 N_VDD_c_37_p N_A1_c_278_n 0.00757793f $X=2.38 $Y=6.44 $X2=2.07 $Y2=0.825
cc_65 VDD N_A1_c_278_n 0.00476261f $X=2.38 $Y=6.42 $X2=2.07 $Y2=0.825
cc_66 N_A_110_115#_c_71_n N_S0_M1004_g 0.0158178f $X=1.09 $Y=1.85 $X2=0.475
+ $Y2=1.075
cc_67 N_A_110_115#_c_73_n N_S0_M1004_g 0.0094215f $X=0.69 $Y=0.825 $X2=0.475
+ $Y2=1.075
cc_68 N_A_110_115#_c_75_n N_S0_M1004_g 0.00637747f $X=0.69 $Y=2.525 $X2=0.475
+ $Y2=1.075
cc_69 N_A_110_115#_c_77_n N_S0_M1004_g 0.00988145f $X=0.925 $Y=1.85 $X2=0.475
+ $Y2=1.075
cc_70 N_A_110_115#_c_72_n N_S0_M1002_g 0.0158178f $X=1.09 $Y=2.69 $X2=0.475
+ $Y2=4.585
cc_71 N_A_110_115#_c_76_n N_S0_M1002_g 0.00938463f $X=0.69 $Y=3.455 $X2=0.475
+ $Y2=4.585
cc_72 N_A_110_115#_c_78_n N_S0_M1002_g 0.00356688f $X=0.925 $Y=2.69 $X2=0.475
+ $Y2=4.585
cc_73 N_A_110_115#_c_66_n N_S0_c_139_n 0.0173318f $X=1.35 $Y=1.79 $X2=1.78
+ $Y2=2.27
cc_74 N_A_110_115#_c_71_n N_S0_c_139_n 0.0203852f $X=1.09 $Y=1.85 $X2=1.78
+ $Y2=2.27
cc_75 N_A_110_115#_c_72_n N_S0_c_139_n 0.0768879f $X=1.09 $Y=2.69 $X2=1.78
+ $Y2=2.27
cc_76 N_A_110_115#_c_75_n N_S0_c_139_n 0.013308f $X=0.69 $Y=2.525 $X2=1.78
+ $Y2=2.27
cc_77 N_A_110_115#_c_77_n N_S0_c_139_n 0.00273434f $X=0.925 $Y=1.85 $X2=1.78
+ $Y2=2.27
cc_78 N_A_110_115#_c_78_n N_S0_c_139_n 0.0028918f $X=0.925 $Y=2.69 $X2=1.78
+ $Y2=2.27
cc_79 N_A_110_115#_c_76_n N_S0_c_146_n 0.00326725f $X=0.69 $Y=3.455 $X2=1.35
+ $Y2=6.235
cc_80 N_A_110_115#_c_67_n N_S0_c_150_n 0.00910076f $X=1.78 $Y=2.63 $X2=1.425
+ $Y2=6.16
cc_81 N_A_110_115#_M1001_g N_S0_c_150_n 0.0195358f $X=1.855 $Y=4.585 $X2=1.425
+ $Y2=6.16
cc_82 N_A_110_115#_M1003_g N_S0_M1000_g 0.0322763f $X=1.425 $Y=1.075 $X2=1.855
+ $Y2=1.075
cc_83 N_A_110_115#_c_71_n N_S0_M1000_g 0.00120661f $X=1.09 $Y=1.85 $X2=1.855
+ $Y2=1.075
cc_84 N_A_110_115#_c_75_n N_S0_c_142_n 0.002234f $X=0.69 $Y=2.525 $X2=0.55
+ $Y2=2.305
cc_85 N_A_110_115#_c_75_n N_S0_c_143_n 0.0202899f $X=0.69 $Y=2.525 $X2=0.27
+ $Y2=2.305
cc_86 N_A_110_115#_c_76_n N_S0_c_143_n 0.0149462f $X=0.69 $Y=3.455 $X2=0.27
+ $Y2=2.305
cc_87 N_A_110_115#_c_78_n N_S0_c_143_n 0.0202357f $X=0.925 $Y=2.69 $X2=0.27
+ $Y2=2.305
cc_88 N_A_110_115#_M1002_d S0 0.00403387f $X=0.55 $Y=3.085 $X2=0.27 $Y2=3.33
cc_89 N_A_110_115#_c_76_n S0 0.00860476f $X=0.69 $Y=3.455 $X2=0.27 $Y2=3.33
cc_90 N_A_110_115#_c_73_n N_A0_c_200_n 0.0398625f $X=0.69 $Y=0.825 $X2=1.21
+ $Y2=0.825
cc_91 N_A_110_115#_c_66_n N_A0_c_202_n 0.0128445f $X=1.35 $Y=1.79 $X2=1.265
+ $Y2=2.96
cc_92 N_A_110_115#_c_67_n N_A0_c_202_n 0.0121009f $X=1.78 $Y=2.63 $X2=1.265
+ $Y2=2.96
cc_93 N_A_110_115#_M1003_g N_A0_c_202_n 0.00851711f $X=1.425 $Y=1.075 $X2=1.265
+ $Y2=2.96
cc_94 N_A_110_115#_c_71_n N_A0_c_202_n 0.0014863f $X=1.09 $Y=1.85 $X2=1.265
+ $Y2=2.96
cc_95 N_A_110_115#_c_72_n N_A0_c_202_n 0.0014863f $X=1.09 $Y=2.69 $X2=1.265
+ $Y2=2.96
cc_96 N_A_110_115#_c_73_n N_A0_c_202_n 0.00721095f $X=0.69 $Y=0.825 $X2=1.265
+ $Y2=2.96
cc_97 N_A_110_115#_c_75_n N_A0_c_202_n 0.019932f $X=0.69 $Y=2.525 $X2=1.265
+ $Y2=2.96
cc_98 N_A_110_115#_c_76_n N_A0_c_202_n 0.00714017f $X=0.69 $Y=3.455 $X2=1.265
+ $Y2=2.96
cc_99 N_A_110_115#_c_77_n N_A0_c_202_n 0.0240775f $X=0.925 $Y=1.85 $X2=1.265
+ $Y2=2.96
cc_100 N_A_110_115#_c_78_n N_A0_c_202_n 0.0247471f $X=0.925 $Y=2.69 $X2=1.265
+ $Y2=2.96
cc_101 N_A_110_115#_c_66_n N_A0_c_220_n 0.00212623f $X=1.35 $Y=1.79 $X2=1.237
+ $Y2=1.505
cc_102 N_A_110_115#_c_67_n N_A0_c_221_n 0.0017221f $X=1.78 $Y=2.63 $X2=1.237
+ $Y2=3.285
cc_103 N_A_110_115#_c_76_n N_A0_c_221_n 0.126077f $X=0.69 $Y=3.455 $X2=1.237
+ $Y2=3.285
cc_104 N_A_110_115#_c_67_n A0 0.00295688f $X=1.78 $Y=2.63 $X2=1.265 $Y2=2.96
cc_105 N_A_110_115#_c_72_n A0 0.00205826f $X=1.09 $Y=2.69 $X2=1.265 $Y2=2.96
cc_106 N_A_110_115#_c_76_n A0 0.00713596f $X=0.69 $Y=3.455 $X2=1.265 $Y2=2.96
cc_107 N_A_110_115#_c_78_n A0 0.00374574f $X=0.925 $Y=2.69 $X2=1.265 $Y2=2.96
cc_108 N_A_110_115#_M1003_g N_Y_c_241_n 0.00125663f $X=1.425 $Y=1.075 $X2=1.64
+ $Y2=0.825
cc_109 N_A_110_115#_c_67_n N_Y_c_243_n 0.0119679f $X=1.78 $Y=2.63 $X2=1.64
+ $Y2=2.22
cc_110 N_A_110_115#_M1001_g N_Y_c_243_n 0.00659127f $X=1.855 $Y=4.585 $X2=1.64
+ $Y2=2.22
cc_111 N_A_110_115#_M1003_g N_Y_c_244_n 0.00411772f $X=1.425 $Y=1.075 $X2=1.64
+ $Y2=2.105
cc_112 N_A_110_115#_M1003_g N_Y_c_245_n 0.00357441f $X=1.425 $Y=1.075 $X2=1.64
+ $Y2=1.48
cc_113 N_A_110_115#_c_67_n Y 5.02602e-19 $X=1.78 $Y=2.63 $X2=1.64 $Y2=2.22
cc_114 N_A_110_115#_c_67_n N_A1_c_278_n 0.0167254f $X=1.78 $Y=2.63 $X2=2.07
+ $Y2=0.825
cc_115 N_A_110_115#_c_67_n A1 0.0110708f $X=1.78 $Y=2.63 $X2=2.07 $Y2=2.59
cc_116 N_S0_c_146_n N_A0_c_204_n 0.00326725f $X=1.35 $Y=6.235 $X2=1.21 $Y2=3.455
cc_117 N_S0_M1004_g N_A0_c_202_n 8.64183e-19 $X=0.475 $Y=1.075 $X2=1.265
+ $Y2=2.96
cc_118 N_S0_M1002_g N_A0_c_202_n 6.2926e-19 $X=0.475 $Y=4.585 $X2=1.265 $Y2=2.96
cc_119 N_S0_c_139_n N_A0_c_202_n 0.011586f $X=1.78 $Y=2.27 $X2=1.265 $Y2=2.96
cc_120 N_S0_c_150_n N_A0_c_202_n 0.00636952f $X=1.425 $Y=6.16 $X2=1.265 $Y2=2.96
cc_121 N_S0_M1000_g N_A0_c_202_n 0.00404578f $X=1.855 $Y=1.075 $X2=1.265
+ $Y2=2.96
cc_122 N_S0_c_150_n A0 0.00517231f $X=1.425 $Y=6.16 $X2=1.265 $Y2=2.96
cc_123 N_S0_c_139_n N_Y_c_241_n 5.10857e-19 $X=1.78 $Y=2.27 $X2=1.64 $Y2=0.825
cc_124 N_S0_M1000_g N_Y_c_241_n 0.00132279f $X=1.855 $Y=1.075 $X2=1.64 $Y2=0.825
cc_125 N_S0_c_139_n N_Y_c_243_n 0.00869293f $X=1.78 $Y=2.27 $X2=1.64 $Y2=2.22
cc_126 N_S0_c_150_n N_Y_c_243_n 0.00194003f $X=1.425 $Y=6.16 $X2=1.64 $Y2=2.22
cc_127 N_S0_M1000_g N_Y_c_243_n 0.00117992f $X=1.855 $Y=1.075 $X2=1.64 $Y2=2.22
cc_128 N_S0_M1000_g N_Y_c_244_n 0.00873611f $X=1.855 $Y=1.075 $X2=1.64 $Y2=2.105
cc_129 N_S0_c_139_n N_Y_c_245_n 2.65725e-19 $X=1.78 $Y=2.27 $X2=1.64 $Y2=1.48
cc_130 N_S0_M1000_g N_Y_c_245_n 0.00370346f $X=1.855 $Y=1.075 $X2=1.64 $Y2=1.48
cc_131 N_S0_c_139_n Y 0.00459363f $X=1.78 $Y=2.27 $X2=1.64 $Y2=2.22
cc_132 N_S0_M1000_g Y 0.00192497f $X=1.855 $Y=1.075 $X2=1.64 $Y2=2.22
cc_133 N_S0_M1000_g N_A1_c_278_n 0.0267327f $X=1.855 $Y=1.075 $X2=2.07 $Y2=0.825
cc_134 N_S0_c_139_n A1 0.00214033f $X=1.78 $Y=2.27 $X2=2.07 $Y2=2.59
cc_135 N_A0_c_220_n N_Y_c_241_n 0.00379296f $X=1.237 $Y=1.505 $X2=1.64 $Y2=0.825
cc_136 N_A0_c_202_n N_Y_c_243_n 0.0552779f $X=1.265 $Y=2.96 $X2=1.64 $Y2=2.22
cc_137 A0 N_Y_c_243_n 0.0068435f $X=1.265 $Y=2.96 $X2=1.64 $Y2=2.22
cc_138 N_A0_c_202_n N_Y_c_244_n 0.0155159f $X=1.265 $Y=2.96 $X2=1.64 $Y2=2.105
cc_139 N_A0_c_220_n N_Y_c_245_n 0.00620538f $X=1.237 $Y=1.505 $X2=1.64 $Y2=1.48
cc_140 N_A0_c_202_n Y 0.00644986f $X=1.265 $Y=2.96 $X2=1.64 $Y2=2.22
cc_141 N_A0_c_202_n N_A1_c_278_n 0.00616016f $X=1.265 $Y=2.96 $X2=2.07 $Y2=0.825
cc_142 N_Y_c_243_n N_A1_c_278_n 0.0451561f $X=1.64 $Y=2.22 $X2=2.07 $Y2=0.825
cc_143 N_Y_c_244_n N_A1_c_278_n 0.0147366f $X=1.64 $Y=2.105 $X2=2.07 $Y2=0.825
cc_144 N_Y_c_245_n N_A1_c_278_n 0.00591748f $X=1.64 $Y=1.48 $X2=2.07 $Y2=0.825
cc_145 Y N_A1_c_278_n 0.00589642f $X=1.64 $Y=2.22 $X2=2.07 $Y2=0.825
cc_146 N_Y_c_243_n A1 0.00751022f $X=1.64 $Y=2.22 $X2=2.07 $Y2=2.59
cc_147 Y A1 0.00272809f $X=1.64 $Y=2.22 $X2=2.07 $Y2=2.59
