* File: sky130_osu_sc_18T_ls__mux2_1.spice
* Created: Thu Oct 29 17:37:02 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ls__mux2_1.pex.spice"
.subckt sky130_osu_sc_18T_ls__mux2_1  GND VDD S0 A0 Y A1
* 
* A1	A1
* Y	Y
* A0	A0
* S0	S0
* VDD	VDD
* GND	GND
MM1004 N_A_110_115#_M1004_d N_S0_M1004_g N_GND_M1004_s N_GND_M1004_b NSHORT
+ L=0.15 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1003_d N_A_110_115#_M1003_g N_A0_M1003_s N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A1_M1000_d N_S0_M1000_g N_Y_M1003_d N_GND_M1004_b NSHORT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_110_115#_M1002_d N_S0_M1002_g N_VDD_M1002_s N_VDD_M1002_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1005 N_Y_M1005_d N_S0_M1005_g N_A0_M1005_s N_VDD_M1002_b PHIGHVT L=0.15 W=3
+ AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2 SB=75000.6
+ A=0.45 P=6.3 MULT=1
MM1001 N_A1_M1001_d N_A_110_115#_M1001_g N_Y_M1005_d N_VDD_M1002_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1002_b NWDIODE A=10.678 P=13.22
pX7_noxref noxref_8 S0 S0 PROBETYPE=1
pX8_noxref noxref_9 A0 A0 PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
pX10_noxref noxref_11 A1 A1 PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__mux2_1.pxi.spice"
*
.ends
*
*
