* File: sky130_osu_sc_15T_hs__nand2_l.pxi.spice
* Created: Fri Nov 12 14:31:49 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__NAND2_L%GND N_GND_M1000_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_9_p GND N_GND_c_3_p PM_SKY130_OSU_SC_15T_HS__NAND2_L%GND
x_PM_SKY130_OSU_SC_15T_HS__NAND2_L%VDD N_VDD_M1001_s N_VDD_M1003_d N_VDD_M1001_b
+ N_VDD_c_26_p N_VDD_c_27_p N_VDD_c_33_p VDD N_VDD_c_28_p
+ PM_SKY130_OSU_SC_15T_HS__NAND2_L%VDD
x_PM_SKY130_OSU_SC_15T_HS__NAND2_L%A N_A_M1002_g N_A_M1001_g N_A_c_44_n
+ N_A_c_45_n A PM_SKY130_OSU_SC_15T_HS__NAND2_L%A
x_PM_SKY130_OSU_SC_15T_HS__NAND2_L%B N_B_M1000_g N_B_M1003_g N_B_c_72_n
+ N_B_c_74_n N_B_c_75_n B PM_SKY130_OSU_SC_15T_HS__NAND2_L%B
x_PM_SKY130_OSU_SC_15T_HS__NAND2_L%Y N_Y_M1002_s N_Y_M1001_d N_Y_c_102_n
+ N_Y_c_105_n N_Y_c_106_n N_Y_c_107_n Y N_Y_c_109_n
+ PM_SKY130_OSU_SC_15T_HS__NAND2_L%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.101322f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.85
cc_4 N_GND_M1002_b N_A_M1001_g 0.00342256f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.195
cc_5 N_GND_M1002_b N_A_c_44_n 0.0490341f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.425
cc_6 N_GND_M1002_b N_A_c_45_n 0.00856875f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.425
cc_7 N_GND_M1002_b N_B_M1000_g 0.0392257f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.85
cc_8 N_GND_c_2_p N_B_M1000_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.85
cc_9 N_GND_c_9_p N_B_M1000_g 0.00502587f $X=1.05 $Y=0.74 $X2=0.835 $Y2=0.85
cc_10 N_GND_c_3_p N_B_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.85
cc_11 N_GND_M1002_b N_B_M1003_g 0.0497877f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.195
cc_12 N_GND_M1002_b N_B_c_72_n 0.0353806f $X=-0.045 $Y=0 $X2=0.915 $Y2=1.675
cc_13 N_GND_c_9_p N_B_c_72_n 0.00239673f $X=1.05 $Y=0.74 $X2=0.915 $Y2=1.675
cc_14 N_GND_M1002_b N_B_c_74_n 0.0293783f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.7
cc_15 N_GND_M1002_b N_B_c_75_n 0.0123076f $X=-0.045 $Y=0 $X2=1.06 $Y2=1.675
cc_16 N_GND_M1002_b B 0.00499588f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.7
cc_17 N_GND_M1002_b N_Y_c_102_n 0.00945075f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.74
cc_18 N_GND_c_2_p N_Y_c_102_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26 $Y2=0.74
cc_19 N_GND_c_3_p N_Y_c_102_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26 $Y2=0.74
cc_20 N_GND_M1002_b N_Y_c_105_n 0.00860362f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.33
cc_21 N_GND_M1002_b N_Y_c_106_n 0.0101912f $X=-0.045 $Y=0 $X2=0.605 $Y2=1.22
cc_22 N_GND_M1002_b N_Y_c_107_n 0.0206417f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.22
cc_23 N_GND_M1002_b Y 0.0166407f $X=-0.045 $Y=0 $X2=0.68 $Y2=2.09
cc_24 N_GND_M1002_b N_Y_c_109_n 0.00535447f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.33
cc_25 N_VDD_M1001_b N_A_M1001_g 0.0762016f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=4.195
cc_26 N_VDD_c_26_p N_A_M1001_g 0.00751602f $X=0.26 $Y=4.565 $X2=0.475 $Y2=4.195
cc_27 N_VDD_c_27_p N_A_M1001_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475 $Y2=4.195
cc_28 N_VDD_c_28_p N_A_M1001_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=4.195
cc_29 N_VDD_M1001_b N_A_c_45_n 0.0153337f $X=-0.045 $Y=2.645 $X2=0.32 $Y2=2.425
cc_30 N_VDD_M1001_b A 0.0208751f $X=-0.045 $Y=2.645 $X2=0.32 $Y2=3.07
cc_31 N_VDD_M1001_b N_B_M1003_g 0.0831768f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=4.195
cc_32 N_VDD_c_27_p N_B_M1003_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905 $Y2=4.195
cc_33 N_VDD_c_33_p N_B_M1003_g 0.00751602f $X=1.12 $Y=4.565 $X2=0.905 $Y2=4.195
cc_34 N_VDD_c_28_p N_B_M1003_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.905 $Y2=4.195
cc_35 N_VDD_M1001_b N_B_c_74_n 0.00391589f $X=-0.045 $Y=2.645 $X2=1.06 $Y2=2.7
cc_36 N_VDD_M1001_b B 0.0168801f $X=-0.045 $Y=2.645 $X2=1.06 $Y2=2.7
cc_37 N_VDD_M1001_b N_Y_c_105_n 0.0216012f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.33
cc_38 N_VDD_c_27_p N_Y_c_105_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69 $Y2=2.33
cc_39 N_VDD_c_28_p N_Y_c_105_n 0.00434939f $X=1.02 $Y=5.36 $X2=0.69 $Y2=2.33
cc_40 N_A_M1002_g N_B_M1000_g 0.0874628f $X=0.475 $Y=0.85 $X2=0.835 $Y2=0.85
cc_41 N_A_M1002_g N_B_M1003_g 0.10588f $X=0.475 $Y=0.85 $X2=0.905 $Y2=4.195
cc_42 N_A_M1002_g N_B_c_74_n 0.00248145f $X=0.475 $Y=0.85 $X2=1.06 $Y2=2.7
cc_43 N_A_M1002_g N_B_c_75_n 0.00282768f $X=0.475 $Y=0.85 $X2=1.06 $Y2=1.675
cc_44 N_A_M1002_g N_Y_c_102_n 0.00971844f $X=0.475 $Y=0.85 $X2=0.26 $Y2=0.74
cc_45 N_A_M1002_g N_Y_c_105_n 0.0202901f $X=0.475 $Y=0.85 $X2=0.69 $Y2=2.33
cc_46 N_A_c_45_n N_Y_c_105_n 0.0513069f $X=0.32 $Y=2.425 $X2=0.69 $Y2=2.33
cc_47 A N_Y_c_105_n 0.00831114f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.33
cc_48 N_A_M1002_g N_Y_c_106_n 0.0136921f $X=0.475 $Y=0.85 $X2=0.605 $Y2=1.22
cc_49 N_A_M1002_g N_Y_c_107_n 0.00393078f $X=0.475 $Y=0.85 $X2=0.405 $Y2=1.22
cc_50 N_A_M1002_g Y 0.0125133f $X=0.475 $Y=0.85 $X2=0.68 $Y2=2.09
cc_51 N_A_M1002_g N_Y_c_109_n 0.00216533f $X=0.475 $Y=0.85 $X2=0.69 $Y2=2.33
cc_52 N_A_c_44_n N_Y_c_109_n 0.00278592f $X=0.32 $Y=2.425 $X2=0.69 $Y2=2.33
cc_53 N_A_c_45_n N_Y_c_109_n 0.00474021f $X=0.32 $Y=2.425 $X2=0.69 $Y2=2.33
cc_54 A N_Y_c_109_n 0.00152954f $X=0.32 $Y=3.07 $X2=0.69 $Y2=2.33
cc_55 N_B_M1003_g N_Y_c_105_n 0.0259548f $X=0.905 $Y=4.195 $X2=0.69 $Y2=2.33
cc_56 N_B_c_74_n N_Y_c_105_n 0.0295869f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_57 N_B_c_75_n N_Y_c_105_n 5.24123e-19 $X=1.06 $Y=1.675 $X2=0.69 $Y2=2.33
cc_58 B N_Y_c_105_n 0.00831114f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_59 N_B_M1000_g N_Y_c_106_n 0.00853825f $X=0.835 $Y=0.85 $X2=0.605 $Y2=1.22
cc_60 N_B_M1000_g Y 0.00770103f $X=0.835 $Y=0.85 $X2=0.68 $Y2=2.09
cc_61 N_B_M1003_g Y 0.00539744f $X=0.905 $Y=4.195 $X2=0.68 $Y2=2.09
cc_62 N_B_c_72_n Y 0.00401356f $X=0.915 $Y=1.675 $X2=0.68 $Y2=2.09
cc_63 N_B_c_74_n Y 0.0183986f $X=1.06 $Y=2.7 $X2=0.68 $Y2=2.09
cc_64 N_B_c_75_n Y 0.0141623f $X=1.06 $Y=1.675 $X2=0.68 $Y2=2.09
cc_65 N_B_M1003_g N_Y_c_109_n 0.00341272f $X=0.905 $Y=4.195 $X2=0.69 $Y2=2.33
cc_66 N_B_c_72_n N_Y_c_109_n 0.00144278f $X=0.915 $Y=1.675 $X2=0.69 $Y2=2.33
cc_67 N_B_c_74_n N_Y_c_109_n 0.00640429f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
cc_68 N_B_c_75_n N_Y_c_109_n 0.00194461f $X=1.06 $Y=1.675 $X2=0.69 $Y2=2.33
cc_69 B N_Y_c_109_n 0.00280435f $X=1.06 $Y=2.7 $X2=0.69 $Y2=2.33
