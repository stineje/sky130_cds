* File: sky130_osu_sc_12T_hs__addh_1.pex.spice
* Created: Fri Nov 12 15:06:27 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%GND 1 2 45 47 55 57 70 86 88
r104 86 88 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r105 72 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r106 68 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r107 68 70 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.755
r108 58 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r109 57 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r110 53 81 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r111 53 55 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.755
r112 47 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r113 45 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r114 45 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r115 45 72 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r116 45 57 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r117 45 58 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r118 45 47 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r119 2 70 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.755
r120 1 55 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%VDD 1 2 3 37 39 46 50 56 58 66 72 80 84
r57 80 84 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=3.74 $Y2=4.287
r58 72 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=4.25
+ $X2=3.74 $Y2=4.25
r59 70 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=4.287
+ $X2=3.05 $Y2=4.287
r60 70 72 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=4.287
+ $X2=3.74 $Y2=4.287
r61 66 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.05 $Y=2.955
+ $X2=3.05 $Y2=3.635
r62 64 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=4.135
+ $X2=3.05 $Y2=4.287
r63 64 69 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.05 $Y=4.135 $X2=3.05
+ $Y2=3.635
r64 61 63 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=4.287
+ $X2=2.38 $Y2=4.287
r65 59 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=4.287
+ $X2=1.61 $Y2=4.287
r66 59 61 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=4.287
+ $X2=1.7 $Y2=4.287
r67 58 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=4.287
+ $X2=3.05 $Y2=4.287
r68 58 63 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=4.287
+ $X2=2.38 $Y2=4.287
r69 54 76 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=4.135
+ $X2=1.61 $Y2=4.287
r70 54 56 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.61 $Y=4.135
+ $X2=1.61 $Y2=3.295
r71 51 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=4.287
+ $X2=0.75 $Y2=4.287
r72 51 53 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=4.287
+ $X2=1.02 $Y2=4.287
r73 50 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=4.287
+ $X2=1.61 $Y2=4.287
r74 50 53 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=4.287
+ $X2=1.02 $Y2=4.287
r75 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.75 $Y=2.955
+ $X2=0.75 $Y2=3.635
r76 44 75 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=4.135
+ $X2=0.75 $Y2=4.287
r77 44 49 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.75 $Y=4.135 $X2=0.75
+ $Y2=3.635
r78 41 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r79 39 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=4.287
+ $X2=0.75 $Y2=4.287
r80 39 41 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=4.287
+ $X2=0.34 $Y2=4.287
r81 37 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r82 37 78 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r83 37 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r84 37 61 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r85 37 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r86 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r87 3 69 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=2.605 $X2=3.05 $Y2=3.635
r88 3 66 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=2.605 $X2=3.05 $Y2=2.955
r89 2 56 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.605 $X2=1.61 $Y2=3.295
r90 1 49 400 $w=1.7e-07 $l=1.12557e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.75 $Y2=3.635
r91 1 46 400 $w=1.7e-07 $l=4.38748e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.75 $Y2=2.955
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%CON 1 7 8 23 26 29 30 36 37 40 44 46 48
+ 51 53 54 58 63 64 68 69 74 77 82 83 88 91
c142 91 0 2.7119e-19 $X=3.42 $Y=1.37
c143 83 0 1.57622e-19 $X=0.78 $Y=1.37
c144 69 0 4.75316e-20 $X=2.99 $Y=0.635
c145 51 0 1.92558e-19 $X=3.42 $Y=1.285
r146 83 85 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.37
+ $X2=0.635 $Y2=1.37
r147 82 88 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.37
+ $X2=2.62 $Y2=1.37
r148 82 83 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.37
+ $X2=0.78 $Y2=1.37
r149 77 80 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.85 $Y=0.635
+ $X2=3.85 $Y2=0.755
r150 76 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.37
+ $X2=3.42 $Y2=1.37
r151 69 72 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.99 $Y=0.635
+ $X2=2.99 $Y2=0.755
r152 67 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.37
+ $X2=2.62 $Y2=1.37
r153 63 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.37
+ $X2=0.635 $Y2=1.37
r154 63 64 4.99498 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=1.385
+ $X2=0.55 $Y2=1.385
r155 58 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.84 $Y=2.955
+ $X2=3.84 $Y2=3.635
r156 56 58 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.84 $Y=2.555
+ $X2=3.84 $Y2=2.955
r157 55 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=0.635
+ $X2=3.42 $Y2=0.635
r158 54 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.85 $Y2=0.635
r159 54 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.505 $Y2=0.635
r160 51 76 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.285
+ $X2=3.42 $Y2=1.37
r161 51 53 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.42 $Y=1.285
+ $X2=3.42 $Y2=0.755
r162 50 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.72
+ $X2=3.42 $Y2=0.635
r163 50 53 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.42 $Y=0.72
+ $X2=3.42 $Y2=0.755
r164 49 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.635
+ $X2=2.99 $Y2=0.635
r165 48 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.635
+ $X2=3.42 $Y2=0.635
r166 48 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.335 $Y=0.635
+ $X2=3.075 $Y2=0.635
r167 47 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.47
+ $X2=2.62 $Y2=2.47
r168 46 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.47
+ $X2=3.84 $Y2=2.555
r169 46 47 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.47
+ $X2=2.705 $Y2=2.47
r170 45 67 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.37
+ $X2=2.62 $Y2=1.37
r171 44 76 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.37
+ $X2=3.42 $Y2=1.37
r172 44 45 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.37
+ $X2=2.705 $Y2=1.37
r173 40 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.62 $Y=2.955
+ $X2=2.62 $Y2=3.635
r174 38 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.555
+ $X2=2.62 $Y2=2.47
r175 38 40 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.62 $Y=2.555
+ $X2=2.62 $Y2=2.955
r176 37 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.385
+ $X2=2.62 $Y2=2.47
r177 36 67 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.455
+ $X2=2.62 $Y2=1.37
r178 36 37 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.455
+ $X2=2.62 $Y2=2.385
r179 34 64 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.35 $Y=1.4 $X2=0.55
+ $Y2=1.4
r180 29 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.4 $X2=0.35 $Y2=1.4
r181 29 31 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.4
+ $X2=0.382 $Y2=1.565
r182 29 30 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.4
+ $X2=0.382 $Y2=1.235
r183 26 31 856.319 $w=1.5e-07 $l=1.67e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=1.565
r184 23 30 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=0.85
+ $X2=0.475 $Y2=1.235
r185 8 60 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=2.605 $X2=3.84 $Y2=3.635
r186 8 58 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=2.605 $X2=3.84 $Y2=2.955
r187 7 42 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.605 $X2=2.62 $Y2=3.635
r188 7 40 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.605 $X2=2.62 $Y2=2.955
r189 1 80 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.755
r190 1 53 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=0.755
r191 1 72 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%B 3 7 11 15 18 22 25 30 39 42 44
c101 44 0 4.99902e-20 $X=3.21 $Y=1.74
c102 22 0 1.42567e-19 $X=3.205 $Y=1.74
c103 18 0 1.57622e-19 $X=0.905 $Y=1.74
c104 11 0 4.75316e-20 $X=3.205 $Y=0.85
r105 41 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=3.205 $Y=1.74
+ $X2=3.21 $Y2=1.74
r106 41 42 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.205 $Y=1.74
+ $X2=3.06 $Y2=1.74
r107 39 42 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=1.742
+ $X2=3.06 $Y2=1.742
r108 37 39 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=1.74
+ $X2=1.05 $Y2=1.74
r109 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=1.74
+ $X2=3.205 $Y2=1.74
r110 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=1.74
+ $X2=0.905 $Y2=1.74
r111 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.74 $X2=3.205 $Y2=1.74
r112 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.74
+ $X2=3.205 $Y2=1.905
r113 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.74 $X2=0.905 $Y2=1.74
r114 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.74
+ $X2=0.905 $Y2=1.905
r115 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.74
+ $X2=0.905 $Y2=1.575
r116 15 23 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.265 $Y=3.235
+ $X2=3.265 $Y2=1.905
r117 9 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.575
+ $X2=3.205 $Y2=1.74
r118 9 11 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=3.205 $Y=1.575
+ $X2=3.205 $Y2=0.85
r119 7 20 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.965 $Y=3.235
+ $X2=0.965 $Y2=1.905
r120 3 19 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=0.965 $Y=0.85
+ $X2=0.965 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%A 3 7 11 15 18 22 26 31 40 42 43
c88 22 0 1.74252e-19 $X=3.685 $Y=2.11
r89 42 43 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.11
+ $X2=3.54 $Y2=2.11
r90 40 43 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.107
+ $X2=3.54 $Y2=2.107
r91 38 40 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.11
+ $X2=1.53 $Y2=2.11
r92 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.11
+ $X2=3.685 $Y2=2.11
r93 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.11
+ $X2=1.385 $Y2=2.11
r94 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.11 $X2=3.685 $Y2=2.11
r95 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.11
+ $X2=3.685 $Y2=2.275
r96 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.11
+ $X2=3.685 $Y2=1.945
r97 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.11 $X2=1.385 $Y2=2.11
r98 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.11
+ $X2=1.385 $Y2=2.275
r99 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.11
+ $X2=1.385 $Y2=1.945
r100 15 23 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=3.635 $Y=0.85
+ $X2=3.635 $Y2=1.945
r101 11 24 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.625 $Y=3.235
+ $X2=3.625 $Y2=2.275
r102 7 20 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.395 $Y=3.235
+ $X2=1.395 $Y2=2.275
r103 3 19 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=1.325 $Y=0.85
+ $X2=1.325 $Y2=1.945
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%A_208_521# 1 3 10 13 15 17 19 21 22 24
+ 26 29 31 36 37 40 42 43 46 49 51
c113 29 0 2.52869e-20 $X=2.835 $Y=3.235
c114 22 0 9.69384e-20 $X=2.7 $Y=1.32
r115 51 53 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.475
+ $X2=1.825 $Y2=1.475
r116 50 51 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.475
+ $X2=1.725 $Y2=1.475
r117 48 51 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.64
+ $X2=1.725 $Y2=1.475
r118 48 49 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=1.64
+ $X2=1.725 $Y2=2.445
r119 44 50 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.31
+ $X2=1.54 $Y2=1.475
r120 44 46 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.54 $Y=1.31
+ $X2=1.54 $Y2=0.755
r121 42 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=2.53
+ $X2=1.725 $Y2=2.445
r122 42 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=2.53
+ $X2=1.265 $Y2=2.53
r123 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=2.615
+ $X2=1.265 $Y2=2.53
r124 38 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.18 $Y=2.615
+ $X2=1.18 $Y2=3.295
r125 34 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.475 $X2=1.825 $Y2=1.475
r126 34 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.475
+ $X2=1.825 $Y2=1.64
r127 31 34 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.32
+ $X2=1.825 $Y2=1.475
r128 27 29 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.835 $Y=2.265
+ $X2=2.835 $Y2=3.235
r129 24 26 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.775 $Y=1.245
+ $X2=2.775 $Y2=0.85
r130 23 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.32
+ $X2=2.285 $Y2=1.32
r131 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.32
+ $X2=2.775 $Y2=1.245
r132 22 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.32 $X2=2.36
+ $Y2=1.32
r133 19 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.245
+ $X2=2.285 $Y2=1.32
r134 19 21 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.285 $Y=1.245
+ $X2=2.285 $Y2=0.85
r135 18 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.19
+ $X2=1.885 $Y2=2.19
r136 17 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.19
+ $X2=2.835 $Y2=2.265
r137 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.19 $X2=1.96
+ $Y2=2.19
r138 16 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.32
+ $X2=1.825 $Y2=1.32
r139 15 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.32
+ $X2=2.285 $Y2=1.32
r140 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.32
+ $X2=1.96 $Y2=1.32
r141 11 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.265
+ $X2=1.885 $Y2=2.19
r142 11 13 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.885 $Y=2.265
+ $X2=1.885 $Y2=3.235
r143 10 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.115
+ $X2=1.885 $Y2=2.19
r144 10 35 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.115
+ $X2=1.885 $Y2=1.64
r145 3 40 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.605 $X2=1.18 $Y2=3.295
r146 1 46 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.4 $Y=0.575
+ $X2=1.54 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%S 1 3 10 16 26 29 32
r34 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=2.735
+ $X2=0.26 $Y2=2.85
r35 24 26 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=2.735
+ $X2=0.26 $Y2=1.905
r36 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.11
+ $X2=0.26 $Y2=0.995
r37 23 26 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.11
+ $X2=0.26 $Y2=1.905
r38 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r39 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.85
+ $X2=0.26 $Y2=2.85
r40 16 19 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.26 $Y=2.85
+ $X2=0.26 $Y2=2.955
r41 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=0.995
+ $X2=0.26 $Y2=0.995
r42 10 13 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.26 $Y=0.755
+ $X2=0.26 $Y2=0.995
r43 3 21 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r44 3 19 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r45 1 10 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__ADDH_1%CO 1 3 11 15 23 26 27 30
c53 26 0 2.52869e-20 $X=2.175 $Y=2.48
r54 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.48
+ $X2=2.175 $Y2=2.48
r55 26 28 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.48
+ $X2=2.137 $Y2=2.565
r56 26 27 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.48
+ $X2=2.137 $Y2=2.395
r57 21 23 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=0.992
+ $X2=2.175 $Y2=0.992
r58 19 23 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.175 $Y=1.08
+ $X2=2.175 $Y2=0.992
r59 19 27 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.08
+ $X2=2.175 $Y2=2.395
r60 15 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.1 $Y=2.955 $X2=2.1
+ $Y2=3.635
r61 15 28 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.1 $Y=2.955 $X2=2.1
+ $Y2=2.565
r62 9 21 0.89264 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.07 $Y=0.905 $X2=2.07
+ $Y2=0.992
r63 9 11 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.07 $Y=0.905 $X2=2.07
+ $Y2=0.755
r64 3 17 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=2.605 $X2=2.1 $Y2=3.635
r65 3 15 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=2.605 $X2=2.1 $Y2=2.955
r66 1 11 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.755
.ends

