magic
tech sky130A
magscale 1 2
timestamp 1612373083
<< nwell >>
rect -10 529 1741 1119
<< nmoslvt >>
rect 80 115 110 199
rect 152 115 182 199
rect 356 115 386 243
rect 428 115 458 243
rect 548 115 578 243
rect 620 115 650 243
rect 706 115 736 243
rect 778 115 808 243
rect 898 115 928 243
rect 970 115 1000 243
rect 1056 115 1086 243
rect 1246 115 1276 199
rect 1318 115 1348 199
rect 1522 115 1552 243
rect 1608 115 1638 243
<< pmos >>
rect 80 713 110 965
rect 166 713 196 965
rect 356 565 386 965
rect 428 565 458 965
rect 548 565 578 965
rect 620 565 650 965
rect 706 565 736 965
rect 778 565 808 965
rect 898 565 928 965
rect 970 565 1000 965
rect 1056 565 1086 965
rect 1246 713 1276 965
rect 1332 713 1362 965
rect 1522 565 1552 965
rect 1608 565 1638 965
<< ndiff >>
rect 303 215 356 243
rect 27 165 80 199
rect 27 131 35 165
rect 69 131 80 165
rect 27 115 80 131
rect 110 115 152 199
rect 182 165 235 199
rect 182 131 193 165
rect 227 131 235 165
rect 182 115 235 131
rect 303 131 311 215
rect 345 131 356 215
rect 303 115 356 131
rect 386 115 428 243
rect 458 215 548 243
rect 458 131 469 215
rect 537 131 548 215
rect 458 115 548 131
rect 578 115 620 243
rect 650 165 706 243
rect 650 131 661 165
rect 695 131 706 165
rect 650 115 706 131
rect 736 115 778 243
rect 808 215 898 243
rect 808 131 819 215
rect 887 131 898 215
rect 808 115 898 131
rect 928 115 970 243
rect 1000 215 1056 243
rect 1000 131 1011 215
rect 1045 131 1056 215
rect 1000 115 1056 131
rect 1086 215 1139 243
rect 1086 131 1097 215
rect 1131 131 1139 215
rect 1086 115 1139 131
rect 1193 165 1246 199
rect 1193 131 1201 165
rect 1235 131 1246 165
rect 1193 115 1246 131
rect 1276 115 1318 199
rect 1348 165 1401 199
rect 1348 131 1359 165
rect 1393 131 1401 165
rect 1348 115 1401 131
rect 1469 165 1522 243
rect 1469 131 1477 165
rect 1511 131 1522 165
rect 1469 115 1522 131
rect 1552 165 1608 243
rect 1552 131 1563 165
rect 1597 131 1608 165
rect 1552 115 1608 131
rect 1638 165 1691 243
rect 1638 131 1649 165
rect 1683 131 1691 165
rect 1638 115 1691 131
<< pdiff >>
rect 27 949 80 965
rect 27 877 35 949
rect 69 877 80 949
rect 27 713 80 877
rect 110 949 166 965
rect 110 877 121 949
rect 155 877 166 949
rect 110 713 166 877
rect 196 949 249 965
rect 196 877 207 949
rect 241 877 249 949
rect 196 713 249 877
rect 303 949 356 965
rect 303 673 311 949
rect 345 673 356 949
rect 303 565 356 673
rect 386 565 428 965
rect 458 949 548 965
rect 458 605 469 949
rect 537 605 548 949
rect 458 565 548 605
rect 578 565 620 965
rect 650 949 706 965
rect 650 673 661 949
rect 695 673 706 949
rect 650 565 706 673
rect 736 565 778 965
rect 808 949 898 965
rect 808 673 819 949
rect 887 673 898 949
rect 808 565 898 673
rect 928 565 970 965
rect 1000 949 1056 965
rect 1000 605 1011 949
rect 1045 605 1056 949
rect 1000 565 1056 605
rect 1086 949 1139 965
rect 1086 605 1097 949
rect 1131 605 1139 949
rect 1193 949 1246 965
rect 1193 877 1201 949
rect 1235 877 1246 949
rect 1193 713 1246 877
rect 1276 949 1332 965
rect 1276 877 1287 949
rect 1321 877 1332 949
rect 1276 713 1332 877
rect 1362 949 1415 965
rect 1362 877 1373 949
rect 1407 877 1415 949
rect 1362 713 1415 877
rect 1469 949 1522 965
rect 1469 809 1477 949
rect 1511 809 1522 949
rect 1086 565 1139 605
rect 1469 565 1522 809
rect 1552 949 1608 965
rect 1552 809 1563 949
rect 1597 809 1608 949
rect 1552 565 1608 809
rect 1638 949 1691 965
rect 1638 809 1649 949
rect 1683 809 1691 949
rect 1638 565 1691 809
<< ndiffc >>
rect 35 131 69 165
rect 193 131 227 165
rect 311 131 345 215
rect 469 131 537 215
rect 661 131 695 165
rect 819 131 887 215
rect 1011 131 1045 215
rect 1097 131 1131 215
rect 1201 131 1235 165
rect 1359 131 1393 165
rect 1477 131 1511 165
rect 1563 131 1597 165
rect 1649 131 1683 165
<< pdiffc >>
rect 35 877 69 949
rect 121 877 155 949
rect 207 877 241 949
rect 311 673 345 949
rect 469 605 537 949
rect 661 673 695 949
rect 819 673 887 949
rect 1011 605 1045 949
rect 1097 605 1131 949
rect 1201 877 1235 949
rect 1287 877 1321 949
rect 1373 877 1407 949
rect 1477 809 1511 949
rect 1563 809 1597 949
rect 1649 809 1683 949
<< psubdiff >>
rect 26 27 50 61
rect 84 27 108 61
rect 162 27 186 61
rect 220 27 244 61
rect 298 27 322 61
rect 356 27 380 61
rect 434 27 458 61
rect 492 27 516 61
rect 570 27 594 61
rect 628 27 652 61
rect 706 27 730 61
rect 764 27 788 61
rect 842 27 866 61
rect 900 27 924 61
rect 978 27 1002 61
rect 1036 27 1060 61
rect 1114 27 1138 61
rect 1172 27 1196 61
rect 1250 27 1274 61
rect 1308 27 1332 61
rect 1386 27 1410 61
rect 1444 27 1468 61
rect 1522 27 1546 61
rect 1580 27 1604 61
<< nsubdiff >>
rect 26 1049 50 1083
rect 84 1049 108 1083
rect 162 1049 186 1083
rect 220 1049 244 1083
rect 298 1049 322 1083
rect 356 1049 380 1083
rect 434 1049 458 1083
rect 492 1049 516 1083
rect 570 1049 594 1083
rect 628 1049 652 1083
rect 706 1049 730 1083
rect 764 1049 788 1083
rect 842 1049 866 1083
rect 900 1049 924 1083
rect 978 1049 1002 1083
rect 1036 1049 1060 1083
rect 1114 1049 1138 1083
rect 1172 1049 1196 1083
rect 1250 1049 1274 1083
rect 1308 1049 1332 1083
rect 1386 1049 1410 1083
rect 1444 1049 1468 1083
rect 1522 1049 1546 1083
rect 1580 1049 1604 1083
<< psubdiffcont >>
rect 50 27 84 61
rect 186 27 220 61
rect 322 27 356 61
rect 458 27 492 61
rect 594 27 628 61
rect 730 27 764 61
rect 866 27 900 61
rect 1002 27 1036 61
rect 1138 27 1172 61
rect 1274 27 1308 61
rect 1410 27 1444 61
rect 1546 27 1580 61
<< nsubdiffcont >>
rect 50 1049 84 1083
rect 186 1049 220 1083
rect 322 1049 356 1083
rect 458 1049 492 1083
rect 594 1049 628 1083
rect 730 1049 764 1083
rect 866 1049 900 1083
rect 1002 1049 1036 1083
rect 1138 1049 1172 1083
rect 1274 1049 1308 1083
rect 1410 1049 1444 1083
rect 1546 1049 1580 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 356 965 386 991
rect 428 965 458 991
rect 548 965 578 991
rect 620 965 650 991
rect 706 965 736 991
rect 778 965 808 991
rect 898 965 928 991
rect 970 965 1000 991
rect 1056 965 1086 991
rect 1246 965 1276 991
rect 1332 965 1362 991
rect 1522 965 1552 991
rect 1608 965 1638 991
rect 80 351 110 713
rect 166 442 196 713
rect 37 335 110 351
rect 37 301 47 335
rect 81 301 110 335
rect 37 285 110 301
rect 80 199 110 285
rect 152 426 233 442
rect 152 392 189 426
rect 223 392 233 426
rect 152 376 233 392
rect 356 425 386 565
rect 428 534 458 565
rect 428 518 482 534
rect 428 484 438 518
rect 472 484 482 518
rect 428 468 482 484
rect 356 409 410 425
rect 548 423 578 565
rect 620 528 650 565
rect 706 528 736 565
rect 620 518 736 528
rect 620 484 652 518
rect 686 484 736 518
rect 620 474 736 484
rect 778 423 808 565
rect 898 534 928 565
rect 874 518 928 534
rect 874 484 884 518
rect 918 484 928 518
rect 874 468 928 484
rect 152 199 182 376
rect 356 375 366 409
rect 400 375 410 409
rect 356 359 410 375
rect 452 393 904 423
rect 356 243 386 359
rect 452 315 482 393
rect 874 351 904 393
rect 970 419 1000 565
rect 1056 534 1086 565
rect 1056 518 1127 534
rect 1056 504 1083 518
rect 1067 484 1083 504
rect 1117 484 1127 518
rect 1067 468 1127 484
rect 970 403 1024 419
rect 970 369 980 403
rect 1014 369 1024 403
rect 970 353 1024 369
rect 428 285 482 315
rect 524 335 578 351
rect 524 301 534 335
rect 568 301 578 335
rect 524 285 578 301
rect 428 243 458 285
rect 548 243 578 285
rect 620 335 736 345
rect 620 301 652 335
rect 686 301 736 335
rect 620 291 736 301
rect 620 243 650 291
rect 706 243 736 291
rect 778 335 832 351
rect 778 301 788 335
rect 822 301 832 335
rect 778 285 832 301
rect 874 335 928 351
rect 874 301 884 335
rect 918 301 928 335
rect 874 285 928 301
rect 778 243 808 285
rect 898 243 928 285
rect 970 243 1000 353
rect 1067 315 1097 468
rect 1246 351 1276 713
rect 1056 285 1097 315
rect 1193 335 1276 351
rect 1193 301 1203 335
rect 1237 301 1276 335
rect 1193 285 1276 301
rect 1056 243 1086 285
rect 1246 199 1276 285
rect 1332 307 1362 713
rect 1522 549 1552 565
rect 1512 519 1552 549
rect 1512 419 1542 519
rect 1608 460 1638 565
rect 1487 403 1542 419
rect 1487 369 1497 403
rect 1531 369 1542 403
rect 1584 444 1638 460
rect 1584 410 1594 444
rect 1628 410 1638 444
rect 1584 394 1638 410
rect 1487 353 1542 369
rect 1512 308 1542 353
rect 1332 291 1399 307
rect 1332 283 1355 291
rect 1318 257 1355 283
rect 1389 257 1399 291
rect 1512 258 1552 308
rect 1318 221 1399 257
rect 1522 243 1552 258
rect 1608 243 1638 394
rect 1318 199 1348 221
rect 80 89 110 115
rect 152 89 182 115
rect 356 89 386 115
rect 428 89 458 115
rect 548 89 578 115
rect 620 89 650 115
rect 706 89 736 115
rect 778 89 808 115
rect 898 89 928 115
rect 970 89 1000 115
rect 1056 89 1086 115
rect 1246 89 1276 115
rect 1318 89 1348 115
rect 1522 89 1552 115
rect 1608 89 1638 115
<< polycont >>
rect 47 301 81 335
rect 189 392 223 426
rect 438 484 472 518
rect 652 484 686 518
rect 884 484 918 518
rect 366 375 400 409
rect 1083 484 1117 518
rect 980 369 1014 403
rect 534 301 568 335
rect 652 301 686 335
rect 788 301 822 335
rect 884 301 918 335
rect 1203 301 1237 335
rect 1497 369 1531 403
rect 1594 410 1628 444
rect 1355 257 1389 291
<< locali >>
rect 0 1089 1738 1110
rect 0 1049 50 1089
rect 84 1049 186 1089
rect 220 1049 322 1089
rect 356 1049 458 1089
rect 492 1049 594 1089
rect 628 1049 730 1089
rect 764 1049 866 1089
rect 900 1049 1002 1089
rect 1036 1049 1138 1089
rect 1172 1049 1274 1089
rect 1308 1049 1410 1089
rect 1444 1049 1546 1089
rect 1580 1049 1738 1089
rect 35 949 69 1049
rect 35 861 69 877
rect 121 949 155 965
rect 47 335 81 351
rect 47 261 81 301
rect 121 335 155 877
rect 207 949 241 1049
rect 207 861 241 877
rect 311 949 345 1049
rect 311 657 345 673
rect 469 949 537 965
rect 661 949 695 1049
rect 661 657 695 673
rect 819 949 887 965
rect 469 602 537 605
rect 819 602 887 673
rect 121 193 155 301
rect 189 568 537 602
rect 720 568 887 602
rect 1011 949 1045 1049
rect 1011 589 1045 605
rect 1097 949 1131 965
rect 1201 949 1235 1049
rect 1201 861 1235 877
rect 1287 949 1321 965
rect 1097 602 1131 605
rect 1097 568 1187 602
rect 189 426 223 568
rect 438 518 472 534
rect 438 483 472 484
rect 652 518 686 534
rect 472 449 568 483
rect 189 318 223 392
rect 366 409 400 425
rect 366 359 400 375
rect 534 335 568 449
rect 652 335 686 484
rect 189 284 500 318
rect 534 285 568 301
rect 652 285 686 301
rect 720 335 754 568
rect 884 518 918 534
rect 884 483 918 484
rect 466 231 500 284
rect 720 251 754 301
rect 788 449 884 483
rect 1083 518 1117 534
rect 1083 483 1117 484
rect 788 335 822 449
rect 1151 415 1187 568
rect 964 369 980 403
rect 1014 369 1030 403
rect 1097 381 1187 415
rect 1287 403 1321 877
rect 1373 949 1407 1049
rect 1373 861 1407 877
rect 1477 949 1511 965
rect 1477 557 1511 809
rect 1563 949 1597 1049
rect 1563 793 1597 809
rect 1649 949 1683 965
rect 1649 631 1683 809
rect 1682 614 1683 631
rect 1682 597 1706 614
rect 1649 580 1706 597
rect 1477 518 1511 523
rect 1477 484 1628 518
rect 1594 444 1628 484
rect 1097 335 1131 381
rect 1287 369 1497 403
rect 1531 369 1547 403
rect 868 301 884 335
rect 918 301 1131 335
rect 1187 301 1203 335
rect 1237 301 1253 335
rect 788 285 822 301
rect 35 165 155 193
rect 311 215 345 231
rect 69 159 155 165
rect 193 165 227 181
rect 35 115 69 131
rect 193 61 227 131
rect 466 215 537 231
rect 720 217 887 251
rect 466 197 469 215
rect 311 61 345 131
rect 819 215 887 217
rect 469 115 537 131
rect 661 165 695 181
rect 661 61 695 131
rect 819 115 887 131
rect 1011 215 1045 231
rect 1011 61 1045 131
rect 1097 215 1131 301
rect 1287 199 1321 369
rect 1594 335 1628 410
rect 1355 291 1389 307
rect 1477 301 1628 335
rect 1097 115 1131 131
rect 1201 165 1321 199
rect 1359 165 1393 181
rect 1201 115 1235 131
rect 1359 61 1393 131
rect 1477 165 1511 301
rect 1672 268 1706 580
rect 1649 234 1706 268
rect 1477 115 1511 131
rect 1563 165 1597 181
rect 1563 61 1597 131
rect 1649 165 1683 234
rect 1649 115 1683 131
rect 0 21 50 61
rect 84 21 186 61
rect 220 21 322 61
rect 356 21 458 61
rect 492 21 594 61
rect 628 21 730 61
rect 764 21 866 61
rect 900 21 1002 61
rect 1036 21 1138 61
rect 1172 21 1274 61
rect 1308 21 1410 61
rect 1444 21 1546 61
rect 1580 21 1738 61
rect 0 0 1738 21
<< viali >>
rect 50 1083 84 1089
rect 50 1055 84 1083
rect 186 1083 220 1089
rect 186 1055 220 1083
rect 322 1083 356 1089
rect 322 1055 356 1083
rect 458 1083 492 1089
rect 458 1055 492 1083
rect 594 1083 628 1089
rect 594 1055 628 1083
rect 730 1083 764 1089
rect 730 1055 764 1083
rect 866 1083 900 1089
rect 866 1055 900 1083
rect 1002 1083 1036 1089
rect 1002 1055 1036 1083
rect 1138 1083 1172 1089
rect 1138 1055 1172 1083
rect 1274 1083 1308 1089
rect 1274 1055 1308 1083
rect 1410 1083 1444 1089
rect 1410 1055 1444 1083
rect 1546 1083 1580 1089
rect 1546 1055 1580 1083
rect 47 227 81 261
rect 121 301 155 335
rect 438 449 472 483
rect 366 375 400 409
rect 634 301 652 335
rect 652 301 668 335
rect 720 301 754 335
rect 884 449 918 483
rect 1083 449 1117 483
rect 980 369 1014 403
rect 1648 597 1682 631
rect 1477 523 1511 557
rect 1497 369 1531 403
rect 1203 301 1237 335
rect 1355 257 1389 261
rect 1355 227 1389 257
rect 50 27 84 55
rect 50 21 84 27
rect 186 27 220 55
rect 186 21 220 27
rect 322 27 356 55
rect 322 21 356 27
rect 458 27 492 55
rect 458 21 492 27
rect 594 27 628 55
rect 594 21 628 27
rect 730 27 764 55
rect 730 21 764 27
rect 866 27 900 55
rect 866 21 900 27
rect 1002 27 1036 55
rect 1002 21 1036 27
rect 1138 27 1172 55
rect 1138 21 1172 27
rect 1274 27 1308 55
rect 1274 21 1308 27
rect 1410 27 1444 55
rect 1410 21 1444 27
rect 1546 27 1580 55
rect 1546 21 1580 27
<< metal1 >>
rect 0 1089 1738 1110
rect 0 1055 50 1089
rect 84 1055 186 1089
rect 220 1055 322 1089
rect 356 1055 458 1089
rect 492 1055 594 1089
rect 628 1055 730 1089
rect 764 1055 866 1089
rect 900 1055 1002 1089
rect 1036 1055 1138 1089
rect 1172 1055 1274 1089
rect 1308 1055 1410 1089
rect 1444 1055 1546 1089
rect 1580 1055 1738 1089
rect 0 1049 1738 1055
rect 1636 631 1694 637
rect 1614 597 1648 631
rect 1682 597 1694 631
rect 1636 591 1694 597
rect 1465 557 1523 563
rect 1442 523 1477 557
rect 1511 523 1523 557
rect 1465 517 1523 523
rect 426 483 484 489
rect 872 483 930 489
rect 1071 483 1129 489
rect 426 449 438 483
rect 472 449 884 483
rect 918 449 1083 483
rect 1117 449 1129 483
rect 426 443 484 449
rect 872 443 930 449
rect 1071 443 1129 449
rect 354 409 412 415
rect 354 375 366 409
rect 400 375 434 409
rect 968 403 1026 409
rect 1485 403 1543 409
rect 354 369 412 375
rect 968 369 980 403
rect 1014 369 1497 403
rect 1531 369 1543 403
rect 968 363 1026 369
rect 1485 363 1543 369
rect 109 335 167 341
rect 622 335 680 341
rect 109 301 121 335
rect 155 301 634 335
rect 668 301 680 335
rect 109 295 167 301
rect 622 295 680 301
rect 708 335 766 341
rect 1191 335 1249 341
rect 708 301 720 335
rect 754 301 1203 335
rect 1237 301 1249 335
rect 708 295 766 301
rect 1191 295 1249 301
rect 35 261 93 267
rect 1343 261 1401 267
rect 35 227 47 261
rect 81 227 1355 261
rect 1389 227 1401 261
rect 35 221 93 227
rect 1343 221 1401 227
rect 0 55 1738 61
rect 0 21 50 55
rect 84 21 186 55
rect 220 21 322 55
rect 356 21 458 55
rect 492 21 594 55
rect 628 21 730 55
rect 764 21 866 55
rect 900 21 1002 55
rect 1036 21 1138 55
rect 1172 21 1274 55
rect 1308 21 1410 55
rect 1444 21 1546 55
rect 1580 21 1738 55
rect 0 0 1738 21
<< labels >>
rlabel viali 383 392 383 392 1 D
port 1 n
rlabel viali 1100 466 1100 466 1 CK
port 2 n
rlabel viali 1665 614 1665 614 1 Q
port 4 n
rlabel viali 1495 540 1495 540 1 QN
port 3 n
rlabel viali 64 244 64 244 1 SN
rlabel viali 67 48 67 48 1 gnd
rlabel viali 67 1062 67 1062 1 vdd
<< end >>
