* File: sky130_osu_sc_12T_hs__buf_1.pex.spice
* Created: Fri Nov 12 15:08:03 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__BUF_1%GND 1 17 19 26 36 39
r27 36 39 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r28 28 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r29 24 34 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r30 24 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r31 19 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r32 17 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r33 17 28 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r34 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r35 1 26 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_1%VDD 1 13 15 21 25 30 33
r21 30 33 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r22 25 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r23 23 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r24 23 25 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r25 19 28 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r26 19 21 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135 $X2=0.69
+ $Y2=3.635
r27 15 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r28 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r29 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r30 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r31 1 21 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_1%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=2.85
+ $X2=0.635 $Y2=2.85
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2 $X2=0.635
+ $Y2=2.85
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635 $Y=2
+ $X2=0.635 $Y2=2
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=2.165
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=1.835
r45 7 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=2.165
r46 3 11 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=0.475 $Y=0.85
+ $X2=0.475 $Y2=1.835
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_1%A_27_115# 1 3 11 13 15 17 22 26 30 34 38
+ 40 43
r55 39 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.455
+ $X2=0.26 $Y2=1.455
r56 38 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.965 $Y2=1.455
r57 38 39 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.345 $Y2=1.455
r58 34 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r59 32 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.54 $X2=0.26
+ $Y2=1.455
r60 32 34 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=0.26 $Y=1.54
+ $X2=0.26 $Y2=2.955
r61 28 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.37 $X2=0.26
+ $Y2=1.455
r62 28 30 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r63 24 26 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.455
+ $X2=1.18 $Y2=2.455
r64 21 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.455 $X2=0.965 $Y2=1.455
r65 21 22 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.455
+ $X2=1.18 $Y2=1.455
r66 18 21 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.455
+ $X2=0.965 $Y2=1.455
r67 17 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.38
+ $X2=1.18 $Y2=2.455
r68 16 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=1.455
r69 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=2.38
r70 13 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=2.455
r71 13 15 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=3.235
r72 9 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=1.455
r73 9 11 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=0.85
r74 3 36 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r75 3 34 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r76 1 30 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_1%Y 1 3 10 16 26 29 32
r33 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=2.48
r34 24 26 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=1.795
r35 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1
r36 23 26 0.65476 $w=1.7e-07 $l=6.8e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1.795
r37 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r38 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.48
r39 16 19 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.955
r40 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1 $X2=1.12
+ $Y2=1
r41 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.12 $Y=0.755
+ $X2=1.12 $Y2=1
r42 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r43 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r44 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
.ends

