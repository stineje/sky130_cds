* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_15T_ls__aoi22_l
** N=15 EP=0 IP=0 FDC=14
M0 9 A0 gnd gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=400 $Y=575 $D=9
M1 Y A1 9 gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=760 $Y=575 $D=9
M2 10 B0 Y gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=1260 $Y=575 $D=9
M3 gnd B1 10 gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=1620 $Y=575 $D=9
M4 vdd A0 7 vdd phighvt L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=400 $Y=2825 $D=89
M5 7 A1 vdd vdd phighvt L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=830 $Y=2825 $D=89
M6 Y B0 7 vdd phighvt L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=1260 $Y=2825 $D=89
M7 7 B1 Y vdd phighvt L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=1690 $Y=2825 $D=89
X8 gnd vdd Dpar a=6.94725 p=10.61 m=1 $[nwdiode] $X=-45 $Y=2645 $D=185
X9 11 A0 Probe probetype=1 $[A0] $X=383 $Y=3068 $D=289
X10 12 A1 Probe probetype=1 $[A1] $X=723 $Y=2698 $D=289
X11 13 B0 Probe probetype=1 $[B0] $X=1163 $Y=2328 $D=289
X12 14 Y Probe probetype=1 $[Y] $X=1603 $Y=1438 $D=289
X13 15 B1 Probe probetype=1 $[B1] $X=1933 $Y=1963 $D=289
.ENDS
***************************************
