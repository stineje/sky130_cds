* File: sky130_osu_sc_15T_ls__xnor2_l.pex.spice
* Created: Fri Nov 12 15:00:45 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%GND 1 2 33 35 43 45 55 67 69
r70 67 69 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r71 53 55 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.74
r72 46 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r73 41 59 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r74 41 43 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r75 35 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r76 33 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r77 33 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r78 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r79 33 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r80 33 45 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r81 33 46 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r82 33 35 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r83 2 55 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.575 $X2=2.44 $Y2=0.74
r84 1 43 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%VDD 1 2 25 27 34 38 46 54 57 61
c40 34 0 1.59951e-19 $X=0.69 $Y=3.205
r41 57 61 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=2.38 $Y2=5.397
r42 54 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=5.36
+ $X2=2.38 $Y2=5.36
r43 46 49 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.44 $Y=3.205
+ $X2=2.44 $Y2=4.565
r44 44 54 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=5.245
+ $X2=2.44 $Y2=5.397
r45 44 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.44 $Y=5.245
+ $X2=2.44 $Y2=4.565
r46 41 43 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=5.397
+ $X2=1.7 $Y2=5.397
r47 39 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r48 39 41 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r49 38 54 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=5.397
+ $X2=2.44 $Y2=5.397
r50 38 43 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=5.397
+ $X2=1.7 $Y2=5.397
r51 34 37 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r52 32 52 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r53 32 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r54 29 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r55 27 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r56 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r57 25 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r58 25 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r59 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r60 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r61 2 49 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.3
+ $Y=2.825 $X2=2.44 $Y2=4.565
r62 2 46 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.3
+ $Y=2.825 $X2=2.44 $Y2=3.205
r63 1 37 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r64 1 34 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%A 3 5 8 9 13 16 18 19 20 21 22 26 30 37
+ 42 44 45 50 53
r114 47 50 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=0.845 $Y=1.22
+ $X2=0.85 $Y2=1.22
r115 45 50 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=0.99 $Y=1.22
+ $X2=0.85 $Y2=1.22
r116 44 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2 $Y=1.22
+ $X2=2.145 $Y2=1.22
r117 44 45 0.972511 $w=1.7e-07 $l=1.01e-06 $layer=MET1_cond $X=2 $Y=1.22
+ $X2=0.99 $Y2=1.22
r118 39 42 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.145 $Y=2.13
+ $X2=2.225 $Y2=2.13
r119 37 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=1.22
+ $X2=2.145 $Y2=1.22
r120 35 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.045
+ $X2=2.145 $Y2=2.13
r121 35 37 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.145 $Y=2.045
+ $X2=2.145 $Y2=1.22
r122 30 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.845 $Y=1.22
+ $X2=0.845 $Y2=1.22
r123 30 33 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.845 $Y=1.22
+ $X2=0.845 $Y2=1.59
r124 28 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=2.13 $X2=2.225 $Y2=2.13
r125 26 28 73.8383 $w=2.35e-07 $l=3.6e-07 $layer=POLY_cond $X=1.865 $Y=2.145
+ $X2=2.225 $Y2=2.145
r126 24 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.59 $X2=0.845 $Y2=1.59
r127 21 24 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=0.845 $Y=1.465
+ $X2=0.845 $Y2=1.59
r128 21 22 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.465
+ $X2=0.845 $Y2=1.39
r129 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.45 $Y=2.6 $X2=0.45
+ $Y2=2.75
r130 14 26 13.2911 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.865 $Y=2.295
+ $X2=1.865 $Y2=2.145
r131 14 16 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=1.865 $Y=2.295
+ $X2=1.865 $Y2=3.825
r132 13 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=1.39
r133 10 18 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=1.465
+ $X2=0.45 $Y2=1.465
r134 9 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=1.465
+ $X2=0.845 $Y2=1.465
r135 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=1.465
+ $X2=0.55 $Y2=1.465
r136 8 20 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.75
r137 3 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.45 $Y2=1.465
r138 3 5 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.475 $Y2=0.945
r139 1 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=1.54
+ $X2=0.45 $Y2=1.465
r140 1 19 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.425 $Y=1.54
+ $X2=0.425 $Y2=2.6
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%A_27_115# 1 3 11 13 15 17 21 25 29 33
+ 39 41
c78 39 0 1.07013e-19 $X=1.765 $Y=1.59
r79 37 39 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.765 $Y=2.045
+ $X2=1.765 $Y2=1.59
r80 34 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.13
+ $X2=0.26 $Y2=2.13
r81 34 36 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=2.13
+ $X2=0.845 $Y2=2.13
r82 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=2.13
+ $X2=1.765 $Y2=2.045
r83 33 36 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.68 $Y=2.13
+ $X2=0.845 $Y2=2.13
r84 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r85 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.215
+ $X2=0.26 $Y2=2.13
r86 27 29 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=0.26 $Y=2.215
+ $X2=0.26 $Y2=3.205
r87 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.045
+ $X2=0.26 $Y2=2.13
r88 23 25 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=0.26 $Y=2.045
+ $X2=0.26 $Y2=0.865
r89 21 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.59 $X2=1.765 $Y2=1.59
r90 21 22 15.9603 $w=3.02e-07 $l=1e-07 $layer=POLY_cond $X=1.765 $Y=1.59
+ $X2=1.865 $Y2=1.59
r91 17 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.13 $X2=0.845 $Y2=2.13
r92 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=2.13
+ $X2=0.845 $Y2=2.295
r93 13 22 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.425
+ $X2=1.865 $Y2=1.59
r94 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.865 $Y=1.425
+ $X2=1.865 $Y2=0.945
r95 11 19 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.295
r96 3 31 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r97 3 29 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r98 1 25 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%A_238_89# 1 3 11 15 18 21 27 31 35
r60 31 33 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.87 $Y=3.205
+ $X2=2.87 $Y2=4.565
r61 29 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.59 $X2=2.87
+ $Y2=2.505
r62 29 31 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.87 $Y=2.59
+ $X2=2.87 $Y2=3.205
r63 25 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.42 $X2=2.87
+ $Y2=2.505
r64 25 27 101.449 $w=1.68e-07 $l=1.555e-06 $layer=LI1_cond $X=2.87 $Y=2.42
+ $X2=2.87 $Y2=0.865
r65 21 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=2.505
+ $X2=2.87 $Y2=2.505
r66 21 23 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=2.505
+ $X2=1.325 $Y2=2.505
r67 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.505 $X2=1.325 $Y2=2.505
r68 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.505
+ $X2=1.325 $Y2=2.67
r69 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.505
+ $X2=1.325 $Y2=2.34
r70 15 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=1.265 $Y=3.825
+ $X2=1.265 $Y2=2.67
r71 11 19 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=1.265 $Y=0.945
+ $X2=1.265 $Y2=2.34
r72 3 33 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=2.825 $X2=2.87 $Y2=4.565
r73 3 31 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=2.825 $X2=2.87 $Y2=3.205
r74 1 27 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.575 $X2=2.87 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 20 21 23 28
c57 20 0 1.07013e-19 $X=2.655 $Y=1.572
r58 23 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.59
+ $X2=2.53 $Y2=1.59
r59 19 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.59 $X2=2.53 $Y2=1.59
r60 19 20 21.9891 $w=2.74e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=1.572
+ $X2=2.655 $Y2=1.572
r61 14 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=2.75
+ $X2=2.655 $Y2=2.675
r62 14 16 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.655 $Y=2.75
+ $X2=2.655 $Y2=3.825
r63 13 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=2.6
+ $X2=2.655 $Y2=2.675
r64 12 20 16.847 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=2.655 $Y=1.755
+ $X2=2.655 $Y2=1.572
r65 12 13 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=2.655 $Y=1.755
+ $X2=2.655 $Y2=2.6
r66 9 20 16.847 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.655 $Y=1.39
+ $X2=2.655 $Y2=1.572
r67 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.655 $Y=1.39
+ $X2=2.655 $Y2=0.945
r68 7 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=2.675
+ $X2=2.655 $Y2=2.675
r69 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=2.675 $X2=2.3
+ $Y2=2.675
r70 4 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=2.75
+ $X2=2.3 $Y2=2.675
r71 4 6 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.225 $Y=2.75
+ $X2=2.225 $Y2=3.825
r72 1 19 53.6533 $w=2.74e-07 $l=3.85402e-07 $layer=POLY_cond $X=2.225 $Y=1.39
+ $X2=2.53 $Y2=1.572
r73 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.225 $Y=1.39
+ $X2=2.225 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XNOR2_L%Y 1 3 11 15 17 19 24 30 33 36
c56 30 0 1.59951e-19 $X=1.42 $Y=1.875
r57 28 36 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=2.955
+ $X2=1.425 $Y2=3.07
r58 28 30 1.03991 $w=1.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.425 $Y=2.955
+ $X2=1.425 $Y2=1.875
r59 27 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.705
+ $X2=1.425 $Y2=1.59
r60 27 30 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.425 $Y=1.705
+ $X2=1.425 $Y2=1.875
r61 26 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=3.07
+ $X2=1.425 $Y2=3.07
r62 23 24 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.537 $Y=0.985
+ $X2=1.537 $Y2=1.155
r63 19 21 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=1.565 $Y=3.205
+ $X2=1.565 $Y2=4.565
r64 17 26 3.84112 $w=3.85e-07 $l=1.28238e-07 $layer=LI1_cond $X=1.565 $Y=3.185
+ $X2=1.537 $Y2=3.07
r65 17 19 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=1.565 $Y=3.185
+ $X2=1.565 $Y2=3.205
r66 15 23 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.565 $Y=0.865
+ $X2=1.565 $Y2=0.985
r67 11 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=1.59
+ $X2=1.425 $Y2=1.59
r68 11 24 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.425 $Y=1.59
+ $X2=1.425 $Y2=1.155
r69 3 21 240 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.565 $Y2=4.565
r70 3 19 240 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.565 $Y2=3.205
r71 1 15 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.865
.ends

