* File: sky130_osu_sc_18T_ms__tnbufi_1.pex.spice
* Created: Thu Oct 29 17:31:56 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__TNBUFI_1%GND 1 12 14 21 26 29
r34 26 29 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r35 23 24 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r36 19 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r37 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r38 14 24 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r39 12 23 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r40 12 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r41 12 14 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r42 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TNBUFI_1%VDD 1 10 12 18 25 28 32
r19 28 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r20 25 28 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r21 22 32 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507 $X2=1.02
+ $Y2=6.507
r22 22 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r23 18 21 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.69 $Y=3.795
+ $X2=0.69 $Y2=5.835
r24 16 23 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r25 16 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r26 12 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r27 12 14 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r28 10 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r29 10 14 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r30 1 21 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r31 1 18 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TNBUFI_1%A_27_115# 1 2 9 13 17 21 23 26 31
r44 27 31 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=2.175
+ $X2=0.905 $Y2=2.175
r45 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.175 $X2=0.69 $Y2=2.175
r46 22 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.175
+ $X2=0.26 $Y2=2.175
r47 21 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=2.175
+ $X2=0.69 $Y2=2.175
r48 21 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=2.175
+ $X2=0.345 $Y2=2.175
r49 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r50 15 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.26 $X2=0.26
+ $Y2=2.175
r51 15 17 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=0.26 $Y=2.26
+ $X2=0.26 $Y2=3.455
r52 11 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.09 $X2=0.26
+ $Y2=2.175
r53 11 13 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=0.26 $Y=2.09
+ $X2=0.26 $Y2=0.825
r54 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.01
+ $X2=0.905 $Y2=2.175
r55 7 9 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.905 $Y=2.01
+ $X2=0.905 $Y2=1.075
r56 2 19 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r57 2 17 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r58 1 13 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TNBUFI_1%OE 3 5 6 8 11 14 17 22
r42 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.765 $X2=0.69 $Y2=2.765
r43 19 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=2.765
r44 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=2.96
r45 12 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.725
+ $X2=0.475 $Y2=1.725
r46 6 23 49.2914 $w=4.58e-07 $l=4.23124e-07 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.587 $Y2=2.765
r47 6 11 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=4.585
r48 6 8 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.475 $Y2=4.585
r49 3 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.475 $Y2=1.725
r50 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.475 $Y2=1.075
r51 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=1.8 $X2=0.27
+ $Y2=1.725
r52 1 6 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.8 $X2=0.27
+ $Y2=2.86
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TNBUFI_1%A 3 7 13 14 17 19
r47 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=3.33
+ $X2=1.14 $Y2=3.33
r48 14 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.09
+ $X2=1.325 $Y2=2.255
r49 14 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.09
+ $X2=1.325 $Y2=1.925
r50 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.09 $X2=1.325 $Y2=2.09
r51 10 19 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=2.175
+ $X2=1.14 $Y2=3.33
r52 9 13 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=2.09
+ $X2=1.325 $Y2=2.09
r53 9 10 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.09 $X2=1.14
+ $Y2=2.175
r54 7 23 1194.74 $w=1.5e-07 $l=2.33e-06 $layer=POLY_cond $X=1.265 $Y=4.585
+ $X2=1.265 $Y2=2.255
r55 3 22 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.265 $Y=1.075
+ $X2=1.265 $Y2=1.925
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TNBUFI_1%Y 1 2 10 13 17 18 21
r32 28 30 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.48 $Y=3.455
+ $X2=1.48 $Y2=5.835
r33 18 28 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.48 $Y=2.59
+ $X2=1.48 $Y2=3.455
r34 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.59
+ $X2=1.48 $Y2=2.59
r35 14 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.48 $Y=1.48
+ $X2=1.48 $Y2=0.825
r36 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.48
+ $X2=1.48 $Y2=1.48
r37 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.475
+ $X2=1.48 $Y2=2.59
r38 8 10 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.475
+ $X2=1.48 $Y2=1.82
r39 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.595
+ $X2=1.48 $Y2=1.48
r40 7 10 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.595
+ $X2=1.48 $Y2=1.82
r41 2 30 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.48 $Y2=5.835
r42 2 28 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.48 $Y2=3.455
r43 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.825
.ends

