* File: sky130_osu_sc_12T_hs__inv_l.pex.spice
* Created: Fri Nov 12 15:11:27 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__INV_L%GND 1 11 15 24 27
r14 24 27 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=0.19
+ $X2=0.495 $Y2=0.24
r15 13 15 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r16 11 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r17 11 13 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r18 1 15 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__INV_L%VDD 1 9 13 18 21
r12 21 24 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=4.19
+ $X2=0.495 $Y2=4.24
r13 18 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=4.24
+ $X2=0.34 $Y2=4.24
r14 11 18 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.125
+ $X2=0.172 $Y2=4.277
r15 11 13 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=4.125
+ $X2=0.26 $Y2=3.605
r16 9 18 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.125 $X2=0.34 $Y2=4.21
r17 1 13 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.015 $X2=0.26 $Y2=3.605
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__INV_L%A 3 7 10 15 17 19 22
r37 17 19 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=1.825
+ $X2=0.535 $Y2=1.825
r38 15 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r39 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.405 $Y2=1.825
r40 13 15 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.32 $Y2=2.85
r41 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.825 $X2=0.535 $Y2=1.825
r42 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.99
r43 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.66
r44 7 12 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=0.475 $Y=3.435
+ $X2=0.475 $Y2=1.99
r45 3 11 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.475 $Y=0.785
+ $X2=0.475 $Y2=1.66
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__INV_L%Y 1 3 10 16 24 27 30
r31 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.48
r32 22 24 0.616245 $w=1.7e-07 $l=6.4e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=1.725
r33 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.485
+ $X2=0.69 $Y2=1.37
r34 21 24 0.231092 $w=1.7e-07 $l=2.4e-07 $layer=MET1_cond $X=0.69 $Y=1.485
+ $X2=0.69 $Y2=1.725
r35 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r36 16 19 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=3.605
r37 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.37
+ $X2=0.69 $Y2=1.37
r38 10 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.69 $Y=0.74
+ $X2=0.69 $Y2=1.37
r39 3 19 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.015 $X2=0.69 $Y2=3.605
r40 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

