* File: sky130_osu_sc_18T_ls__buf_2.pxi.spice
* Created: Fri Nov 12 14:14:47 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__BUF_2%GND N_GND_M1003_d N_GND_M1001_s N_GND_M1003_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p N_GND_c_15_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_LS__BUF_2%GND
x_PM_SKY130_OSU_SC_18T_LS__BUF_2%VDD N_VDD_M1002_d N_VDD_M1005_d N_VDD_M1002_b
+ N_VDD_c_36_p N_VDD_c_37_p N_VDD_c_46_p N_VDD_c_51_p VDD N_VDD_c_38_p
+ PM_SKY130_OSU_SC_18T_LS__BUF_2%VDD
x_PM_SKY130_OSU_SC_18T_LS__BUF_2%A N_A_M1003_g N_A_M1002_g N_A_c_66_n N_A_c_67_n
+ A PM_SKY130_OSU_SC_18T_LS__BUF_2%A
x_PM_SKY130_OSU_SC_18T_LS__BUF_2%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1002_s N_A_27_115#_M1000_g N_A_27_115#_c_120_n
+ N_A_27_115#_M1004_g N_A_27_115#_c_105_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_124_n N_A_27_115#_M1005_g N_A_27_115#_c_110_n
+ N_A_27_115#_c_111_n N_A_27_115#_c_112_n N_A_27_115#_c_115_n
+ N_A_27_115#_c_116_n N_A_27_115#_c_118_n N_A_27_115#_c_119_n
+ PM_SKY130_OSU_SC_18T_LS__BUF_2%A_27_115#
x_PM_SKY130_OSU_SC_18T_LS__BUF_2%Y N_Y_M1000_d N_Y_M1004_s N_Y_c_170_n
+ N_Y_c_178_n Y N_Y_c_174_n N_Y_c_177_n PM_SKY130_OSU_SC_18T_LS__BUF_2%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1003_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1003_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_A_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.075
cc_5 N_GND_M1003_b N_A_M1002_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_6 N_GND_M1003_b N_A_c_66_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_7 N_GND_M1003_b N_A_c_67_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_8 N_GND_M1003_b N_A_27_115#_M1000_g 0.0207501f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=1.075
cc_9 N_GND_c_3_p N_A_27_115#_M1000_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=1.075
cc_10 N_GND_c_10_p N_A_27_115#_M1000_g 0.00606474f $X=1.465 $Y=0.152 $X2=0.905
+ $Y2=1.075
cc_11 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=1.075
cc_12 N_GND_M1003_b N_A_27_115#_c_105_n 0.0597491f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.86
cc_13 N_GND_M1003_b N_A_27_115#_M1001_g 0.0264941f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_14 N_GND_c_10_p N_A_27_115#_M1001_g 0.00606474f $X=1.465 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_15 N_GND_c_15_p N_A_27_115#_M1001_g 0.00713292f $X=1.55 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_16 N_GND_c_4_p N_A_27_115#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_M1003_b N_A_27_115#_c_110_n 0.0268682f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=2.935
cc_18 N_GND_M1003_b N_A_27_115#_c_111_n 0.0617719f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=1.935
cc_19 N_GND_M1003_b N_A_27_115#_c_112_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_20 N_GND_c_2_p N_A_27_115#_c_112_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_21 N_GND_c_4_p N_A_27_115#_c_112_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_22 N_GND_M1003_b N_A_27_115#_c_115_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.455
cc_23 N_GND_M1003_b N_A_27_115#_c_116_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.935
cc_24 N_GND_c_3_p N_A_27_115#_c_116_n 0.00702738f $X=0.69 $Y=0.825 $X2=0.88
+ $Y2=1.935
cc_25 N_GND_M1003_b N_A_27_115#_c_118_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.935
cc_26 N_GND_M1003_b N_A_27_115#_c_119_n 0.00592383f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.935
cc_27 N_GND_M1003_b N_Y_c_170_n 0.00155118f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.825
cc_28 N_GND_c_10_p N_Y_c_170_n 0.00734006f $X=1.465 $Y=0.152 $X2=1.12 $Y2=0.825
cc_29 N_GND_c_4_p N_Y_c_170_n 0.00475776f $X=1.02 $Y=0.19 $X2=1.12 $Y2=0.825
cc_30 N_GND_M1003_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=2.27
cc_31 N_GND_M1003_b N_Y_c_174_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.48
cc_32 N_GND_c_3_p N_Y_c_174_n 0.00125659f $X=0.69 $Y=0.825 $X2=1.12 $Y2=1.48
cc_33 N_GND_c_15_p N_Y_c_174_n 0.00125659f $X=1.55 $Y=0.825 $X2=1.12 $Y2=1.48
cc_34 N_GND_M1003_b N_Y_c_177_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.96
cc_35 N_VDD_M1002_b N_A_M1002_g 0.0245629f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_36 N_VDD_c_36_p N_A_M1002_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475 $Y2=4.585
cc_37 N_VDD_c_37_p N_A_M1002_g 0.00354579f $X=0.69 $Y=4.135 $X2=0.475 $Y2=4.585
cc_38 N_VDD_c_38_p N_A_M1002_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=4.585
cc_39 N_VDD_M1002_d N_A_c_67_n 0.00628533f $X=0.55 $Y=3.085 $X2=0.635 $Y2=2.48
cc_40 N_VDD_M1002_b N_A_c_67_n 0.00328912f $X=-0.045 $Y=2.905 $X2=0.635 $Y2=2.48
cc_41 N_VDD_c_37_p N_A_c_67_n 0.00264661f $X=0.69 $Y=4.135 $X2=0.635 $Y2=2.48
cc_42 N_VDD_M1002_d A 0.00797576f $X=0.55 $Y=3.085 $X2=0.635 $Y2=3.33
cc_43 N_VDD_c_37_p A 0.00510982f $X=0.69 $Y=4.135 $X2=0.635 $Y2=3.33
cc_44 N_VDD_M1002_b N_A_27_115#_c_120_n 0.014249f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=3.01
cc_45 N_VDD_c_37_p N_A_27_115#_c_120_n 0.00354579f $X=0.69 $Y=4.135 $X2=0.905
+ $Y2=3.01
cc_46 N_VDD_c_46_p N_A_27_115#_c_120_n 0.00606474f $X=1.465 $Y=6.507 $X2=0.905
+ $Y2=3.01
cc_47 N_VDD_c_38_p N_A_27_115#_c_120_n 0.00468827f $X=1.02 $Y=6.47 $X2=0.905
+ $Y2=3.01
cc_48 N_VDD_M1002_b N_A_27_115#_c_124_n 0.0169732f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=3.01
cc_49 N_VDD_c_37_p N_A_27_115#_c_124_n 3.67508e-19 $X=0.69 $Y=4.135 $X2=1.335
+ $Y2=3.01
cc_50 N_VDD_c_46_p N_A_27_115#_c_124_n 0.00610567f $X=1.465 $Y=6.507 $X2=1.335
+ $Y2=3.01
cc_51 N_VDD_c_51_p N_A_27_115#_c_124_n 0.00732698f $X=1.55 $Y=3.455 $X2=1.335
+ $Y2=3.01
cc_52 N_VDD_c_38_p N_A_27_115#_c_124_n 0.00470215f $X=1.02 $Y=6.47 $X2=1.335
+ $Y2=3.01
cc_53 N_VDD_M1002_b N_A_27_115#_c_110_n 0.0170554f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.935
cc_54 N_VDD_M1002_b N_A_27_115#_c_115_n 0.00996008f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.455
cc_55 N_VDD_c_36_p N_A_27_115#_c_115_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=3.455
cc_56 N_VDD_c_38_p N_A_27_115#_c_115_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26
+ $Y2=3.455
cc_57 N_VDD_M1002_b N_Y_c_178_n 0.00290209f $X=-0.045 $Y=2.905 $X2=1.12 $Y2=2.96
cc_58 N_VDD_c_46_p N_Y_c_178_n 0.00734006f $X=1.465 $Y=6.507 $X2=1.12 $Y2=2.96
cc_59 N_VDD_c_38_p N_Y_c_178_n 0.00475776f $X=1.02 $Y=6.47 $X2=1.12 $Y2=2.96
cc_60 N_VDD_M1002_b N_Y_c_177_n 0.00409378f $X=-0.045 $Y=2.905 $X2=1.12 $Y2=2.96
cc_61 A N_A_27_115#_M1002_s 0.00414531f $X=0.635 $Y=3.33 $X2=0.135 $Y2=3.085
cc_62 N_A_M1003_g N_A_27_115#_M1000_g 0.0386421f $X=0.475 $Y=1.075 $X2=0.905
+ $Y2=1.075
cc_63 A N_A_27_115#_c_120_n 0.00419145f $X=0.635 $Y=3.33 $X2=0.905 $Y2=3.01
cc_64 N_A_M1003_g N_A_27_115#_c_105_n 0.00260138f $X=0.475 $Y=1.075 $X2=1.18
+ $Y2=2.86
cc_65 N_A_M1002_g N_A_27_115#_c_105_n 0.00209773f $X=0.475 $Y=4.585 $X2=1.18
+ $Y2=2.86
cc_66 N_A_c_66_n N_A_27_115#_c_105_n 0.0139096f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_67 N_A_c_67_n N_A_27_115#_c_105_n 0.00361737f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_68 N_A_M1002_g N_A_27_115#_c_110_n 0.049829f $X=0.475 $Y=4.585 $X2=1.335
+ $Y2=2.935
cc_69 N_A_c_67_n N_A_27_115#_c_110_n 0.00473532f $X=0.635 $Y=2.48 $X2=1.335
+ $Y2=2.935
cc_70 N_A_M1003_g N_A_27_115#_c_112_n 0.0148408f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_71 N_A_M1003_g N_A_27_115#_c_115_n 0.0337582f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=3.455
cc_72 N_A_c_67_n N_A_27_115#_c_115_n 0.0548951f $X=0.635 $Y=2.48 $X2=0.26
+ $Y2=3.455
cc_73 A N_A_27_115#_c_115_n 0.0155137f $X=0.635 $Y=3.33 $X2=0.26 $Y2=3.455
cc_74 N_A_M1003_g N_A_27_115#_c_116_n 0.0207696f $X=0.475 $Y=1.075 $X2=0.88
+ $Y2=1.935
cc_75 N_A_c_66_n N_A_27_115#_c_116_n 0.00273049f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_76 N_A_c_67_n N_A_27_115#_c_116_n 0.00886797f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_77 N_A_M1003_g N_A_27_115#_c_119_n 6.59135e-19 $X=0.475 $Y=1.075 $X2=0.965
+ $Y2=1.935
cc_78 N_A_c_67_n N_Y_c_178_n 0.0135622f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_79 A N_Y_c_178_n 0.00731851f $X=0.635 $Y=3.33 $X2=1.12 $Y2=2.96
cc_80 N_A_M1003_g Y 0.00310306f $X=0.475 $Y=1.075 $X2=1.055 $Y2=2.27
cc_81 N_A_c_66_n Y 0.00441844f $X=0.635 $Y=2.48 $X2=1.055 $Y2=2.27
cc_82 N_A_c_67_n Y 0.0200396f $X=0.635 $Y=2.48 $X2=1.055 $Y2=2.27
cc_83 N_A_M1003_g N_Y_c_174_n 7.99941e-19 $X=0.475 $Y=1.075 $X2=1.12 $Y2=1.48
cc_84 N_A_c_67_n N_Y_c_177_n 0.00609526f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_85 N_A_27_115#_M1000_g N_Y_c_170_n 0.00231637f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_86 N_A_27_115#_M1001_g N_Y_c_170_n 0.00231637f $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_87 N_A_27_115#_c_111_n N_Y_c_170_n 0.0030245f $X=1.18 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_88 N_A_27_115#_c_119_n N_Y_c_170_n 7.32051e-19 $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_89 N_A_27_115#_c_120_n N_Y_c_178_n 0.00155107f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_90 N_A_27_115#_c_124_n N_Y_c_178_n 0.00250481f $X=1.335 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_91 N_A_27_115#_c_110_n N_Y_c_178_n 0.0121869f $X=1.335 $Y=2.935 $X2=1.12
+ $Y2=2.96
cc_92 N_A_27_115#_M1000_g Y 0.00251111f $X=0.905 $Y=1.075 $X2=1.055 $Y2=2.27
cc_93 N_A_27_115#_c_105_n Y 0.0310322f $X=1.18 $Y=2.86 $X2=1.055 $Y2=2.27
cc_94 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.055 $Y2=2.27
cc_95 N_A_27_115#_c_111_n Y 0.0153085f $X=1.18 $Y=1.935 $X2=1.055 $Y2=2.27
cc_96 N_A_27_115#_c_116_n Y 8.73078e-19 $X=0.88 $Y=1.935 $X2=1.055 $Y2=2.27
cc_97 N_A_27_115#_c_119_n Y 0.0121742f $X=0.965 $Y=1.935 $X2=1.055 $Y2=2.27
cc_98 N_A_27_115#_M1000_g N_Y_c_174_n 0.00526938f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=1.48
cc_99 N_A_27_115#_M1001_g N_Y_c_174_n 0.00908199f $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=1.48
cc_100 N_A_27_115#_c_119_n N_Y_c_174_n 0.00278861f $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=1.48
cc_101 N_A_27_115#_c_120_n N_Y_c_177_n 0.0011906f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_102 N_A_27_115#_c_105_n N_Y_c_177_n 0.00226191f $X=1.18 $Y=2.86 $X2=1.12
+ $Y2=2.96
cc_103 N_A_27_115#_c_124_n N_Y_c_177_n 0.00303932f $X=1.335 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_104 N_A_27_115#_c_110_n N_Y_c_177_n 0.00877967f $X=1.335 $Y=2.935 $X2=1.12
+ $Y2=2.96
