* File: sky130_osu_sc_18T_hs__and2_l.pxi.spice
* Created: Fri Nov 12 13:47:11 2021
* 
x_PM_SKY130_OSU_SC_18T_HS__AND2_L%GND N_GND_M1001_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_8_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_HS__AND2_L%GND
x_PM_SKY130_OSU_SC_18T_HS__AND2_L%VDD N_VDD_M1005_s N_VDD_M1003_d N_VDD_M1005_b
+ N_VDD_c_35_p N_VDD_c_36_p N_VDD_c_43_p N_VDD_c_49_p VDD N_VDD_c_37_p
+ PM_SKY130_OSU_SC_18T_HS__AND2_L%VDD
x_PM_SKY130_OSU_SC_18T_HS__AND2_L%A N_A_M1002_g N_A_M1005_g N_A_c_62_n
+ N_A_c_63_n A PM_SKY130_OSU_SC_18T_HS__AND2_L%A
x_PM_SKY130_OSU_SC_18T_HS__AND2_L%B N_B_M1001_g N_B_M1003_g N_B_c_92_n
+ N_B_c_93_n B PM_SKY130_OSU_SC_18T_HS__AND2_L%B
x_PM_SKY130_OSU_SC_18T_HS__AND2_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1005_d N_A_27_115#_M1000_g N_A_27_115#_M1004_g
+ N_A_27_115#_c_129_n N_A_27_115#_c_130_n N_A_27_115#_c_131_n
+ N_A_27_115#_c_132_n N_A_27_115#_c_135_n N_A_27_115#_c_136_n
+ N_A_27_115#_c_145_n N_A_27_115#_c_137_n N_A_27_115#_c_138_n
+ N_A_27_115#_c_139_n N_A_27_115#_c_161_n
+ PM_SKY130_OSU_SC_18T_HS__AND2_L%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__AND2_L%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_194_n
+ N_Y_c_196_n Y N_Y_c_198_n N_Y_c_199_n PM_SKY130_OSU_SC_18T_HS__AND2_L%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.0945332f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1002_b N_A_c_62_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_5 N_GND_M1002_b N_A_c_63_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.765
cc_6 N_GND_M1002_b N_B_M1001_g 0.0600862f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_7 N_GND_c_2_p N_B_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.945
cc_8 N_GND_c_8_p N_B_M1001_g 0.00376152f $X=1.05 $Y=0.825 $X2=0.835 $Y2=0.945
cc_9 N_GND_c_3_p N_B_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.945
cc_10 N_GND_M1002_b N_B_M1003_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=5.085
cc_11 N_GND_M1002_b N_B_c_92_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_12 N_GND_M1002_b N_B_c_93_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_13 N_GND_M1002_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.96
cc_14 N_GND_M1002_b N_A_27_115#_M1000_g 0.0525555f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.945
cc_15 N_GND_c_8_p N_A_27_115#_M1000_g 0.00733906f $X=1.05 $Y=0.825 $X2=1.335
+ $Y2=0.945
cc_16 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=0.945
cc_17 N_GND_M1002_b N_A_27_115#_c_129_n 0.0373102f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.1
cc_18 N_GND_M1002_b N_A_27_115#_c_130_n 0.0470206f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.81
cc_19 N_GND_M1002_b N_A_27_115#_c_131_n 0.0076653f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.96
cc_20 N_GND_M1002_b N_A_27_115#_c_132_n 0.0272477f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_21 N_GND_c_2_p N_A_27_115#_c_132_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_22 N_GND_c_3_p N_A_27_115#_c_132_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_23 N_GND_M1002_b N_A_27_115#_c_135_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.935
cc_24 N_GND_M1002_b N_A_27_115#_c_136_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.935
cc_25 N_GND_M1002_b N_A_27_115#_c_137_n 0.0275781f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_26 N_GND_M1002_b N_A_27_115#_c_138_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.935
cc_27 N_GND_M1002_b N_A_27_115#_c_139_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=4.225
cc_28 N_GND_M1002_b N_Y_c_194_n 0.0191683f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_29 N_GND_c_3_p N_Y_c_194_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.825
cc_30 N_GND_M1002_b N_Y_c_196_n 0.0163869f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_31 N_GND_M1002_b Y 0.0401139f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_32 N_GND_M1002_b N_Y_c_198_n 0.0157042f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.48
cc_33 N_GND_M1002_b N_Y_c_199_n 0.0141689f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_34 N_VDD_M1005_b N_A_M1005_g 0.0888934f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_35 N_VDD_c_35_p N_A_M1005_g 0.00713292f $X=0.26 $Y=4.475 $X2=0.475 $Y2=5.085
cc_36 N_VDD_c_36_p N_A_M1005_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=5.085
cc_37 N_VDD_c_37_p N_A_M1005_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=5.085
cc_38 N_VDD_M1005_b N_A_c_62_n 0.0111025f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=2.765
cc_39 N_VDD_M1005_b N_A_c_63_n 0.0185679f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.765
cc_40 N_VDD_M1005_b A 0.0210226f $X=-0.045 $Y=2.905 $X2=0.275 $Y2=3.33
cc_41 N_VDD_M1005_b N_B_M1003_g 0.0726621f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=5.085
cc_42 N_VDD_c_36_p N_B_M1003_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=5.085
cc_43 N_VDD_c_43_p N_B_M1003_g 0.00354579f $X=1.12 $Y=4.475 $X2=0.905 $Y2=5.085
cc_44 N_VDD_c_37_p N_B_M1003_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.905 $Y2=5.085
cc_45 N_VDD_M1005_b N_B_c_93_n 0.00170274f $X=-0.045 $Y=2.905 $X2=0.95 $Y2=2.425
cc_46 N_VDD_M1005_b B 0.012052f $X=-0.045 $Y=2.905 $X2=0.955 $Y2=2.96
cc_47 N_VDD_M1005_b N_A_27_115#_M1004_g 0.077807f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=5.085
cc_48 N_VDD_c_43_p N_A_27_115#_M1004_g 0.00354579f $X=1.12 $Y=4.475 $X2=1.335
+ $Y2=5.085
cc_49 N_VDD_c_49_p N_A_27_115#_M1004_g 0.00606474f $X=1.12 $Y=6.507 $X2=1.335
+ $Y2=5.085
cc_50 N_VDD_c_37_p N_A_27_115#_M1004_g 0.00468827f $X=1.02 $Y=6.47 $X2=1.335
+ $Y2=5.085
cc_51 N_VDD_M1005_b N_A_27_115#_c_131_n 0.00525234f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.96
cc_52 N_VDD_M1005_b N_A_27_115#_c_145_n 0.00155118f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=4.475
cc_53 N_VDD_c_36_p N_A_27_115#_c_145_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69
+ $Y2=4.475
cc_54 N_VDD_c_37_p N_A_27_115#_c_145_n 0.00475776f $X=1.02 $Y=6.47 $X2=0.69
+ $Y2=4.475
cc_55 N_VDD_M1005_b N_A_27_115#_c_139_n 0.0102128f $X=-0.045 $Y=2.905 $X2=0.65
+ $Y2=4.225
cc_56 N_VDD_M1005_b N_Y_c_196_n 0.0596585f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.59
cc_57 N_VDD_c_49_p N_Y_c_196_n 0.00757793f $X=1.12 $Y=6.507 $X2=1.55 $Y2=2.59
cc_58 N_VDD_c_37_p N_Y_c_196_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.55 $Y2=2.59
cc_59 N_A_M1002_g N_B_M1001_g 0.130464f $X=0.475 $Y=0.945 $X2=0.835 $Y2=0.945
cc_60 N_A_M1002_g N_B_M1003_g 0.0772393f $X=0.475 $Y=0.945 $X2=0.905 $Y2=5.085
cc_61 N_A_M1002_g N_B_c_93_n 7.8234e-19 $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.425
cc_62 N_A_M1002_g N_A_27_115#_c_132_n 0.0274292f $X=0.475 $Y=0.945 $X2=0.26
+ $Y2=0.825
cc_63 N_A_M1002_g N_A_27_115#_c_135_n 0.0160984f $X=0.475 $Y=0.945 $X2=0.525
+ $Y2=1.935
cc_64 N_A_c_62_n N_A_27_115#_c_135_n 0.00117122f $X=0.475 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_65 N_A_c_63_n N_A_27_115#_c_135_n 2.65873e-19 $X=0.27 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_66 N_A_c_62_n N_A_27_115#_c_136_n 0.00133457f $X=0.475 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_67 N_A_c_63_n N_A_27_115#_c_136_n 0.0055861f $X=0.27 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_68 N_A_M1002_g N_A_27_115#_c_138_n 0.00322084f $X=0.475 $Y=0.945 $X2=0.61
+ $Y2=1.935
cc_69 N_A_M1002_g N_A_27_115#_c_139_n 0.0265302f $X=0.475 $Y=0.945 $X2=0.65
+ $Y2=4.225
cc_70 N_A_M1005_g N_A_27_115#_c_139_n 0.0464097f $X=0.475 $Y=5.085 $X2=0.65
+ $Y2=4.225
cc_71 N_A_c_62_n N_A_27_115#_c_139_n 0.00766302f $X=0.475 $Y=2.765 $X2=0.65
+ $Y2=4.225
cc_72 N_A_c_63_n N_A_27_115#_c_139_n 0.0541092f $X=0.27 $Y=2.765 $X2=0.65
+ $Y2=4.225
cc_73 A N_A_27_115#_c_139_n 0.00758489f $X=0.275 $Y=3.33 $X2=0.65 $Y2=4.225
cc_74 N_A_M1005_g N_A_27_115#_c_161_n 0.00355211f $X=0.475 $Y=5.085 $X2=0.65
+ $Y2=4.395
cc_75 N_B_M1001_g N_A_27_115#_M1000_g 0.0429232f $X=0.835 $Y=0.945 $X2=1.335
+ $Y2=0.945
cc_76 N_B_M1001_g N_A_27_115#_c_129_n 0.0104742f $X=0.835 $Y=0.945 $X2=1.37
+ $Y2=2.1
cc_77 N_B_M1003_g N_A_27_115#_c_130_n 0.00773101f $X=0.905 $Y=5.085 $X2=1.352
+ $Y2=2.81
cc_78 N_B_c_92_n N_A_27_115#_c_130_n 0.0206104f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.81
cc_79 N_B_c_93_n N_A_27_115#_c_130_n 0.0033451f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.81
cc_80 N_B_M1003_g N_A_27_115#_c_131_n 0.0684885f $X=0.905 $Y=5.085 $X2=1.352
+ $Y2=2.96
cc_81 N_B_c_93_n N_A_27_115#_c_131_n 0.00156524f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.96
cc_82 B N_A_27_115#_c_131_n 0.0037561f $X=0.955 $Y=2.96 $X2=1.352 $Y2=2.96
cc_83 N_B_M1001_g N_A_27_115#_c_137_n 0.0182215f $X=0.835 $Y=0.945 $X2=1.43
+ $Y2=1.935
cc_84 N_B_c_92_n N_A_27_115#_c_137_n 0.00258465f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_85 N_B_c_93_n N_A_27_115#_c_137_n 0.0101796f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_86 N_B_M1001_g N_A_27_115#_c_139_n 0.00755919f $X=0.835 $Y=0.945 $X2=0.65
+ $Y2=4.225
cc_87 N_B_M1003_g N_A_27_115#_c_139_n 0.0279997f $X=0.905 $Y=5.085 $X2=0.65
+ $Y2=4.225
cc_88 N_B_c_93_n N_A_27_115#_c_139_n 0.0541375f $X=0.95 $Y=2.425 $X2=0.65
+ $Y2=4.225
cc_89 B N_A_27_115#_c_139_n 0.00866797f $X=0.955 $Y=2.96 $X2=0.65 $Y2=4.225
cc_90 N_B_c_93_n N_Y_c_196_n 0.0153635f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_91 B N_Y_c_196_n 0.00659455f $X=0.955 $Y=2.96 $X2=1.55 $Y2=2.59
cc_92 N_B_M1001_g Y 6.71108e-19 $X=0.835 $Y=0.945 $X2=1.555 $Y2=2.22
cc_93 N_B_c_93_n Y 0.00695761f $X=0.95 $Y=2.425 $X2=1.555 $Y2=2.22
cc_94 N_B_M1001_g N_Y_c_198_n 0.00101796f $X=0.835 $Y=0.945 $X2=1.55 $Y2=1.48
cc_95 N_B_c_92_n N_Y_c_199_n 5.70769e-19 $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_96 N_B_c_93_n N_Y_c_199_n 0.00532157f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_97 N_A_27_115#_M1000_g N_Y_c_194_n 0.0152627f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=0.825
cc_98 N_A_27_115#_c_129_n N_Y_c_194_n 0.00168f $X=1.37 $Y=2.1 $X2=1.55 $Y2=0.825
cc_99 N_A_27_115#_c_137_n N_Y_c_194_n 0.00530006f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_100 N_A_27_115#_M1004_g N_Y_c_196_n 0.0472737f $X=1.335 $Y=5.085 $X2=1.55
+ $Y2=2.59
cc_101 N_A_27_115#_c_129_n N_Y_c_196_n 0.00125776f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_102 N_A_27_115#_c_130_n N_Y_c_196_n 0.0115869f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_103 N_A_27_115#_c_137_n N_Y_c_196_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_104 N_A_27_115#_M1000_g Y 0.00406656f $X=1.335 $Y=0.945 $X2=1.555 $Y2=2.22
cc_105 N_A_27_115#_c_129_n Y 0.00711756f $X=1.37 $Y=2.1 $X2=1.555 $Y2=2.22
cc_106 N_A_27_115#_c_130_n Y 0.00892438f $X=1.352 $Y=2.81 $X2=1.555 $Y2=2.22
cc_107 N_A_27_115#_c_137_n Y 0.0152626f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_108 N_A_27_115#_M1000_g N_Y_c_198_n 0.00725105f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=1.48
cc_109 N_A_27_115#_c_129_n N_Y_c_198_n 0.00154864f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=1.48
cc_110 N_A_27_115#_c_137_n N_Y_c_198_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.48
cc_111 N_A_27_115#_c_129_n N_Y_c_199_n 4.58687e-19 $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_112 N_A_27_115#_c_130_n N_Y_c_199_n 0.00721849f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_113 N_A_27_115#_c_137_n N_Y_c_199_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
