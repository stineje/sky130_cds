* File: sky130_osu_sc_18T_ms__and2_2.pex.spice
* Created: Thu Oct 29 17:27:21 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__AND2_2%GND 1 2 19 23 27 30 34 39 41
r44 39 41 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r45 25 34 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.895 $Y2=0.152
r46 25 27 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r47 21 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r48 19 34 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r49 19 29 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r50 19 30 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r51 19 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.17 $X2=1.7
+ $Y2=0.17
r52 19 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r53 19 21 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r54 19 30 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r55 19 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r56 2 27 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r57 1 23 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_2%VDD 1 2 3 19 23 27 33 39 45 47 52
r36 52 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.49 $X2=1.7
+ $Y2=6.49
r37 47 52 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r38 47 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r39 45 56 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r40 43 56 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r41 43 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r42 39 42 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r43 37 45 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.895 $Y2=6.507
r44 37 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r45 33 36 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r46 31 44 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r47 31 36 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r48 28 50 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r49 28 30 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r50 27 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r51 27 30 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r52 23 26 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r53 21 50 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r54 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r55 19 50 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r56 19 56 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r57 19 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r58 3 42 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r59 3 39 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r60 2 36 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r61 2 33 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r62 1 26 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r63 1 23 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_2%A 3 7 12 15 18
r32 16 18 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.765
+ $X2=0.475 $Y2=2.765
r33 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.765 $X2=0.27 $Y2=2.765
r34 11 15 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=2.765
r35 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r36 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=2.765
r37 5 7 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=4.585
r38 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=2.765
r39 1 3 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_2%B 3 7 12 15 16
c41 7 0 1.37149e-19 $X=0.905 $Y=4.585
r42 16 18 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.59
r43 16 17 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.26
r44 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.425 $X2=0.95 $Y2=2.425
r45 11 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.425
r46 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.96
r47 7 18 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.59
r48 3 17 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_2%A_27_115# 1 2 9 11 13 15 16 20 22 24 25
+ 28 30 31 36 42 43 45 46 47
r87 48 49 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.935
+ $X2=1.37 $Y2=1.935
r88 46 47 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.545
+ $X2=0.65 $Y2=3.715
r89 43 49 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.43 $Y=1.935 $X2=1.37
+ $Y2=1.935
r90 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r91 40 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=0.61 $Y2=1.935
r92 40 42 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=1.43 $Y2=1.935
r93 36 38 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.69 $Y=3.795
+ $X2=0.69 $Y2=5.835
r94 36 47 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.795 $X2=0.69
+ $Y2=3.715
r95 32 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=2.02 $X2=0.61
+ $Y2=1.935
r96 32 46 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r97 30 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.61 $Y2=1.935
r98 30 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.345 $Y2=1.935
r99 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.345 $Y2=1.935
r100 26 28 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r101 22 24 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r102 18 43 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.43 $Y2=1.935
r103 18 20 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r104 17 25 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.885
+ $X2=1.352 $Y2=2.885
r105 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.96
r106 16 17 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.445 $Y2=2.885
r107 15 25 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.81
+ $X2=1.352 $Y2=2.885
r108 14 49 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=1.935
r109 14 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=2.81
r110 11 25 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.352 $Y2=2.885
r111 11 13 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r112 7 48 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.935
r113 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r114 2 38 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r115 2 36 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.795
r116 1 28 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__AND2_2%Y 1 2 10 13 17 18 21
c42 18 0 1.37149e-19 $X=1.55 $Y=2.59
r43 28 30 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r44 18 28 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r45 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r46 14 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r47 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r48 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r49 8 10 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r50 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r51 7 10 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r52 2 30 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r53 2 28 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r54 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

