* File: sky130_osu_sc_15T_hs__nor2_l.pex.spice
* Created: Fri Nov 12 14:32:06 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__NOR2_L%GND 1 2 21 25 27 35 41 44
r23 41 44 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r24 33 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.74
r25 27 33 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.305
r26 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r27 21 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r28 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r29 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r30 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r31 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r32 2 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.74
r33 1 25 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NOR2_L%VDD 1 13 15 21 27 30
r15 27 30 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r16 24 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r17 19 24 4.25596 $w=1.7e-07 $l=2.13185e-07 $layer=LI1_cond $X=1.05 $Y=5.245
+ $X2=1.197 $Y2=5.397
r18 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.05 $Y=5.245
+ $X2=1.05 $Y2=4.225
r19 15 24 3.30228 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=0.965 $Y=5.397
+ $X2=1.197 $Y2=5.397
r20 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=5.397
+ $X2=0.34 $Y2=5.397
r21 13 24 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r22 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r23 1 21 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=3.565 $X2=1.05 $Y2=4.225
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NOR2_L%B 3 7 10 13 19 22
r47 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.65 $Y=2.7 $X2=0.65
+ $Y2=2.7
r48 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.65 $Y=1.915
+ $X2=0.65 $Y2=2.7
r49 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=1.83
+ $X2=0.65 $Y2=1.915
r50 13 15 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.565 $Y=1.83
+ $X2=0.415 $Y2=1.83
r51 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.83 $X2=0.415 $Y2=1.83
r52 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.83
+ $X2=0.415 $Y2=1.995
r53 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.83
+ $X2=0.415 $Y2=1.665
r54 7 12 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.475 $Y=4.195
+ $X2=0.475 $Y2=1.995
r55 3 11 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=0.475 $Y=0.85
+ $X2=0.475 $Y2=1.665
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NOR2_L%A 3 7 10 14 20
r32 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=3.07
+ $X2=0.99 $Y2=3.07
r33 14 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.99 $Y=2.495
+ $X2=0.99 $Y2=3.07
r34 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.495 $X2=0.99 $Y2=2.495
r35 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.495
+ $X2=0.942 $Y2=2.66
r36 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.495
+ $X2=0.942 $Y2=2.33
r37 7 11 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=0.905 $Y=0.85
+ $X2=0.905 $Y2=2.33
r38 3 12 787.096 $w=1.5e-07 $l=1.535e-06 $layer=POLY_cond $X=0.835 $Y=4.195
+ $X2=0.835 $Y2=2.66
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NOR2_L%Y 1 3 10 16 21 22 26 32
r39 24 26 0.519956 $w=1.7e-07 $l=5.4e-07 $layer=MET1_cond $X=0.69 $Y=2.245
+ $X2=0.69 $Y2=1.705
r40 23 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.22
r41 23 26 0.356266 $w=1.7e-07 $l=3.7e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.705
r42 22 29 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=2.33
+ $X2=0.26 $Y2=2.33
r43 21 24 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=2.33
+ $X2=0.69 $Y2=2.245
r44 21 22 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=2.33
+ $X2=0.405 $Y2=2.33
r45 19 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.22
+ $X2=0.69 $Y2=1.22
r46 16 19 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.69 $Y=0.74
+ $X2=0.69 $Y2=1.22
r47 10 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.33
+ $X2=0.26 $Y2=2.33
r48 10 13 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=0.26 $Y=2.33
+ $X2=0.26 $Y2=4.225
r49 3 13 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.225
r50 1 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

