* File: sky130_osu_sc_12T_hs__tbufi_l.pex.spice
* Created: Fri Nov 12 15:13:25 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__TBUFI_L%GND 1 17 19 26 35 38
r36 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r37 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r38 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r39 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r40 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r41 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r42 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r43 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r44 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__TBUFI_L%VDD 1 13 15 21 25 29 32
r24 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r25 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r26 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r27 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287 $X2=1.02
+ $Y2=4.287
r28 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r29 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.275
r30 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r31 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r32 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r33 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r34 1 21 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.025 $X2=0.69 $Y2=3.275
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__TBUFI_L%OE 2 5 7 9 12 16 21 24 31 34
c62 31 0 2.60266e-19 $X=0.69 $Y=1.74
r63 28 31 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.855
+ $X2=0.69 $Y2=1.74
r64 28 34 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=0.69 $Y=1.855
+ $X2=0.69 $Y2=2.365
r65 24 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.74
+ $X2=0.69 $Y2=1.74
r66 21 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.74 $X2=0.69 $Y2=1.74
r67 14 16 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.825
+ $X2=0.475 $Y2=2.825
r68 10 21 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.69 $Y2=1.722
r69 10 12 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.905 $Y2=0.785
r70 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=2.825
r71 7 9 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=3.445
r72 3 21 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.69 $Y2=1.722
r73 3 5 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=0.785
r74 2 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.75 $X2=0.27
+ $Y2=2.825
r75 1 3 44.3094 $w=2.23e-07 $l=2.69768e-07 $layer=POLY_cond $X=0.27 $Y=1.69
+ $X2=0.475 $Y2=1.54
r76 1 2 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.69 $X2=0.27
+ $Y2=2.75
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__TBUFI_L%A_27_115# 1 3 11 16 20 24 26 28 31
r53 27 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.37
+ $X2=0.26 $Y2=2.37
r54 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.37
+ $X2=0.8 $Y2=2.37
r55 26 27 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=2.37
+ $X2=0.345 $Y2=2.37
r56 22 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.455
+ $X2=0.26 $Y2=2.37
r57 22 24 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.26 $Y=2.455
+ $X2=0.26 $Y2=3.275
r58 18 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.285
+ $X2=0.26 $Y2=2.37
r59 18 20 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=0.26 $Y=2.285
+ $X2=0.26 $Y2=0.74
r60 14 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=2.37 $X2=0.8 $Y2=2.37
r61 14 16 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.8 $Y=2.37
+ $X2=0.905 $Y2=2.37
r62 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.535
+ $X2=0.905 $Y2=2.37
r63 9 11 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=0.905 $Y=2.535
+ $X2=0.905 $Y2=3.445
r64 3 24 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.275
r65 1 20 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__TBUFI_L%A 3 7 10 15 20 23
c47 10 0 1.90743e-19 $X=1.325 $Y=1.98
c48 3 0 6.95226e-20 $X=1.265 $Y=0.785
r49 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.98
+ $X2=1.325 $Y2=1.98
r50 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=2.85
+ $X2=1.14 $Y2=2.85
r51 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.065
+ $X2=1.14 $Y2=1.98
r52 13 15 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.14 $Y=2.065
+ $X2=1.14 $Y2=2.85
r53 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.98 $X2=1.325 $Y2=1.98
r54 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.98
+ $X2=1.325 $Y2=2.145
r55 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.98
+ $X2=1.325 $Y2=1.815
r56 7 12 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=1.265 $Y=3.445
+ $X2=1.265 $Y2=2.145
r57 3 11 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=1.265 $Y=0.785
+ $X2=1.265 $Y2=1.815
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__TBUFI_L%Y 1 3 10 16 24 27 30
r34 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.365
+ $X2=1.48 $Y2=2.48
r35 22 24 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.365
+ $X2=1.48 $Y2=1.71
r36 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.485
+ $X2=1.48 $Y2=1.37
r37 21 24 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.485
+ $X2=1.48 $Y2=1.71
r38 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.48
+ $X2=1.48 $Y2=2.48
r39 16 19 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.48 $Y=2.48
+ $X2=1.48 $Y2=3.275
r40 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.37
+ $X2=1.48 $Y2=1.37
r41 10 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.48 $Y=0.74
+ $X2=1.48 $Y2=1.37
r42 3 19 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=3.025 $X2=1.48 $Y2=3.275
r43 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.74
.ends

