* File: sky130_osu_sc_12T_hs__inv_l.pxi.spice
* Created: Fri Nov 12 15:11:27 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__INV_L%GND N_GND_M1001_s N_GND_M1001_b N_GND_c_2_p
+ N_GND_c_3_p GND PM_SKY130_OSU_SC_12T_HS__INV_L%GND
x_PM_SKY130_OSU_SC_12T_HS__INV_L%VDD N_VDD_M1000_s N_VDD_M1000_b N_VDD_c_16_p
+ N_VDD_c_17_p VDD PM_SKY130_OSU_SC_12T_HS__INV_L%VDD
x_PM_SKY130_OSU_SC_12T_HS__INV_L%A N_A_M1001_g N_A_M1000_g N_A_c_31_n N_A_c_32_n
+ N_A_c_33_n N_A_c_34_n A PM_SKY130_OSU_SC_12T_HS__INV_L%A
x_PM_SKY130_OSU_SC_12T_HS__INV_L%Y N_Y_M1001_d N_Y_M1000_d N_Y_c_64_n N_Y_c_66_n
+ Y N_Y_c_68_n N_Y_c_69_n PM_SKY130_OSU_SC_12T_HS__INV_L%Y
cc_1 N_GND_M1001_b N_A_M1001_g 0.0817697f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.785
cc_2 N_GND_c_2_p N_A_M1001_g 0.00502587f $X=0.26 $Y=0.74 $X2=0.475 $Y2=0.785
cc_3 N_GND_c_3_p N_A_M1001_g 0.00468827f $X=0.34 $Y=0.19 $X2=0.475 $Y2=0.785
cc_4 N_GND_M1001_b N_A_M1000_g 0.0337175f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.435
cc_5 N_GND_M1001_b N_A_c_31_n 0.0392496f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_6 N_GND_M1001_b N_A_c_32_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.85
cc_7 N_GND_M1001_b N_A_c_33_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.825
cc_8 N_GND_M1001_b N_A_c_34_n 0.00255951f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_9 N_GND_M1001_b N_Y_c_64_n 0.0298613f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.74
cc_10 N_GND_c_3_p N_Y_c_64_n 0.00476261f $X=0.34 $Y=0.19 $X2=0.69 $Y2=0.74
cc_11 N_GND_M1001_b N_Y_c_66_n 0.00237997f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.48
cc_12 N_GND_M1001_b Y 0.0385097f $X=-0.045 $Y=0 $X2=0.755 $Y2=1.725
cc_13 N_GND_M1001_b N_Y_c_68_n 0.0157042f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.37
cc_14 N_GND_M1001_b N_Y_c_69_n 0.00507896f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.48
cc_15 N_VDD_M1000_b N_A_M1000_g 0.0589931f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.435
cc_16 N_VDD_c_16_p N_A_M1000_g 0.00713292f $X=0.26 $Y=3.605 $X2=0.475 $Y2=3.435
cc_17 N_VDD_c_17_p N_A_M1000_g 0.00606474f $X=0.34 $Y=4.24 $X2=0.475 $Y2=3.435
cc_18 VDD N_A_M1000_g 0.00468827f $X=0.34 $Y=4.19 $X2=0.475 $Y2=3.435
cc_19 N_VDD_M1000_b N_A_c_32_n 0.0147005f $X=-0.045 $Y=2.425 $X2=0.32 $Y2=2.85
cc_20 N_VDD_c_16_p N_A_c_32_n 0.00307077f $X=0.26 $Y=3.605 $X2=0.32 $Y2=2.85
cc_21 N_VDD_M1000_b A 0.0174587f $X=-0.045 $Y=2.425 $X2=0.32 $Y2=2.85
cc_22 N_VDD_c_16_p A 0.00542885f $X=0.26 $Y=3.605 $X2=0.32 $Y2=2.85
cc_23 N_VDD_M1000_b N_Y_c_66_n 0.0247014f $X=-0.045 $Y=2.425 $X2=0.69 $Y2=2.48
cc_24 N_VDD_c_17_p N_Y_c_66_n 0.00757793f $X=0.34 $Y=4.24 $X2=0.69 $Y2=2.48
cc_25 VDD N_Y_c_66_n 0.00476261f $X=0.34 $Y=4.19 $X2=0.69 $Y2=2.48
cc_26 N_VDD_M1000_b N_Y_c_69_n 0.00914195f $X=-0.045 $Y=2.425 $X2=0.69 $Y2=2.48
cc_27 N_A_M1001_g N_Y_c_64_n 0.0178582f $X=0.475 $Y=0.785 $X2=0.69 $Y2=0.74
cc_28 N_A_c_31_n N_Y_c_64_n 0.00108606f $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.74
cc_29 N_A_c_34_n N_Y_c_64_n 0.00388848f $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.74
cc_30 N_A_M1000_g N_Y_c_66_n 0.0226192f $X=0.475 $Y=3.435 $X2=0.69 $Y2=2.48
cc_31 N_A_c_31_n N_Y_c_66_n 8.13098e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_32 N_A_c_32_n N_Y_c_66_n 0.0305887f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_33 N_A_c_34_n N_Y_c_66_n 0.00202105f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_34 A N_Y_c_66_n 0.0149533f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_35 N_A_M1001_g Y 0.00406656f $X=0.475 $Y=0.785 $X2=0.755 $Y2=1.725
cc_36 N_A_M1000_g Y 0.00874077f $X=0.475 $Y=3.435 $X2=0.755 $Y2=1.725
cc_37 N_A_c_31_n Y 0.00700152f $X=0.535 $Y=1.825 $X2=0.755 $Y2=1.725
cc_38 N_A_c_32_n Y 0.0183799f $X=0.32 $Y=2.85 $X2=0.755 $Y2=1.725
cc_39 N_A_c_34_n Y 0.016989f $X=0.535 $Y=1.825 $X2=0.755 $Y2=1.725
cc_40 N_A_M1001_g N_Y_c_68_n 0.0118358f $X=0.475 $Y=0.785 $X2=0.69 $Y2=1.37
cc_41 N_A_c_31_n N_Y_c_68_n 0.0014188f $X=0.535 $Y=1.825 $X2=0.69 $Y2=1.37
cc_42 N_A_c_34_n N_Y_c_68_n 0.00238892f $X=0.535 $Y=1.825 $X2=0.69 $Y2=1.37
cc_43 N_A_M1000_g N_Y_c_69_n 0.00478745f $X=0.475 $Y=3.435 $X2=0.69 $Y2=2.48
cc_44 N_A_c_31_n N_Y_c_69_n 0.00126139f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_45 N_A_c_32_n N_Y_c_69_n 0.00640429f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_46 N_A_c_34_n N_Y_c_69_n 0.00194461f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_47 A N_Y_c_69_n 0.00827053f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
