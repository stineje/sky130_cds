magic
tech sky130A
magscale 1 2
timestamp 1612371642
<< nwell >>
rect -9 529 638 1119
<< nmoslvt >>
rect 80 115 110 243
rect 152 115 182 243
rect 252 115 282 243
rect 338 115 368 243
rect 424 115 454 243
rect 510 115 540 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
rect 338 565 368 965
rect 424 565 454 965
rect 510 565 540 965
<< ndiff >>
rect 27 229 80 243
rect 27 131 35 229
rect 69 131 80 229
rect 27 115 80 131
rect 110 115 152 243
rect 182 229 252 243
rect 182 131 193 229
rect 227 131 252 229
rect 182 115 252 131
rect 282 229 338 243
rect 282 131 293 229
rect 327 131 338 229
rect 282 115 338 131
rect 368 229 424 243
rect 368 131 379 229
rect 413 131 424 229
rect 368 115 424 131
rect 454 229 510 243
rect 454 131 465 229
rect 499 131 510 229
rect 454 115 510 131
rect 540 229 593 243
rect 540 131 551 229
rect 585 131 593 229
rect 540 115 593 131
<< pdiff >>
rect 27 949 80 965
rect 27 745 35 949
rect 69 745 80 949
rect 27 565 80 745
rect 110 949 166 965
rect 110 677 121 949
rect 155 677 166 949
rect 110 565 166 677
rect 196 949 252 965
rect 196 677 207 949
rect 241 677 252 949
rect 196 565 252 677
rect 282 949 338 965
rect 282 609 293 949
rect 327 609 338 949
rect 282 565 338 609
rect 368 949 424 965
rect 368 609 379 949
rect 413 609 424 949
rect 368 565 424 609
rect 454 949 510 965
rect 454 609 465 949
rect 499 609 510 949
rect 454 565 510 609
rect 540 949 593 965
rect 540 609 551 949
rect 585 609 593 949
rect 540 565 593 609
<< ndiffc >>
rect 35 131 69 229
rect 193 131 227 229
rect 293 131 327 229
rect 379 131 413 229
rect 465 131 499 229
rect 551 131 585 229
<< pdiffc >>
rect 35 745 69 949
rect 121 677 155 949
rect 207 677 241 949
rect 293 609 327 949
rect 379 609 413 949
rect 465 609 499 949
rect 551 609 585 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 991
rect 338 965 368 992
rect 424 965 454 991
rect 510 965 540 991
rect 80 534 110 565
rect 27 518 110 534
rect 27 484 37 518
rect 71 484 110 518
rect 27 468 110 484
rect 80 243 110 468
rect 166 466 196 565
rect 252 540 282 565
rect 338 540 368 565
rect 424 540 454 565
rect 510 540 540 565
rect 252 510 540 540
rect 152 450 217 466
rect 152 416 173 450
rect 207 416 217 450
rect 152 400 217 416
rect 152 243 182 400
rect 259 368 289 510
rect 259 352 313 368
rect 259 332 269 352
rect 252 318 269 332
rect 303 332 313 352
rect 303 318 540 332
rect 252 302 540 318
rect 252 243 282 302
rect 338 243 368 302
rect 424 243 454 302
rect 510 243 540 302
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
rect 338 89 368 115
rect 424 89 454 115
rect 510 89 540 115
<< polycont >>
rect 37 484 71 518
rect 173 416 207 450
rect 269 318 303 352
<< locali >>
rect 0 1089 638 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 638 1089
rect 35 949 69 1049
rect 35 729 69 745
rect 121 949 155 965
rect 105 677 121 695
rect 105 661 155 677
rect 207 949 241 1049
rect 207 661 241 677
rect 293 949 327 965
rect 37 518 71 597
rect 37 468 71 484
rect 105 352 139 661
rect 173 450 207 523
rect 293 483 327 609
rect 379 949 413 1049
rect 379 593 413 609
rect 465 949 499 965
rect 465 483 499 609
rect 551 949 585 1049
rect 551 593 585 609
rect 173 400 207 416
rect 35 318 269 352
rect 303 318 319 352
rect 35 229 69 318
rect 35 115 69 131
rect 193 229 227 249
rect 193 61 227 131
rect 293 115 327 131
rect 379 229 413 249
rect 379 61 413 131
rect 465 115 499 131
rect 551 229 585 249
rect 551 61 585 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 638 61
rect 0 0 638 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 37 597 71 631
rect 173 523 207 557
rect 293 449 327 483
rect 465 449 499 483
rect 293 229 327 261
rect 293 227 327 229
rect 465 229 499 261
rect 465 227 499 229
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1089 638 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 638 1089
rect 0 1049 638 1055
rect 25 631 83 637
rect 25 597 37 631
rect 71 597 105 631
rect 25 591 83 597
rect 161 557 219 563
rect 140 523 173 557
rect 207 523 219 557
rect 161 517 219 523
rect 281 483 339 489
rect 453 483 511 489
rect 281 449 293 483
rect 327 449 465 483
rect 499 449 511 483
rect 281 443 339 449
rect 453 443 511 449
rect 293 267 327 443
rect 465 267 499 443
rect 281 261 339 267
rect 453 261 511 267
rect 281 227 293 261
rect 327 227 465 261
rect 499 227 511 261
rect 281 221 339 227
rect 453 221 511 227
rect 0 55 638 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 638 55
rect 0 0 638 21
<< labels >>
rlabel metal1 311 392 311 392 1 Y
port 1 n
rlabel viali 55 614 55 614 1 A
port 2 n
rlabel viali 191 540 191 540 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
