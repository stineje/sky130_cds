* File: sky130_osu_sc_12T_ms__and2_6.pxi.spice
* Created: Fri Nov 12 15:20:34 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__AND2_6%GND N_GND_M1002_d N_GND_M1009_s N_GND_M1013_s
+ N_GND_M1015_s N_GND_M1005_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p N_GND_c_23_p
+ N_GND_c_30_p N_GND_c_36_p N_GND_c_43_p N_GND_c_50_p GND N_GND_c_3_p
+ PM_SKY130_OSU_SC_12T_MS__AND2_6%GND
x_PM_SKY130_OSU_SC_12T_MS__AND2_6%VDD N_VDD_M1001_s N_VDD_M1010_d N_VDD_M1004_s
+ N_VDD_M1007_s N_VDD_M1012_s N_VDD_M1001_b N_VDD_c_114_p N_VDD_c_115_p
+ N_VDD_c_126_p N_VDD_c_133_p N_VDD_c_139_p N_VDD_c_145_p N_VDD_c_150_p
+ N_VDD_c_156_p N_VDD_c_161_p VDD N_VDD_c_116_p
+ PM_SKY130_OSU_SC_12T_MS__AND2_6%VDD
x_PM_SKY130_OSU_SC_12T_MS__AND2_6%A N_A_M1005_g N_A_M1001_g N_A_c_186_n
+ N_A_c_187_n A PM_SKY130_OSU_SC_12T_MS__AND2_6%A
x_PM_SKY130_OSU_SC_12T_MS__AND2_6%B N_B_M1002_g N_B_M1010_g N_B_c_217_n
+ N_B_c_218_n B PM_SKY130_OSU_SC_12T_MS__AND2_6%B
x_PM_SKY130_OSU_SC_12T_MS__AND2_6%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1001_d N_A_27_115#_M1000_g N_A_27_115#_c_254_n
+ N_A_27_115#_c_305_n N_A_27_115#_M1003_g N_A_27_115#_c_255_n
+ N_A_27_115#_c_256_n N_A_27_115#_M1009_g N_A_27_115#_c_310_n
+ N_A_27_115#_M1004_g N_A_27_115#_c_261_n N_A_27_115#_c_263_n
+ N_A_27_115#_M1011_g N_A_27_115#_c_317_n N_A_27_115#_M1006_g
+ N_A_27_115#_c_268_n N_A_27_115#_c_269_n N_A_27_115#_M1013_g
+ N_A_27_115#_c_322_n N_A_27_115#_M1007_g N_A_27_115#_c_274_n
+ N_A_27_115#_c_276_n N_A_27_115#_M1014_g N_A_27_115#_c_281_n
+ N_A_27_115#_c_328_n N_A_27_115#_M1008_g N_A_27_115#_c_282_n
+ N_A_27_115#_c_283_n N_A_27_115#_M1015_g N_A_27_115#_c_333_n
+ N_A_27_115#_M1012_g N_A_27_115#_c_288_n N_A_27_115#_c_289_n
+ N_A_27_115#_c_290_n N_A_27_115#_c_291_n N_A_27_115#_c_292_n
+ N_A_27_115#_c_293_n N_A_27_115#_c_294_n N_A_27_115#_c_295_n
+ N_A_27_115#_c_296_n N_A_27_115#_c_297_n N_A_27_115#_c_298_n
+ N_A_27_115#_c_301_n N_A_27_115#_c_343_n N_A_27_115#_c_302_n
+ N_A_27_115#_c_303_n N_A_27_115#_c_355_n
+ PM_SKY130_OSU_SC_12T_MS__AND2_6%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__AND2_6%Y N_Y_M1000_d N_Y_M1011_d N_Y_M1014_d
+ N_Y_M1003_d N_Y_M1006_d N_Y_M1008_d N_Y_c_438_n N_Y_c_443_n N_Y_c_444_n
+ N_Y_c_449_n N_Y_c_450_n N_Y_c_454_n N_Y_c_455_n N_Y_c_459_n Y N_Y_c_461_n
+ N_Y_c_465_n N_Y_c_466_n N_Y_c_467_n N_Y_c_471_n N_Y_c_475_n N_Y_c_476_n
+ N_Y_c_477_n N_Y_c_481_n PM_SKY130_OSU_SC_12T_MS__AND2_6%Y
cc_1 N_GND_M1005_b N_A_M1005_g 0.0805447f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1005_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_A_M1005_g 0.00468827f $X=3.06 $Y=0.19 $X2=0.475 $Y2=0.835
cc_4 N_GND_M1005_b N_A_c_186_n 0.0447183f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.285
cc_5 N_GND_M1005_b N_A_c_187_n 0.00329519f $X=-0.045 $Y=0 $X2=0.235 $Y2=2.285
cc_6 N_GND_M1005_b N_B_M1002_g 0.0456699f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.835
cc_7 N_GND_c_2_p N_B_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.835
cc_8 N_GND_c_8_p N_B_M1002_g 0.00319969f $X=1.05 $Y=0.755 $X2=0.835 $Y2=0.835
cc_9 N_GND_c_3_p N_B_M1002_g 0.00468827f $X=3.06 $Y=0.19 $X2=0.835 $Y2=0.835
cc_10 N_GND_M1005_b N_B_M1010_g 0.0145087f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_11 N_GND_M1005_b N_B_c_217_n 0.0304191f $X=-0.045 $Y=0 $X2=0.915 $Y2=1.945
cc_12 N_GND_M1005_b N_B_c_218_n 0.00352155f $X=-0.045 $Y=0 $X2=0.915 $Y2=1.945
cc_13 N_GND_M1005_b B 0.00685421f $X=-0.045 $Y=0 $X2=0.92 $Y2=2.48
cc_14 N_GND_M1005_b N_A_27_115#_M1000_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.835
cc_15 N_GND_c_8_p N_A_27_115#_M1000_g 0.00610843f $X=1.05 $Y=0.755 $X2=1.335
+ $Y2=0.835
cc_16 N_GND_c_16_p N_A_27_115#_M1000_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.835
cc_17 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=3.06 $Y=0.19 $X2=1.335
+ $Y2=0.835
cc_18 N_GND_M1005_b N_A_27_115#_c_254_n 0.0465667f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=2.33
cc_19 N_GND_M1005_b N_A_27_115#_c_255_n 0.00863342f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.405
cc_20 N_GND_M1005_b N_A_27_115#_c_256_n 0.0104564f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.365
cc_21 N_GND_M1005_b N_A_27_115#_M1009_g 0.0202142f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.835
cc_22 N_GND_c_16_p N_A_27_115#_M1009_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.835
cc_23 N_GND_c_23_p N_A_27_115#_M1009_g 0.00311745f $X=1.98 $Y=0.755 $X2=1.765
+ $Y2=0.835
cc_24 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=3.06 $Y=0.19 $X2=1.765
+ $Y2=0.835
cc_25 N_GND_M1005_b N_A_27_115#_c_261_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.365
cc_26 N_GND_c_23_p N_A_27_115#_c_261_n 0.00256938f $X=1.98 $Y=0.755 $X2=2.12
+ $Y2=1.365
cc_27 N_GND_M1005_b N_A_27_115#_c_263_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.405
cc_28 N_GND_M1005_b N_A_27_115#_M1011_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.835
cc_29 N_GND_c_23_p N_A_27_115#_M1011_g 0.00311745f $X=1.98 $Y=0.755 $X2=2.195
+ $Y2=0.835
cc_30 N_GND_c_30_p N_A_27_115#_M1011_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.835
cc_31 N_GND_c_3_p N_A_27_115#_M1011_g 0.00468827f $X=3.06 $Y=0.19 $X2=2.195
+ $Y2=0.835
cc_32 N_GND_M1005_b N_A_27_115#_c_268_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.365
cc_33 N_GND_M1005_b N_A_27_115#_c_269_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.405
cc_34 N_GND_M1005_b N_A_27_115#_M1013_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.835
cc_35 N_GND_c_30_p N_A_27_115#_M1013_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.835
cc_36 N_GND_c_36_p N_A_27_115#_M1013_g 0.00311745f $X=2.84 $Y=0.755 $X2=2.625
+ $Y2=0.835
cc_37 N_GND_c_3_p N_A_27_115#_M1013_g 0.00468827f $X=3.06 $Y=0.19 $X2=2.625
+ $Y2=0.835
cc_38 N_GND_M1005_b N_A_27_115#_c_274_n 0.0181078f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.365
cc_39 N_GND_c_36_p N_A_27_115#_c_274_n 0.00256938f $X=2.84 $Y=0.755 $X2=2.98
+ $Y2=1.365
cc_40 N_GND_M1005_b N_A_27_115#_c_276_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.405
cc_41 N_GND_M1005_b N_A_27_115#_M1014_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.835
cc_42 N_GND_c_36_p N_A_27_115#_M1014_g 0.00311745f $X=2.84 $Y=0.755 $X2=3.055
+ $Y2=0.835
cc_43 N_GND_c_43_p N_A_27_115#_M1014_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.055
+ $Y2=0.835
cc_44 N_GND_c_3_p N_A_27_115#_M1014_g 0.00468827f $X=3.06 $Y=0.19 $X2=3.055
+ $Y2=0.835
cc_45 N_GND_M1005_b N_A_27_115#_c_281_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.33
cc_46 N_GND_M1005_b N_A_27_115#_c_282_n 0.0369419f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.365
cc_47 N_GND_M1005_b N_A_27_115#_c_283_n 0.0268552f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.405
cc_48 N_GND_M1005_b N_A_27_115#_M1015_g 0.0264941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=0.835
cc_49 N_GND_c_43_p N_A_27_115#_M1015_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.485
+ $Y2=0.835
cc_50 N_GND_c_50_p N_A_27_115#_M1015_g 0.00502587f $X=3.7 $Y=0.755 $X2=3.485
+ $Y2=0.835
cc_51 N_GND_c_3_p N_A_27_115#_M1015_g 0.00468827f $X=3.06 $Y=0.19 $X2=3.485
+ $Y2=0.835
cc_52 N_GND_M1005_b N_A_27_115#_c_288_n 0.0264756f $X=-0.045 $Y=0 $X2=1.395
+ $Y2=1.365
cc_53 N_GND_M1005_b N_A_27_115#_c_289_n 0.00339913f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=2.405
cc_54 N_GND_M1005_b N_A_27_115#_c_290_n 0.00873941f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.365
cc_55 N_GND_M1005_b N_A_27_115#_c_291_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.405
cc_56 N_GND_M1005_b N_A_27_115#_c_292_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.365
cc_57 N_GND_M1005_b N_A_27_115#_c_293_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.405
cc_58 N_GND_M1005_b N_A_27_115#_c_294_n 0.00873941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.365
cc_59 N_GND_M1005_b N_A_27_115#_c_295_n 0.00735657f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.405
cc_60 N_GND_M1005_b N_A_27_115#_c_296_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.365
cc_61 N_GND_M1005_b N_A_27_115#_c_297_n 0.00151234f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.405
cc_62 N_GND_M1005_b N_A_27_115#_c_298_n 0.0148636f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_63 N_GND_c_2_p N_A_27_115#_c_298_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_64 N_GND_c_3_p N_A_27_115#_c_298_n 0.00476261f $X=3.06 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_65 N_GND_M1005_b N_A_27_115#_c_301_n 0.00626966f $X=-0.045 $Y=0 $X2=0.575
+ $Y2=3.065
cc_66 N_GND_M1005_b N_A_27_115#_c_302_n 0.0164401f $X=-0.045 $Y=0 $X2=0.66
+ $Y2=1.455
cc_67 N_GND_M1005_b N_A_27_115#_c_303_n 0.0251886f $X=-0.045 $Y=0 $X2=1.395
+ $Y2=1.455
cc_68 N_GND_c_8_p N_A_27_115#_c_303_n 0.00704977f $X=1.05 $Y=0.755 $X2=1.395
+ $Y2=1.455
cc_69 N_GND_M1005_b N_Y_c_438_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_70 N_GND_c_8_p N_Y_c_438_n 0.00806382f $X=1.05 $Y=0.755 $X2=1.55 $Y2=0.755
cc_71 N_GND_c_16_p N_Y_c_438_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_72 N_GND_c_23_p N_Y_c_438_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=0.755
cc_73 N_GND_c_3_p N_Y_c_438_n 0.0047139f $X=3.06 $Y=0.19 $X2=1.55 $Y2=0.755
cc_74 N_GND_M1005_b N_Y_c_443_n 0.0110121f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_75 N_GND_M1005_b N_Y_c_444_n 0.00154299f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.755
cc_76 N_GND_c_23_p N_Y_c_444_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=2.41 $Y2=0.755
cc_77 N_GND_c_30_p N_Y_c_444_n 0.00718527f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.755
cc_78 N_GND_c_36_p N_Y_c_444_n 8.14297e-19 $X=2.84 $Y=0.755 $X2=2.41 $Y2=0.755
cc_79 N_GND_c_3_p N_Y_c_444_n 0.0047139f $X=3.06 $Y=0.19 $X2=2.41 $Y2=0.755
cc_80 N_GND_M1005_b N_Y_c_449_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.11
cc_81 N_GND_M1005_b N_Y_c_450_n 0.00154299f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.755
cc_82 N_GND_c_36_p N_Y_c_450_n 8.14297e-19 $X=2.84 $Y=0.755 $X2=3.27 $Y2=0.755
cc_83 N_GND_c_43_p N_Y_c_450_n 0.00729945f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.755
cc_84 N_GND_c_3_p N_Y_c_450_n 0.0047139f $X=3.06 $Y=0.19 $X2=3.27 $Y2=0.755
cc_85 N_GND_M1005_b N_Y_c_454_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.11
cc_86 N_GND_M1005_b N_Y_c_455_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.115
cc_87 N_GND_c_8_p N_Y_c_455_n 0.00127231f $X=1.05 $Y=0.755 $X2=1.55 $Y2=1.115
cc_88 N_GND_c_16_p N_Y_c_455_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.55 $Y2=1.115
cc_89 N_GND_c_23_p N_Y_c_455_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=1.115
cc_90 N_GND_M1005_b N_Y_c_459_n 0.00675046f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.995
cc_91 N_GND_M1005_b Y 0.030773f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.74
cc_92 N_GND_M1009_s N_Y_c_461_n 0.0100329f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1
cc_93 N_GND_c_16_p N_Y_c_461_n 0.0028844f $X=1.895 $Y=0.152 $X2=2.265 $Y2=1
cc_94 N_GND_c_23_p N_Y_c_461_n 0.0142303f $X=1.98 $Y=0.755 $X2=2.265 $Y2=1
cc_95 N_GND_c_30_p N_Y_c_461_n 0.0028844f $X=2.755 $Y=0.152 $X2=2.265 $Y2=1
cc_96 N_GND_M1005_b N_Y_c_465_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.11
cc_97 N_GND_M1005_b N_Y_c_466_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.995
cc_98 N_GND_M1013_s N_Y_c_467_n 0.0100329f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1
cc_99 N_GND_c_30_p N_Y_c_467_n 0.0028844f $X=2.755 $Y=0.152 $X2=3.125 $Y2=1
cc_100 N_GND_c_36_p N_Y_c_467_n 0.0142303f $X=2.84 $Y=0.755 $X2=3.125 $Y2=1
cc_101 N_GND_c_43_p N_Y_c_467_n 0.0028844f $X=3.615 $Y=0.152 $X2=3.125 $Y2=1
cc_102 N_GND_M1005_b N_Y_c_471_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1
cc_103 N_GND_c_23_p N_Y_c_471_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=2.555 $Y2=1
cc_104 N_GND_c_30_p N_Y_c_471_n 0.00245319f $X=2.755 $Y=0.152 $X2=2.555 $Y2=1
cc_105 N_GND_c_36_p N_Y_c_471_n 7.53951e-19 $X=2.84 $Y=0.755 $X2=2.555 $Y2=1
cc_106 N_GND_M1005_b N_Y_c_475_n 0.0144211f $X=-0.045 $Y=0 $X2=3.125 $Y2=2.11
cc_107 N_GND_M1005_b N_Y_c_476_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.11
cc_108 N_GND_M1005_b N_Y_c_477_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.115
cc_109 N_GND_c_36_p N_Y_c_477_n 7.53951e-19 $X=2.84 $Y=0.755 $X2=3.27 $Y2=1.115
cc_110 N_GND_c_43_p N_Y_c_477_n 0.00245319f $X=3.615 $Y=0.152 $X2=3.27 $Y2=1.115
cc_111 N_GND_c_50_p N_Y_c_477_n 0.00134236f $X=3.7 $Y=0.755 $X2=3.27 $Y2=1.115
cc_112 N_GND_M1005_b N_Y_c_481_n 0.0485933f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.995
cc_113 N_VDD_M1001_b N_A_M1001_g 0.0189715f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_114 N_VDD_c_114_p N_A_M1001_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_115 N_VDD_c_115_p N_A_M1001_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_116 N_VDD_c_116_p N_A_M1001_g 0.00468827f $X=3.06 $Y=4.25 $X2=0.475 $Y2=3.235
cc_117 N_VDD_M1001_b N_A_c_186_n 0.0124943f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.285
cc_118 N_VDD_M1001_s N_A_c_187_n 0.0150633f $X=0.135 $Y=2.605 $X2=0.235
+ $Y2=2.285
cc_119 N_VDD_M1001_b N_A_c_187_n 0.00613107f $X=-0.045 $Y=2.425 $X2=0.235
+ $Y2=2.285
cc_120 N_VDD_c_114_p N_A_c_187_n 0.00337102f $X=0.26 $Y=3.635 $X2=0.235
+ $Y2=2.285
cc_121 N_VDD_M1001_s A 0.00790556f $X=0.135 $Y=2.605 $X2=0.24 $Y2=2.85
cc_122 N_VDD_M1001_b A 0.0115315f $X=-0.045 $Y=2.425 $X2=0.24 $Y2=2.85
cc_123 N_VDD_c_114_p A 0.00459217f $X=0.26 $Y=3.635 $X2=0.24 $Y2=2.85
cc_124 N_VDD_M1001_b N_B_M1010_g 0.0187479f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_125 N_VDD_c_115_p N_B_M1010_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905
+ $Y2=3.235
cc_126 N_VDD_c_126_p N_B_M1010_g 0.00337744f $X=1.12 $Y=3.295 $X2=0.905
+ $Y2=3.235
cc_127 N_VDD_c_116_p N_B_M1010_g 0.00468827f $X=3.06 $Y=4.25 $X2=0.905 $Y2=3.235
cc_128 N_VDD_M1001_b N_B_c_218_n 0.00130234f $X=-0.045 $Y=2.425 $X2=0.915
+ $Y2=1.945
cc_129 N_VDD_M1001_b B 0.00872506f $X=-0.045 $Y=2.425 $X2=0.92 $Y2=2.48
cc_130 N_VDD_c_126_p B 9.65504e-19 $X=1.12 $Y=3.295 $X2=0.92 $Y2=2.48
cc_131 N_VDD_M1001_b N_A_27_115#_c_305_n 0.0171069f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.48
cc_132 N_VDD_c_126_p N_A_27_115#_c_305_n 0.00337744f $X=1.12 $Y=3.295 $X2=1.335
+ $Y2=2.48
cc_133 N_VDD_c_133_p N_A_27_115#_c_305_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335
+ $Y2=2.48
cc_134 N_VDD_c_116_p N_A_27_115#_c_305_n 0.00468827f $X=3.06 $Y=4.25 $X2=1.335
+ $Y2=2.48
cc_135 N_VDD_M1001_b N_A_27_115#_c_255_n 0.00448664f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_136 N_VDD_M1001_b N_A_27_115#_c_310_n 0.017006f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.48
cc_137 N_VDD_c_126_p N_A_27_115#_c_310_n 3.67508e-19 $X=1.12 $Y=3.295 $X2=1.765
+ $Y2=2.48
cc_138 N_VDD_c_133_p N_A_27_115#_c_310_n 0.00610567f $X=1.895 $Y=4.287 $X2=1.765
+ $Y2=2.48
cc_139 N_VDD_c_139_p N_A_27_115#_c_310_n 0.0035715f $X=1.98 $Y=2.955 $X2=1.765
+ $Y2=2.48
cc_140 N_VDD_c_116_p N_A_27_115#_c_310_n 0.00470215f $X=3.06 $Y=4.25 $X2=1.765
+ $Y2=2.48
cc_141 N_VDD_M1001_b N_A_27_115#_c_263_n 0.00396043f $X=-0.045 $Y=2.425 $X2=2.12
+ $Y2=2.405
cc_142 N_VDD_c_139_p N_A_27_115#_c_263_n 0.00379272f $X=1.98 $Y=2.955 $X2=2.12
+ $Y2=2.405
cc_143 N_VDD_M1001_b N_A_27_115#_c_317_n 0.0166898f $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.48
cc_144 N_VDD_c_139_p N_A_27_115#_c_317_n 0.00337744f $X=1.98 $Y=2.955 $X2=2.195
+ $Y2=2.48
cc_145 N_VDD_c_145_p N_A_27_115#_c_317_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.195
+ $Y2=2.48
cc_146 N_VDD_c_116_p N_A_27_115#_c_317_n 0.00468827f $X=3.06 $Y=4.25 $X2=2.195
+ $Y2=2.48
cc_147 N_VDD_M1001_b N_A_27_115#_c_269_n 0.00448664f $X=-0.045 $Y=2.425 $X2=2.55
+ $Y2=2.405
cc_148 N_VDD_M1001_b N_A_27_115#_c_322_n 0.0166898f $X=-0.045 $Y=2.425 $X2=2.625
+ $Y2=2.48
cc_149 N_VDD_c_145_p N_A_27_115#_c_322_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.625
+ $Y2=2.48
cc_150 N_VDD_c_150_p N_A_27_115#_c_322_n 0.00337744f $X=2.84 $Y=2.955 $X2=2.625
+ $Y2=2.48
cc_151 N_VDD_c_116_p N_A_27_115#_c_322_n 0.00468827f $X=3.06 $Y=4.25 $X2=2.625
+ $Y2=2.48
cc_152 N_VDD_M1001_b N_A_27_115#_c_276_n 0.00396043f $X=-0.045 $Y=2.425 $X2=2.98
+ $Y2=2.405
cc_153 N_VDD_c_150_p N_A_27_115#_c_276_n 0.00379272f $X=2.84 $Y=2.955 $X2=2.98
+ $Y2=2.405
cc_154 N_VDD_M1001_b N_A_27_115#_c_328_n 0.0166898f $X=-0.045 $Y=2.425 $X2=3.055
+ $Y2=2.48
cc_155 N_VDD_c_150_p N_A_27_115#_c_328_n 0.00337744f $X=2.84 $Y=2.955 $X2=3.055
+ $Y2=2.48
cc_156 N_VDD_c_156_p N_A_27_115#_c_328_n 0.00606474f $X=3.615 $Y=4.287 $X2=3.055
+ $Y2=2.48
cc_157 N_VDD_c_116_p N_A_27_115#_c_328_n 0.00468827f $X=3.06 $Y=4.25 $X2=3.055
+ $Y2=2.48
cc_158 N_VDD_M1001_b N_A_27_115#_c_283_n 0.00840215f $X=-0.045 $Y=2.425 $X2=3.41
+ $Y2=2.405
cc_159 N_VDD_M1001_b N_A_27_115#_c_333_n 0.0209036f $X=-0.045 $Y=2.425 $X2=3.485
+ $Y2=2.48
cc_160 N_VDD_c_156_p N_A_27_115#_c_333_n 0.00606474f $X=3.615 $Y=4.287 $X2=3.485
+ $Y2=2.48
cc_161 N_VDD_c_161_p N_A_27_115#_c_333_n 0.00636672f $X=3.7 $Y=2.955 $X2=3.485
+ $Y2=2.48
cc_162 N_VDD_c_116_p N_A_27_115#_c_333_n 0.00468827f $X=3.06 $Y=4.25 $X2=3.485
+ $Y2=2.48
cc_163 N_VDD_M1001_b N_A_27_115#_c_289_n 0.00196792f $X=-0.045 $Y=2.425
+ $X2=1.335 $Y2=2.405
cc_164 N_VDD_M1001_b N_A_27_115#_c_291_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=1.765 $Y2=2.405
cc_165 N_VDD_M1001_b N_A_27_115#_c_293_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=2.195 $Y2=2.405
cc_166 N_VDD_M1001_b N_A_27_115#_c_295_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=2.625 $Y2=2.405
cc_167 N_VDD_M1001_b N_A_27_115#_c_297_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=3.055 $Y2=2.405
cc_168 N_VDD_M1001_b N_A_27_115#_c_301_n 8.35397e-19 $X=-0.045 $Y=2.425
+ $X2=0.575 $Y2=3.065
cc_169 N_VDD_M1001_b N_A_27_115#_c_343_n 0.001549f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=3.295
cc_170 N_VDD_c_115_p N_A_27_115#_c_343_n 0.00751386f $X=1.035 $Y=4.287 $X2=0.69
+ $Y2=3.295
cc_171 N_VDD_c_116_p N_A_27_115#_c_343_n 0.00474587f $X=3.06 $Y=4.25 $X2=0.69
+ $Y2=3.295
cc_172 N_VDD_M1001_b N_Y_c_443_n 0.00347838f $X=-0.045 $Y=2.425 $X2=1.55
+ $Y2=2.11
cc_173 N_VDD_c_133_p N_Y_c_443_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.11
cc_174 N_VDD_c_116_p N_Y_c_443_n 0.00475776f $X=3.06 $Y=4.25 $X2=1.55 $Y2=2.11
cc_175 N_VDD_M1001_b N_Y_c_449_n 0.00380347f $X=-0.045 $Y=2.425 $X2=2.41
+ $Y2=2.11
cc_176 N_VDD_c_145_p N_Y_c_449_n 0.00734006f $X=2.755 $Y=4.287 $X2=2.41 $Y2=2.11
cc_177 N_VDD_c_116_p N_Y_c_449_n 0.00475776f $X=3.06 $Y=4.25 $X2=2.41 $Y2=2.11
cc_178 N_VDD_M1001_b N_Y_c_454_n 0.00380347f $X=-0.045 $Y=2.425 $X2=3.27
+ $Y2=2.11
cc_179 N_VDD_c_156_p N_Y_c_454_n 0.00745425f $X=3.615 $Y=4.287 $X2=3.27 $Y2=2.11
cc_180 N_VDD_c_116_p N_Y_c_454_n 0.00475776f $X=3.06 $Y=4.25 $X2=3.27 $Y2=2.11
cc_181 N_VDD_c_139_p N_Y_c_465_n 0.00634153f $X=1.98 $Y=2.955 $X2=2.265 $Y2=2.11
cc_182 N_VDD_c_150_p N_Y_c_475_n 0.00634153f $X=2.84 $Y=2.955 $X2=3.125 $Y2=2.11
cc_183 N_A_M1005_g N_B_M1002_g 0.101444f $X=0.475 $Y=0.835 $X2=0.835 $Y2=0.835
cc_184 N_A_M1005_g N_B_M1010_g 0.0482865f $X=0.475 $Y=0.835 $X2=0.905 $Y2=3.235
cc_185 N_A_M1005_g N_B_c_218_n 8.69605e-19 $X=0.475 $Y=0.835 $X2=0.915 $Y2=1.945
cc_186 N_A_M1005_g N_A_27_115#_c_298_n 0.0134311f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.755
cc_187 N_A_M1005_g N_A_27_115#_c_301_n 0.0278506f $X=0.475 $Y=0.835 $X2=0.575
+ $Y2=3.065
cc_188 N_A_M1001_g N_A_27_115#_c_301_n 0.0152191f $X=0.475 $Y=3.235 $X2=0.575
+ $Y2=3.065
cc_189 N_A_c_186_n N_A_27_115#_c_301_n 0.00844699f $X=0.475 $Y=2.285 $X2=0.575
+ $Y2=3.065
cc_190 N_A_c_187_n N_A_27_115#_c_301_n 0.053763f $X=0.235 $Y=2.285 $X2=0.575
+ $Y2=3.065
cc_191 A N_A_27_115#_c_301_n 0.00781918f $X=0.24 $Y=2.85 $X2=0.575 $Y2=3.065
cc_192 N_A_M1005_g N_A_27_115#_c_302_n 0.0178909f $X=0.475 $Y=0.835 $X2=0.66
+ $Y2=1.455
cc_193 N_A_c_186_n N_A_27_115#_c_302_n 0.00272689f $X=0.475 $Y=2.285 $X2=0.66
+ $Y2=1.455
cc_194 N_A_c_187_n N_A_27_115#_c_302_n 0.00451097f $X=0.235 $Y=2.285 $X2=0.66
+ $Y2=1.455
cc_195 N_A_M1001_g N_A_27_115#_c_355_n 0.0107221f $X=0.475 $Y=3.235 $X2=0.69
+ $Y2=3.15
cc_196 N_B_M1002_g N_A_27_115#_M1000_g 0.0390746f $X=0.835 $Y=0.835 $X2=1.335
+ $Y2=0.835
cc_197 N_B_M1010_g N_A_27_115#_c_254_n 0.0478471f $X=0.905 $Y=3.235 $X2=1.335
+ $Y2=2.33
cc_198 N_B_c_217_n N_A_27_115#_c_254_n 0.0207593f $X=0.915 $Y=1.945 $X2=1.335
+ $Y2=2.33
cc_199 N_B_c_218_n N_A_27_115#_c_254_n 0.00498982f $X=0.915 $Y=1.945 $X2=1.335
+ $Y2=2.33
cc_200 B N_A_27_115#_c_289_n 0.00380362f $X=0.92 $Y=2.48 $X2=1.335 $Y2=2.405
cc_201 N_B_M1002_g N_A_27_115#_c_301_n 0.00719886f $X=0.835 $Y=0.835 $X2=0.575
+ $Y2=3.065
cc_202 N_B_M1010_g N_A_27_115#_c_301_n 0.01267f $X=0.905 $Y=3.235 $X2=0.575
+ $Y2=3.065
cc_203 N_B_c_218_n N_A_27_115#_c_301_n 0.0541394f $X=0.915 $Y=1.945 $X2=0.575
+ $Y2=3.065
cc_204 B N_A_27_115#_c_301_n 0.00871807f $X=0.92 $Y=2.48 $X2=0.575 $Y2=3.065
cc_205 N_B_M1002_g N_A_27_115#_c_303_n 0.0171085f $X=0.835 $Y=0.835 $X2=1.395
+ $Y2=1.455
cc_206 N_B_c_217_n N_A_27_115#_c_303_n 0.00235847f $X=0.915 $Y=1.945 $X2=1.395
+ $Y2=1.455
cc_207 N_B_c_218_n N_A_27_115#_c_303_n 0.0100447f $X=0.915 $Y=1.945 $X2=1.395
+ $Y2=1.455
cc_208 B N_A_27_115#_c_355_n 0.00385574f $X=0.92 $Y=2.48 $X2=0.69 $Y2=3.15
cc_209 N_B_c_218_n N_Y_c_443_n 0.0138653f $X=0.915 $Y=1.945 $X2=1.55 $Y2=2.11
cc_210 B N_Y_c_443_n 0.00632423f $X=0.92 $Y=2.48 $X2=1.55 $Y2=2.11
cc_211 N_B_M1002_g N_Y_c_455_n 7.93934e-19 $X=0.835 $Y=0.835 $X2=1.55 $Y2=1.115
cc_212 N_B_c_217_n N_Y_c_459_n 5.80618e-19 $X=0.915 $Y=1.945 $X2=1.55 $Y2=1.995
cc_213 N_B_c_218_n N_Y_c_459_n 0.00573285f $X=0.915 $Y=1.945 $X2=1.55 $Y2=1.995
cc_214 N_B_M1002_g Y 6.5988e-19 $X=0.835 $Y=0.835 $X2=1.555 $Y2=1.74
cc_215 N_B_c_218_n Y 0.00671947f $X=0.915 $Y=1.945 $X2=1.555 $Y2=1.74
cc_216 N_A_27_115#_M1000_g N_Y_c_438_n 0.00184843f $X=1.335 $Y=0.835 $X2=1.55
+ $Y2=0.755
cc_217 N_A_27_115#_M1009_g N_Y_c_438_n 0.00182852f $X=1.765 $Y=0.835 $X2=1.55
+ $Y2=0.755
cc_218 N_A_27_115#_c_288_n N_Y_c_438_n 0.0020555f $X=1.395 $Y=1.365 $X2=1.55
+ $Y2=0.755
cc_219 N_A_27_115#_c_303_n N_Y_c_438_n 0.00363898f $X=1.395 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_220 N_A_27_115#_c_254_n N_Y_c_443_n 0.00711959f $X=1.335 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_221 N_A_27_115#_c_305_n N_Y_c_443_n 0.00265429f $X=1.335 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_222 N_A_27_115#_c_255_n N_Y_c_443_n 0.0163883f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_223 N_A_27_115#_c_256_n N_Y_c_443_n 0.00122399f $X=1.69 $Y=1.365 $X2=1.55
+ $Y2=2.11
cc_224 N_A_27_115#_c_310_n N_Y_c_443_n 0.00375894f $X=1.765 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_225 N_A_27_115#_c_288_n N_Y_c_443_n 6.59752e-19 $X=1.395 $Y=1.365 $X2=1.55
+ $Y2=2.11
cc_226 N_A_27_115#_c_303_n N_Y_c_443_n 0.00202105f $X=1.395 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_227 N_A_27_115#_M1011_g N_Y_c_444_n 0.00182852f $X=2.195 $Y=0.835 $X2=2.41
+ $Y2=0.755
cc_228 N_A_27_115#_c_268_n N_Y_c_444_n 0.00274041f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=0.755
cc_229 N_A_27_115#_M1013_g N_Y_c_444_n 0.00182852f $X=2.625 $Y=0.835 $X2=2.41
+ $Y2=0.755
cc_230 N_A_27_115#_c_317_n N_Y_c_449_n 0.00375894f $X=2.195 $Y=2.48 $X2=2.41
+ $Y2=2.11
cc_231 N_A_27_115#_c_268_n N_Y_c_449_n 0.00250559f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=2.11
cc_232 N_A_27_115#_c_269_n N_Y_c_449_n 0.021445f $X=2.55 $Y=2.405 $X2=2.41
+ $Y2=2.11
cc_233 N_A_27_115#_c_322_n N_Y_c_449_n 0.00375894f $X=2.625 $Y=2.48 $X2=2.41
+ $Y2=2.11
cc_234 N_A_27_115#_c_281_n N_Y_c_449_n 0.00361281f $X=3.055 $Y=2.33 $X2=2.41
+ $Y2=2.11
cc_235 N_A_27_115#_M1014_g N_Y_c_450_n 0.00182852f $X=3.055 $Y=0.835 $X2=3.27
+ $Y2=0.755
cc_236 N_A_27_115#_c_282_n N_Y_c_450_n 0.00274041f $X=3.41 $Y=1.365 $X2=3.27
+ $Y2=0.755
cc_237 N_A_27_115#_M1015_g N_Y_c_450_n 0.00182852f $X=3.485 $Y=0.835 $X2=3.27
+ $Y2=0.755
cc_238 N_A_27_115#_c_281_n N_Y_c_454_n 0.00721971f $X=3.055 $Y=2.33 $X2=3.27
+ $Y2=2.11
cc_239 N_A_27_115#_c_328_n N_Y_c_454_n 0.00375894f $X=3.055 $Y=2.48 $X2=3.27
+ $Y2=2.11
cc_240 N_A_27_115#_c_282_n N_Y_c_454_n 0.00250559f $X=3.41 $Y=1.365 $X2=3.27
+ $Y2=2.11
cc_241 N_A_27_115#_c_283_n N_Y_c_454_n 0.0206674f $X=3.41 $Y=2.405 $X2=3.27
+ $Y2=2.11
cc_242 N_A_27_115#_c_333_n N_Y_c_454_n 0.00375894f $X=3.485 $Y=2.48 $X2=3.27
+ $Y2=2.11
cc_243 N_A_27_115#_M1000_g N_Y_c_455_n 0.00493416f $X=1.335 $Y=0.835 $X2=1.55
+ $Y2=1.115
cc_244 N_A_27_115#_M1009_g N_Y_c_455_n 0.00198614f $X=1.765 $Y=0.835 $X2=1.55
+ $Y2=1.115
cc_245 N_A_27_115#_c_303_n N_Y_c_455_n 0.00238892f $X=1.395 $Y=1.455 $X2=1.55
+ $Y2=1.115
cc_246 N_A_27_115#_c_254_n N_Y_c_459_n 0.00638728f $X=1.335 $Y=2.33 $X2=1.55
+ $Y2=1.995
cc_247 N_A_27_115#_c_255_n N_Y_c_459_n 0.00186325f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=1.995
cc_248 N_A_27_115#_c_256_n N_Y_c_459_n 0.00140336f $X=1.69 $Y=1.365 $X2=1.55
+ $Y2=1.995
cc_249 N_A_27_115#_c_288_n N_Y_c_459_n 0.00144278f $X=1.395 $Y=1.365 $X2=1.55
+ $Y2=1.995
cc_250 N_A_27_115#_c_303_n N_Y_c_459_n 0.00194461f $X=1.395 $Y=1.455 $X2=1.55
+ $Y2=1.995
cc_251 N_A_27_115#_M1000_g Y 0.00251111f $X=1.335 $Y=0.835 $X2=1.555 $Y2=1.74
cc_252 N_A_27_115#_c_254_n Y 0.00874077f $X=1.335 $Y=2.33 $X2=1.555 $Y2=1.74
cc_253 N_A_27_115#_c_256_n Y 0.00840707f $X=1.69 $Y=1.365 $X2=1.555 $Y2=1.74
cc_254 N_A_27_115#_M1009_g Y 0.00251111f $X=1.765 $Y=0.835 $X2=1.555 $Y2=1.74
cc_255 N_A_27_115#_c_288_n Y 0.00487273f $X=1.395 $Y=1.365 $X2=1.555 $Y2=1.74
cc_256 N_A_27_115#_c_303_n Y 0.0132141f $X=1.395 $Y=1.455 $X2=1.555 $Y2=1.74
cc_257 N_A_27_115#_M1009_g N_Y_c_461_n 0.00873177f $X=1.765 $Y=0.835 $X2=2.265
+ $Y2=1
cc_258 N_A_27_115#_c_261_n N_Y_c_461_n 0.00213861f $X=2.12 $Y=1.365 $X2=2.265
+ $Y2=1
cc_259 N_A_27_115#_M1011_g N_Y_c_461_n 0.00873177f $X=2.195 $Y=0.835 $X2=2.265
+ $Y2=1
cc_260 N_A_27_115#_c_290_n N_Y_c_465_n 0.0121767f $X=1.765 $Y=1.365 $X2=2.265
+ $Y2=2.11
cc_261 N_A_27_115#_c_291_n N_Y_c_465_n 0.0158479f $X=1.765 $Y=2.405 $X2=2.265
+ $Y2=2.11
cc_262 N_A_27_115#_M1011_g N_Y_c_466_n 0.00251111f $X=2.195 $Y=0.835 $X2=2.41
+ $Y2=1.995
cc_263 N_A_27_115#_c_268_n N_Y_c_466_n 0.0177725f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=1.995
cc_264 N_A_27_115#_M1013_g N_Y_c_466_n 0.00251111f $X=2.625 $Y=0.835 $X2=2.41
+ $Y2=1.995
cc_265 N_A_27_115#_c_281_n N_Y_c_466_n 0.00843025f $X=3.055 $Y=2.33 $X2=2.41
+ $Y2=1.995
cc_266 N_A_27_115#_M1013_g N_Y_c_467_n 0.00873177f $X=2.625 $Y=0.835 $X2=3.125
+ $Y2=1
cc_267 N_A_27_115#_c_274_n N_Y_c_467_n 0.00213861f $X=2.98 $Y=1.365 $X2=3.125
+ $Y2=1
cc_268 N_A_27_115#_M1014_g N_Y_c_467_n 0.00938169f $X=3.055 $Y=0.835 $X2=3.125
+ $Y2=1
cc_269 N_A_27_115#_M1011_g N_Y_c_471_n 0.00198614f $X=2.195 $Y=0.835 $X2=2.555
+ $Y2=1
cc_270 N_A_27_115#_M1013_g N_Y_c_471_n 0.00198614f $X=2.625 $Y=0.835 $X2=2.555
+ $Y2=1
cc_271 N_A_27_115#_c_281_n N_Y_c_475_n 0.0155956f $X=3.055 $Y=2.33 $X2=3.125
+ $Y2=2.11
cc_272 N_A_27_115#_c_294_n N_Y_c_475_n 0.00894336f $X=2.625 $Y=1.365 $X2=3.125
+ $Y2=2.11
cc_273 N_A_27_115#_c_295_n N_Y_c_475_n 0.00903839f $X=2.625 $Y=2.405 $X2=3.125
+ $Y2=2.11
cc_274 N_A_27_115#_c_268_n N_Y_c_476_n 0.00140336f $X=2.55 $Y=1.365 $X2=2.555
+ $Y2=2.11
cc_275 N_A_27_115#_c_281_n N_Y_c_476_n 0.0012308f $X=3.055 $Y=2.33 $X2=2.555
+ $Y2=2.11
cc_276 N_A_27_115#_c_292_n N_Y_c_476_n 0.00140336f $X=2.195 $Y=1.365 $X2=2.555
+ $Y2=2.11
cc_277 N_A_27_115#_c_293_n N_Y_c_476_n 0.00372651f $X=2.195 $Y=2.405 $X2=2.555
+ $Y2=2.11
cc_278 N_A_27_115#_M1014_g N_Y_c_477_n 0.00201073f $X=3.055 $Y=0.835 $X2=3.27
+ $Y2=1.115
cc_279 N_A_27_115#_M1015_g N_Y_c_477_n 0.00878256f $X=3.485 $Y=0.835 $X2=3.27
+ $Y2=1.115
cc_280 N_A_27_115#_M1014_g N_Y_c_481_n 0.00251111f $X=3.055 $Y=0.835 $X2=3.27
+ $Y2=1.995
cc_281 N_A_27_115#_c_281_n N_Y_c_481_n 0.0163934f $X=3.055 $Y=2.33 $X2=3.27
+ $Y2=1.995
cc_282 N_A_27_115#_c_282_n N_Y_c_481_n 0.0196907f $X=3.41 $Y=1.365 $X2=3.27
+ $Y2=1.995
cc_283 N_A_27_115#_c_283_n N_Y_c_481_n 0.00357274f $X=3.41 $Y=2.405 $X2=3.27
+ $Y2=1.995
cc_284 N_A_27_115#_M1015_g N_Y_c_481_n 0.00251111f $X=3.485 $Y=0.835 $X2=3.27
+ $Y2=1.995
