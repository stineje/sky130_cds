* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_12T_hs__dffr_1
** N=28 EP=0 IP=0 FDC=38
M0 4 RN gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=400 $Y=575 $D=19
M1 8 4 gnd gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1350 $Y=575 $D=19
M2 gnd 5 8 gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1780 $Y=575 $D=19
M3 20 D gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=2730 $Y=575 $D=19
M4 5 9 20 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=3090 $Y=575 $D=19
M5 21 CK 5 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=3690 $Y=575 $D=19
M6 gnd 8 21 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=4050 $Y=575 $D=19
M7 22 8 gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=4480 $Y=575 $D=19
M8 11 CK 22 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=4840 $Y=575 $D=19
M9 23 9 11 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=5440 $Y=575 $D=19
M10 gnd 10 23 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=5800 $Y=575 $D=19
M11 9 CK gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=6230 $Y=575 $D=19
M12 10 11 gnd gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7180 $Y=575 $D=19
M13 gnd 4 10 gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7610 $Y=575 $D=19
M14 gnd 10 QN gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=8560 $Y=575 $D=19
M15 Q QN gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=8990 $Y=575 $D=19
M16 4 RN vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=400 $Y=2605 $D=79
M17 13 4 8 vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=1350 $Y=3025 $D=79
M18 vdd 5 13 vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=1710 $Y=3025 $D=79
M19 14 D vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=2730 $Y=2605 $D=79
M20 5 CK 14 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=3090 $Y=2605 $D=79
M21 15 9 5 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=3690 $Y=2605 $D=79
M22 vdd 8 15 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=4050 $Y=2605 $D=79
M23 16 8 vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=4480 $Y=2605 $D=79
M24 11 9 16 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=4840 $Y=2605 $D=79
M25 17 CK 11 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=5440 $Y=2605 $D=79
M26 vdd 10 17 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=5800 $Y=2605 $D=79
M27 9 CK vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=6230 $Y=2605 $D=79
M28 18 11 10 vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=7180 $Y=3025 $D=79
M29 vdd 4 18 vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=7540 $Y=3025 $D=79
M30 vdd 10 QN vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=8560 $Y=2605 $D=79
M31 Q QN vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=8990 $Y=2605 $D=79
X32 gnd vdd Dpar a=19.8481 p=23.39 m=1 $[nwdiode] $X=-50 $Y=2425 $D=185
X33 24 RN Probe probetype=1 $[RN] $X=323 $Y=2848 $D=289
X34 25 D Probe probetype=1 $[D] $X=2863 $Y=1738 $D=289
X35 26 CK Probe probetype=1 $[CK] $X=6448 $Y=2108 $D=289
X36 27 QN Probe probetype=1 $[QN] $X=8423 $Y=2478 $D=289
X37 28 Q Probe probetype=1 $[Q] $X=9273 $Y=2848 $D=289
.ENDS
***************************************
