* File: sky130_osu_sc_12T_ms__dffnr_1.pex.spice
* Created: Fri Feb 12 20:30:12 2021
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%GND 1 2 3 4 5 6 7 8 9 84 88 90 97 99
+ 106 108 115 117 127 129 139 141 148 150 157 159 166 185 187
c248 157 0 5.73867e-20 $X=7.9 $Y=0.74
c249 139 0 1.71621e-19 $X=6.09 $Y=0.755
c250 115 0 3.07651e-19 $X=2.59 $Y=0.755
c251 97 0 5.44281e-20 $X=1.21 $Y=0.74
c252 84 0 1.61973e-19 $X=-0.05 $Y=0
r253 185 187 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.175 $Y2=0.152
r254 179 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.152
+ $X2=8.85 $Y2=0.152
r255 164 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.152
r256 164 166 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.74
r257 159 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.152
+ $X2=8.85 $Y2=0.152
r258 155 157 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.74
r259 151 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.152
+ $X2=7.04 $Y2=0.152
r260 146 175 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.152
r261 146 148 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.74
r262 142 174 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.152
+ $X2=6.09 $Y2=0.152
r263 141 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.152
+ $X2=7.04 $Y2=0.152
r264 137 174 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.152
r265 137 139 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.755
r266 129 174 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.152
+ $X2=6.09 $Y2=0.152
r267 125 127 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.34 $Y=0.305
+ $X2=4.34 $Y2=0.74
r268 118 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.152
+ $X2=2.59 $Y2=0.152
r269 113 170 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.152
r270 113 115 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.755
r271 109 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.152
+ $X2=2.07 $Y2=0.152
r272 108 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.152
+ $X2=2.59 $Y2=0.152
r273 104 169 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.152
r274 104 106 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.74
r275 100 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.152
+ $X2=1.21 $Y2=0.152
r276 99 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.152
+ $X2=2.07 $Y2=0.152
r277 95 168 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.152
r278 95 97 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.74
r279 90 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.152
+ $X2=1.21 $Y2=0.152
r280 86 88 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r281 84 86 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r282 84 91 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r283 84 179 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.935 $Y2=0.152
r284 84 187 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175 $Y=0.19
+ $X2=9.175 $Y2=0.19
r285 84 185 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r286 84 155 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r287 84 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r288 84 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.985 $Y2=0.152
r289 84 125 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.34 $Y2=0.305
r290 84 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.255 $Y2=0.152
r291 84 130 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.425 $Y2=0.152
r292 84 159 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.765 $Y2=0.152
r293 84 160 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=7.985 $Y2=0.152
r294 84 150 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r295 84 151 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.125 $Y2=0.152
r296 84 141 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.955 $Y2=0.152
r297 84 142 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.175 $Y2=0.152
r298 84 129 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.005 $Y2=0.152
r299 84 130 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.425 $Y2=0.152
r300 84 117 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=4.255 $Y2=0.152
r301 84 118 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=2.675 $Y2=0.152
r302 84 108 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.505 $Y2=0.152
r303 84 109 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.155 $Y2=0.152
r304 84 99 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.985 $Y2=0.152
r305 84 100 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.295 $Y2=0.152
r306 84 90 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.125 $Y2=0.152
r307 84 91 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r308 9 166 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.575 $X2=8.85 $Y2=0.74
r309 8 157 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.74
r310 7 148 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.575 $X2=7.04 $Y2=0.74
r311 6 139 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.575 $X2=6.09 $Y2=0.755
r312 5 127 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.575 $X2=4.34 $Y2=0.74
r313 4 115 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.575 $X2=2.59 $Y2=0.755
r314 3 106 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.74
r315 2 97 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.74
r316 1 88 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%VDD 1 2 3 4 5 6 7 64 68 70 78 86 88 96
+ 98 106 108 116 118 124 136 141 145
c124 124 0 1.98165e-19 $X=8.85 $Y=3.265
r125 141 145 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=4.25 $X2=9.175 $Y2=4.25
r126 136 141 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=4.287
+ $X2=9.175 $Y2=4.287
r127 136 139 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=4.25 $X2=0.335 $Y2=4.25
r128 133 145 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=8.935 $Y=4.287
+ $X2=9.175 $Y2=4.287
r129 133 134 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=4.287
+ $X2=8.85 $Y2=4.287
r130 122 134 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.85 $Y=4.135
+ $X2=8.85 $Y2=4.287
r131 122 124 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.85 $Y=4.135
+ $X2=8.85 $Y2=3.265
r132 119 132 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=4.287
+ $X2=7.83 $Y2=4.287
r133 119 121 21.9153 $w=3.03e-07 $l=5.8e-07 $layer=LI1_cond $X=7.915 $Y=4.287
+ $X2=8.495 $Y2=4.287
r134 118 134 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=4.287
+ $X2=8.85 $Y2=4.287
r135 118 121 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.765 $Y=4.287
+ $X2=8.495 $Y2=4.287
r136 114 132 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.83 $Y=4.135
+ $X2=7.83 $Y2=4.287
r137 114 116 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=7.83 $Y=4.135
+ $X2=7.83 $Y2=3.275
r138 111 113 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.455 $Y=4.287
+ $X2=7.135 $Y2=4.287
r139 109 130 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.09 $Y2=4.287
r140 109 111 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.455 $Y2=4.287
r141 108 132 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=4.287
+ $X2=7.83 $Y2=4.287
r142 108 113 23.0489 $w=3.03e-07 $l=6.1e-07 $layer=LI1_cond $X=7.745 $Y=4.287
+ $X2=7.135 $Y2=4.287
r143 104 130 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=4.287
r144 104 106 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=3.21
r145 101 103 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=4.287
+ $X2=5.775 $Y2=4.287
r146 99 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=4.287
+ $X2=4.34 $Y2=4.287
r147 99 101 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.425 $Y=4.287
+ $X2=5.095 $Y2=4.287
r148 98 130 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=6.09 $Y2=4.287
r149 98 103 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=5.775 $Y2=4.287
r150 94 129 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.34 $Y=4.135
+ $X2=4.34 $Y2=4.287
r151 94 96 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.34 $Y=4.135
+ $X2=4.34 $Y2=3.295
r152 91 93 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=4.287
+ $X2=3.735 $Y2=4.287
r153 89 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=4.287
+ $X2=2.59 $Y2=4.287
r154 89 91 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.675 $Y=4.287
+ $X2=3.055 $Y2=4.287
r155 88 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=4.287
+ $X2=4.34 $Y2=4.287
r156 88 93 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=4.255 $Y=4.287
+ $X2=3.735 $Y2=4.287
r157 84 127 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.59 $Y=4.135
+ $X2=2.59 $Y2=4.287
r158 84 86 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.59 $Y=4.135
+ $X2=2.59 $Y2=3.295
r159 81 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=4.287
+ $X2=2 $Y2=4.287
r160 81 83 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=2.085 $Y=4.287
+ $X2=2.375 $Y2=4.287
r161 80 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=4.287
+ $X2=2.59 $Y2=4.287
r162 80 83 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=4.287
+ $X2=2.375 $Y2=4.287
r163 76 126 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2 $Y=4.135 $X2=2
+ $Y2=4.287
r164 76 78 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2 $Y=4.135 $X2=2
+ $Y2=3.275
r165 73 75 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=4.287
+ $X2=1.695 $Y2=4.287
r166 71 139 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r167 71 73 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.015 $Y2=4.287
r168 70 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=4.287
+ $X2=2 $Y2=4.287
r169 70 75 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.915 $Y=4.287
+ $X2=1.695 $Y2=4.287
r170 66 139 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r171 66 68 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r172 64 139 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=4.135 $X2=0.335 $Y2=4.22
r173 64 145 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=4.135 $X2=9.175 $Y2=4.22
r174 64 132 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=4.135 $X2=7.815 $Y2=4.22
r175 64 129 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=4.135 $X2=4.415 $Y2=4.22
r176 64 121 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=4.135 $X2=8.495 $Y2=4.22
r177 64 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=4.135 $X2=7.135 $Y2=4.22
r178 64 111 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=4.135 $X2=6.455 $Y2=4.22
r179 64 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=4.135 $X2=5.775 $Y2=4.22
r180 64 101 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=4.135 $X2=5.095 $Y2=4.22
r181 64 93 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=4.135 $X2=3.735 $Y2=4.22
r182 64 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=4.135 $X2=3.055 $Y2=4.22
r183 64 83 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=4.135 $X2=2.375 $Y2=4.22
r184 64 75 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=4.135 $X2=1.695 $Y2=4.22
r185 64 73 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=4.135 $X2=1.015 $Y2=4.22
r186 7 124 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=2.605 $X2=8.85 $Y2=3.265
r187 6 116 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=3.025 $X2=7.83 $Y2=3.275
r188 5 106 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=5.95
+ $Y=2.605 $X2=6.09 $Y2=3.21
r189 4 96 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=2.605 $X2=4.34 $Y2=3.295
r190 3 86 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.605 $X2=2.59 $Y2=3.295
r191 2 78 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=3.025 $X2=2 $Y2=3.275
r192 1 68 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%RN 3 5 7 9 16 17
c38 17 0 7.50258e-20 $X=0.325 $Y=2.85
r39 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.825 $X2=0.53 $Y2=1.825
r41 10 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=1.99 $X2=0.32
+ $Y2=2.85
r42 9 12 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.53 $Y2=1.825
r43 9 10 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.32 $Y2=1.99
r44 5 13 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.53 $Y2=1.825
r45 5 7 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=3.235
r46 1 13 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.53 $Y2=1.825
r47 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%A_110_115# 1 2 7 9 12 14 16 18 20 23 27
+ 32 33 34 39 42 43 44 46 48 52 57 59 63
c198 52 0 5.73867e-20 $X=7.89 $Y=1.37
c199 48 0 5.44281e-20 $X=1.22 $Y=1.37
c200 39 0 7.50258e-20 $X=0.87 $Y=2.26
c201 14 0 1.71863e-19 $X=7.615 $Y=1.52
r202 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.21 $X2=7.89 $Y2=1.21
r203 56 59 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.22 $Y=1.21
+ $X2=1.425 $Y2=1.21
r204 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.21 $X2=1.22 $Y2=1.21
r205 52 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.89 $Y=1.37
+ $X2=7.89 $Y2=1.37
r206 48 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.22 $Y=1.37
+ $X2=1.22 $Y2=1.37
r207 46 52 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=7.89 $Y=1.255
+ $X2=7.89 $Y2=1.37
r208 45 46 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=7.89 $Y=1.085
+ $X2=7.89 $Y2=1.255
r209 43 45 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=7.805 $Y=1
+ $X2=7.89 $Y2=1.085
r210 43 44 6.25874 $w=1.7e-07 $l=6.5e-06 $layer=MET1_cond $X=7.805 $Y=1
+ $X2=1.305 $Y2=1
r211 42 48 0.0829981 $w=2.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.22 $Y=1.255
+ $X2=1.22 $Y2=1.37
r212 41 44 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.22 $Y=1.085
+ $X2=1.305 $Y2=1
r213 41 42 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.22 $Y=1.085
+ $X2=1.22 $Y2=1.255
r214 37 39 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.26
+ $X2=0.87 $Y2=2.26
r215 35 36 10.0734 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.87 $Y2=1.16
r216 34 36 5.3812 $w=2.18e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.955 $Y=1.21
+ $X2=0.87 $Y2=1.16
r217 33 57 2.00497 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.135 $Y=1.21
+ $X2=1.26 $Y2=1.21
r218 33 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.135 $Y=1.21
+ $X2=0.955 $Y2=1.21
r219 32 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=2.26
r220 31 36 2.19618 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.16
r221 31 32 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=2.175
r222 27 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.95
+ $X2=0.69 $Y2=3.63
r223 25 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.26
r224 25 27 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.95
r225 21 35 2.19618 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=1.16
r226 21 23 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=0.755
r227 18 62 38.8445 $w=3.55e-07 $l=2.07918e-07 $layer=POLY_cond $X=7.685 $Y=1.045
+ $X2=7.782 $Y2=1.21
r228 18 20 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.685 $Y=1.045
+ $X2=7.685 $Y2=0.755
r229 14 62 58.5319 $w=3.55e-07 $l=3.84539e-07 $layer=POLY_cond $X=7.615 $Y=1.52
+ $X2=7.782 $Y2=1.21
r230 14 16 987.074 $w=1.5e-07 $l=1.925e-06 $layer=POLY_cond $X=7.615 $Y=1.52
+ $X2=7.615 $Y2=3.445
r231 10 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.375
+ $X2=1.425 $Y2=1.21
r232 10 12 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=1.425 $Y=1.375
+ $X2=1.425 $Y2=3.445
r233 7 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.045
+ $X2=1.425 $Y2=1.21
r234 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.425 $Y=1.045
+ $X2=1.425 $Y2=0.755
r235 2 29 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.63
r236 2 27 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.95
r237 1 23 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%A_342_442# 1 2 9 13 16 17 19 20 22 25
+ 30 31 33
c83 33 0 1.72079e-19 $X=3.365 $Y=0.755
c84 19 0 1.29912e-19 $X=3.28 $Y=1.285
r85 33 35 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=3.365 $Y=0.755
+ $X2=3.465 $Y2=0.755
r86 31 38 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.375
+ $X2=1.892 $Y2=2.54
r87 31 37 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.375
+ $X2=1.892 $Y2=2.21
r88 30 32 15.1353 $w=2.66e-07 $l=3.3e-07 $layer=LI1_cond $X=2.025 $Y=2.375
+ $X2=2.025 $Y2=2.705
r89 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.375 $X2=1.94 $Y2=2.375
r90 25 27 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=3.465 $Y=2.955
+ $X2=3.465 $Y2=3.635
r91 23 25 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=2.79
+ $X2=3.465 $Y2=2.955
r92 21 33 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.365 $Y=0.935
+ $X2=3.365 $Y2=0.755
r93 21 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=0.935
+ $X2=3.365 $Y2=1.2
r94 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=1.285
+ $X2=3.365 $Y2=1.2
r95 19 20 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.28 $Y=1.285
+ $X2=2.2 $Y2=1.285
r96 18 32 3.35683 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.195 $Y=2.705
+ $X2=2.025 $Y2=2.705
r97 17 23 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.295 $Y=2.705
+ $X2=3.465 $Y2=2.79
r98 17 18 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.295 $Y=2.705
+ $X2=2.195 $Y2=2.705
r99 16 30 9.15133 $w=2.66e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.11 $Y=2.21
+ $X2=2.025 $Y2=2.375
r100 15 20 6.81649 $w=1.7e-07 $l=2.25555e-07 $layer=LI1_cond $X=2.11 $Y=1.47
+ $X2=2.2 $Y2=1.285
r101 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.11 $Y=1.47
+ $X2=2.11 $Y2=2.21
r102 13 37 746.074 $w=1.5e-07 $l=1.455e-06 $layer=POLY_cond $X=1.855 $Y=0.755
+ $X2=1.855 $Y2=2.21
r103 9 38 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.785 $Y=3.445
+ $X2=1.785 $Y2=2.54
r104 2 27 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.605 $X2=3.465 $Y2=3.635
r105 2 25 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.605 $X2=3.465 $Y2=2.955
r106 1 35 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.575 $X2=3.465 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%D 3 7 10 13 15
c42 15 0 1.12321e-19 $X=2.865 $Y=1.74
c43 10 0 1.41836e-19 $X=2.865 $Y=1.74
r44 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.905
r45 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.575
r46 13 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.74 $X2=2.865 $Y2=1.74
r47 10 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.74
r48 7 18 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=2.805 $Y=3.235
+ $X2=2.805 $Y2=1.905
r49 3 17 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.805 $Y=0.835
+ $X2=2.805 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%A_618_424# 1 2 9 13 16 19 21 25 26 30
+ 31 33 34 37 42 43 44 48 52 56 57 58 59 62 66 68 69 72 77 80 83
c258 83 0 4.72879e-20 $X=5.455 $Y=2.285
c259 77 0 1.29912e-19 $X=3.705 $Y=1.205
c260 72 0 1.41836e-19 $X=3.225 $Y=2.285
c261 68 0 1.59924e-19 $X=6.87 $Y=2.11
c262 56 0 1.89675e-19 $X=5.31 $Y=2.11
c263 34 0 6.79641e-20 $X=5.06 $Y=2.11
c264 33 0 1.70195e-19 $X=5.37 $Y=2.11
c265 25 0 1.98654e-19 $X=3.705 $Y=1.37
c266 21 0 1.86602e-19 $X=3.62 $Y=2.11
r267 83 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=2.285
+ $X2=5.455 $Y2=2.45
r268 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=2.285 $X2=5.455 $Y2=2.285
r269 72 75 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.285
+ $X2=3.225 $Y2=2.45
r270 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=2.285 $X2=3.225 $Y2=2.285
r271 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.87 $Y=2.11
+ $X2=6.87 $Y2=2.11
r272 66 84 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.455 $Y=2.11
+ $X2=5.455 $Y2=2.285
r273 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=2.11
+ $X2=5.455 $Y2=2.11
r274 62 73 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.225 $Y=2.11
+ $X2=3.225 $Y2=2.285
r275 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.225 $Y=2.11
+ $X2=3.225 $Y2=2.11
r276 59 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=2.11
+ $X2=5.455 $Y2=2.11
r277 58 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.725 $Y=2.11
+ $X2=6.87 $Y2=2.11
r278 58 59 1.08324 $w=1.7e-07 $l=1.125e-06 $layer=MET1_cond $X=6.725 $Y=2.11
+ $X2=5.6 $Y2=2.11
r279 57 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.37 $Y=2.11
+ $X2=3.225 $Y2=2.11
r280 56 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.31 $Y=2.11
+ $X2=5.455 $Y2=2.11
r281 56 57 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.31 $Y=2.11
+ $X2=3.37 $Y2=2.11
r282 55 69 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.87 $Y=2.62
+ $X2=6.87 $Y2=2.11
r283 53 69 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.87 $Y=1.93
+ $X2=6.87 $Y2=2.11
r284 52 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.87 $Y=1.845
+ $X2=6.87 $Y2=1.93
r285 50 52 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.69 $Y=1.845
+ $X2=6.87 $Y2=1.845
r286 46 48 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=0.755
+ $X2=6.69 $Y2=0.755
r287 43 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.705
+ $X2=6.87 $Y2=2.62
r288 43 44 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.785 $Y=2.705
+ $X2=6.605 $Y2=2.705
r289 42 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.69 $Y=1.76
+ $X2=6.69 $Y2=1.845
r290 41 48 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.69 $Y=0.855 $X2=6.69
+ $Y2=0.755
r291 41 42 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.69 $Y=0.855
+ $X2=6.69 $Y2=1.76
r292 37 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.52 $Y=2.955
+ $X2=6.52 $Y2=3.635
r293 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.52 $Y=2.79
+ $X2=6.605 $Y2=2.705
r294 35 37 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=2.79
+ $X2=6.52 $Y2=2.955
r295 33 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.11
+ $X2=5.455 $Y2=2.11
r296 33 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.37 $Y=2.11
+ $X2=5.06 $Y2=2.11
r297 31 80 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.37
+ $X2=4.975 $Y2=1.205
r298 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.37 $X2=4.975 $Y2=1.37
r299 28 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=2.025
+ $X2=5.06 $Y2=2.11
r300 28 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.975 $Y=2.025
+ $X2=4.975 $Y2=1.37
r301 26 77 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.37
+ $X2=3.705 $Y2=1.205
r302 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.37 $X2=3.705 $Y2=1.37
r303 23 25 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.705 $Y=2.025
+ $X2=3.705 $Y2=1.37
r304 22 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.11
+ $X2=3.225 $Y2=2.11
r305 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.11
+ $X2=3.705 $Y2=2.025
r306 21 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.62 $Y=2.11
+ $X2=3.31 $Y2=2.11
r307 19 86 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.515 $Y=3.235
+ $X2=5.515 $Y2=2.45
r308 16 80 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.915 $Y=0.835
+ $X2=4.915 $Y2=1.205
r309 13 77 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.765 $Y=0.835
+ $X2=3.765 $Y2=1.205
r310 9 75 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.165 $Y=3.235
+ $X2=3.165 $Y2=2.45
r311 2 39 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=3.635
r312 2 37 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=2.955
r313 1 46 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%A_217_605# 1 2 9 13 17 21 23 24 25 26
+ 29 31 32 35 39 45 47 48 55
c138 39 0 1.35571e-19 $X=4.06 $Y=1.37
c139 35 0 1.5821e-19 $X=4.295 $Y=2.285
c140 26 0 6.79641e-20 $X=4.48 $Y=2.285
c141 24 0 1.86602e-19 $X=4.2 $Y=2.285
c142 21 0 6.36774e-20 $X=4.555 $Y=3.235
c143 13 0 6.36774e-20 $X=4.125 $Y=3.235
r144 48 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.37 $X2=4.295 $Y2=1.37
r145 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=1.37
+ $X2=4.205 $Y2=1.37
r146 43 55 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.64 $Y=1.37
+ $X2=1.64 $Y2=0.74
r147 42 45 0.0982977 $w=2.45e-07 $l=1.4e-07 $layer=MET1_cond $X=1.64 $Y=1.372
+ $X2=1.78 $Y2=1.372
r148 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.37
+ $X2=1.64 $Y2=1.37
r149 39 47 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.37
+ $X2=4.205 $Y2=1.37
r150 39 45 2.19537 $w=1.7e-07 $l=2.28e-06 $layer=MET1_cond $X=4.06 $Y=1.37
+ $X2=1.78 $Y2=1.37
r151 38 43 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.64 $Y=1.725
+ $X2=1.64 $Y2=1.37
r152 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=2.285 $X2=4.295 $Y2=2.285
r153 33 48 2.3025 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.295 $Y=1.455
+ $X2=4.205 $Y2=1.33
r154 33 35 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.295 $Y=1.455
+ $X2=4.295 $Y2=2.285
r155 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.64 $Y2=1.725
r156 31 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.295 $Y2=1.81
r157 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.895
+ $X2=1.295 $Y2=1.81
r158 27 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.21 $Y=1.895
+ $X2=1.21 $Y2=3.275
r159 26 36 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=2.285
+ $X2=4.295 $Y2=2.285
r160 25 51 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=1.37
+ $X2=4.295 $Y2=1.37
r161 24 36 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=2.285
+ $X2=4.295 $Y2=2.285
r162 23 51 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=1.37
+ $X2=4.295 $Y2=1.37
r163 19 26 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.48 $Y2=2.285
r164 19 21 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.555 $Y2=3.235
r165 15 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.235
+ $X2=4.48 $Y2=1.37
r166 15 17 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.555 $Y=1.235
+ $X2=4.555 $Y2=0.835
r167 11 24 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=2.42
+ $X2=4.2 $Y2=2.285
r168 11 13 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.125 $Y=2.42
+ $X2=4.125 $Y2=3.235
r169 7 23 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=1.235
+ $X2=4.2 $Y2=1.37
r170 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.125 $Y=1.235
+ $X2=4.125 $Y2=0.835
r171 2 29 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=3.025 $X2=1.21 $Y2=3.275
r172 1 55 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%CK 1 3 5 6 7 10 12 16 18 22 24 26 27 29
+ 32 35 37 38 41 47 50 51 58 59 63 64
c204 64 0 1.89675e-19 $X=5.455 $Y=1.725
c205 58 0 7.96265e-20 $X=6.305 $Y=1.74
c206 51 0 4.36612e-19 $X=5.6 $Y=1.74
c207 50 0 2.9867e-19 $X=6.16 $Y=1.74
c208 35 0 1.98654e-19 $X=3.285 $Y=1.28
c209 10 0 1.12321e-19 $X=3.765 $Y=3.235
r210 63 66 18.9959 $w=3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.47 $Y=1.725
+ $X2=5.47 $Y2=1.82
r211 63 65 55.9777 $w=3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.47 $Y=1.725
+ $X2=5.47 $Y2=1.52
r212 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.725 $X2=5.455 $Y2=1.725
r213 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.305 $Y=1.74
+ $X2=6.305 $Y2=1.74
r214 53 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=1.74
+ $X2=5.455 $Y2=1.74
r215 51 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=1.74
+ $X2=5.455 $Y2=1.74
r216 50 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.16 $Y=1.74
+ $X2=6.305 $Y2=1.74
r217 50 51 0.539214 $w=1.7e-07 $l=5.6e-07 $layer=MET1_cond $X=6.16 $Y=1.74
+ $X2=5.6 $Y2=1.74
r218 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=2.285 $X2=6.45 $Y2=2.285
r219 44 58 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.305 $Y=2.12
+ $X2=6.305 $Y2=1.74
r220 43 47 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.305 $Y=2.285
+ $X2=6.45 $Y2=2.285
r221 43 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=2.285
+ $X2=6.305 $Y2=2.12
r222 39 41 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=6.305 $Y=1.28
+ $X2=6.385 $Y2=1.28
r223 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.165 $Y=1.28
+ $X2=3.285 $Y2=1.28
r224 32 48 38.571 $w=3.25e-07 $l=1.75656e-07 $layer=POLY_cond $X=6.385 $Y=2.12
+ $X2=6.407 $Y2=2.285
r225 31 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.385 $Y=1.355
+ $X2=6.385 $Y2=1.28
r226 31 32 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.385 $Y=1.355
+ $X2=6.385 $Y2=2.12
r227 27 48 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.305 $Y=2.45
+ $X2=6.407 $Y2=2.285
r228 27 29 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.305 $Y=2.45
+ $X2=6.305 $Y2=3.235
r229 24 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=1.28
r230 24 26 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=0.835
r231 22 65 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=5.515 $Y=0.835
+ $X2=5.515 $Y2=1.52
r232 19 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.99 $Y=1.82
+ $X2=4.915 $Y2=1.82
r233 18 66 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.32 $Y=1.82
+ $X2=5.47 $Y2=1.82
r234 18 19 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.32 $Y=1.82
+ $X2=4.99 $Y2=1.82
r235 14 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.915 $Y=1.895
+ $X2=4.915 $Y2=1.82
r236 14 16 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=4.915 $Y=1.895
+ $X2=4.915 $Y2=3.235
r237 13 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.82
+ $X2=3.765 $Y2=1.82
r238 12 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=1.82
+ $X2=4.915 $Y2=1.82
r239 12 13 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.84 $Y=1.82 $X2=3.84
+ $Y2=1.82
r240 8 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.895
+ $X2=3.765 $Y2=1.82
r241 8 10 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=3.765 $Y=1.895
+ $X2=3.765 $Y2=3.235
r242 6 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=1.82
+ $X2=3.765 $Y2=1.82
r243 6 7 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.69 $Y=1.82 $X2=3.36
+ $Y2=1.82
r244 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.285 $Y=1.745
+ $X2=3.36 $Y2=1.82
r245 4 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.355
+ $X2=3.285 $Y2=1.28
r246 4 5 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.285 $Y=1.355
+ $X2=3.285 $Y2=1.745
r247 1 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.205
+ $X2=3.165 $Y2=1.28
r248 1 3 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.165 $Y=1.205
+ $X2=3.165 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%A_1160_89# 1 2 9 12 24 27 28 29 30 31
+ 32 33 34 35 38 40 41 44 47 48 51 53 54 55 57 59 62 65 66 67 70 73 75
c208 73 0 2.20611e-19 $X=8.52 $Y=1.74
c209 70 0 1.31857e-19 $X=5.965 $Y=1.605
c210 54 0 7.96265e-20 $X=7.155 $Y=2.48
c211 51 0 9.09695e-20 $X=5.965 $Y=1.77
c212 34 0 8.77106e-20 $X=8.61 $Y=2.375
c213 31 0 1.50225e-19 $X=5.89 $Y=2.255
c214 29 0 2.82071e-19 $X=5.89 $Y=1.365
r215 73 76 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.74
+ $X2=8.522 $Y2=1.905
r216 73 75 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.74
+ $X2=8.522 $Y2=1.575
r217 66 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.52
+ $Y=1.74 $X2=8.52 $Y2=1.74
r218 65 67 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.52 $Y=1.74
+ $X2=8.375 $Y2=1.74
r219 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.52 $Y=1.74
+ $X2=8.52 $Y2=1.74
r220 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.935 $Y=2.48
+ $X2=5.935 $Y2=2.48
r221 59 67 0.941289 $w=1.75e-07 $l=1.04e-06 $layer=MET1_cond $X=7.335 $Y=1.737
+ $X2=8.375 $Y2=1.737
r222 56 59 0.0698591 $w=1.75e-07 $l=1.2657e-07 $layer=MET1_cond $X=7.245
+ $Y=1.825 $X2=7.335 $Y2=1.737
r223 56 57 0.501568 $w=1.8e-07 $l=5.7e-07 $layer=MET1_cond $X=7.245 $Y=1.825
+ $X2=7.245 $Y2=2.395
r224 55 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=2.48
+ $X2=5.935 $Y2=2.48
r225 54 57 0.0699153 $w=1.7e-07 $l=1.25499e-07 $layer=MET1_cond $X=7.155 $Y=2.48
+ $X2=7.245 $Y2=2.395
r226 54 55 1.0351 $w=1.7e-07 $l=1.075e-06 $layer=MET1_cond $X=7.155 $Y=2.48
+ $X2=6.08 $Y2=2.48
r227 52 66 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.555 $Y=1.74
+ $X2=8.52 $Y2=1.74
r228 52 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=1.74
+ $X2=7.47 $Y2=1.74
r229 51 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=1.77
+ $X2=5.965 $Y2=1.935
r230 51 70 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=1.77
+ $X2=5.965 $Y2=1.605
r231 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.965
+ $Y=1.77 $X2=5.965 $Y2=1.77
r232 48 62 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.935 $Y=2.025
+ $X2=5.935 $Y2=2.48
r233 48 50 17.1635 $w=1.82e-07 $l=2.62393e-07 $layer=LI1_cond $X=5.935 $Y=2.025
+ $X2=5.95 $Y2=1.77
r234 46 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.825
+ $X2=7.47 $Y2=1.74
r235 46 47 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=7.47 $Y=1.825
+ $X2=7.47 $Y2=2.96
r236 42 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.655
+ $X2=7.47 $Y2=1.74
r237 42 44 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.47 $Y=1.655
+ $X2=7.47 $Y2=0.74
r238 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=3.045
+ $X2=7.47 $Y2=2.96
r239 40 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.385 $Y=3.045
+ $X2=7.125 $Y2=3.045
r240 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=3.13
+ $X2=7.125 $Y2=3.045
r241 36 38 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.04 $Y=3.13
+ $X2=7.04 $Y2=3.275
r242 34 35 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=2.375
+ $X2=8.61 $Y2=2.525
r243 34 76 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=8.585 $Y=2.375
+ $X2=8.585 $Y2=1.905
r244 33 75 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.585 $Y=1.32
+ $X2=8.585 $Y2=1.575
r245 32 33 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=1.17 $X2=8.61
+ $Y2=1.32
r246 30 31 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.89 $Y=2.105
+ $X2=5.89 $Y2=2.255
r247 30 71 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.905 $Y=2.105
+ $X2=5.905 $Y2=1.935
r248 29 70 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.905 $Y=1.365
+ $X2=5.905 $Y2=1.605
r249 28 29 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=5.89 $Y=1.205
+ $X2=5.89 $Y2=1.365
r250 27 35 228.147 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=8.635 $Y=3.235
+ $X2=8.635 $Y2=2.525
r251 24 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.635 $Y=0.835
+ $X2=8.635 $Y2=1.17
r252 12 31 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=5.875 $Y=3.235
+ $X2=5.875 $Y2=2.255
r253 9 28 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.875 $Y=0.835
+ $X2=5.875 $Y2=1.205
r254 2 38 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=3.025 $X2=7.04 $Y2=3.275
r255 1 44 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.575 $X2=7.47 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%A_998_115# 1 2 9 13 15 16 19 24 27 28
+ 29 30 33 37 39 40 46
c147 46 0 1.59924e-19 $X=7.255 $Y=1.37
c148 40 0 1.71863e-19 $X=7.05 $Y=1.37
c149 37 0 9.35412e-20 $X=5.315 $Y=1.37
c150 33 0 1.57671e-19 $X=4.635 $Y=1.37
c151 30 0 2.65484e-19 $X=5.44 $Y=1.37
c152 28 0 1.5821e-19 $X=4.78 $Y=1.37
c153 24 0 1.71621e-19 $X=5.215 $Y=0.755
r154 43 46 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=7.05 $Y=1.37
+ $X2=7.255 $Y2=1.37
r155 40 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.05
+ $Y=1.37 $X2=7.05 $Y2=1.37
r156 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.05 $Y=1.37
+ $X2=7.05 $Y2=1.37
r157 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=1.37
+ $X2=5.315 $Y2=1.37
r158 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.37
+ $X2=4.635 $Y2=1.37
r159 30 36 0.0905432 $w=2.3e-07 $l=1.25e-07 $layer=MET1_cond $X=5.44 $Y=1.37
+ $X2=5.315 $Y2=1.37
r160 29 39 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.905 $Y=1.37
+ $X2=7.05 $Y2=1.37
r161 29 30 1.41062 $w=1.7e-07 $l=1.465e-06 $layer=MET1_cond $X=6.905 $Y=1.37
+ $X2=5.44 $Y2=1.37
r162 28 32 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.78 $Y=1.37
+ $X2=4.635 $Y2=1.37
r163 27 36 0.0969593 $w=2.3e-07 $l=1.35e-07 $layer=MET1_cond $X=5.18 $Y=1.37
+ $X2=5.315 $Y2=1.37
r164 27 28 0.385153 $w=1.7e-07 $l=4e-07 $layer=MET1_cond $X=5.18 $Y=1.37
+ $X2=4.78 $Y2=1.37
r165 26 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.315 $Y=1.035
+ $X2=5.315 $Y2=1.37
r166 24 26 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=5.222 $Y=0.755
+ $X2=5.222 $Y2=1.035
r167 21 33 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.635 $Y=2.62
+ $X2=4.635 $Y2=1.37
r168 17 19 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=5.215 $Y=2.79
+ $X2=5.215 $Y2=3.295
r169 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.72 $Y=2.705
+ $X2=4.635 $Y2=2.62
r170 15 17 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=2.705
+ $X2=5.215 $Y2=2.79
r171 15 16 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=2.705
+ $X2=4.72 $Y2=2.705
r172 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.255 $Y=1.535
+ $X2=7.255 $Y2=1.37
r173 11 13 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=7.255 $Y=1.535
+ $X2=7.255 $Y2=3.445
r174 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.255 $Y=1.205
+ $X2=7.255 $Y2=1.37
r175 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.255 $Y=1.205
+ $X2=7.255 $Y2=0.755
r176 2 19 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.605 $X2=5.215 $Y2=3.295
r177 1 24 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.575 $X2=5.215 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%QN 1 2 9 13 17 19 20 21 22 26 27 31 32
c86 32 0 8.77106e-20 $X=8.425 $Y=2.48
c87 27 0 1.98165e-19 $X=9.005 $Y=1.915
c88 21 0 1.02575e-19 $X=8.92 $Y=2.285
c89 19 0 1.18035e-19 $X=8.92 $Y=1.37
r90 31 39 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=3.265
r91 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.48
r92 28 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.42 $Y=2.37
+ $X2=8.42 $Y2=2.48
r93 27 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.915
+ $X2=9.005 $Y2=2.08
r94 27 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.915
+ $X2=9.005 $Y2=1.75
r95 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=1.915 $X2=9.005 $Y2=1.915
r96 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.005 $Y=2.2
+ $X2=9.005 $Y2=1.915
r97 23 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.005 $Y=1.455
+ $X2=9.005 $Y2=1.915
r98 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.505 $Y=2.285
+ $X2=8.42 $Y2=2.37
r99 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=2.285
+ $X2=9.005 $Y2=2.2
r100 21 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=2.285
+ $X2=8.505 $Y2=2.285
r101 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=1.37
+ $X2=9.005 $Y2=1.455
r102 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=1.37
+ $X2=8.505 $Y2=1.37
r103 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=1.285
+ $X2=8.505 $Y2=1.37
r104 15 17 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.42 $Y=1.285
+ $X2=8.42 $Y2=0.74
r105 13 36 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.065 $Y=3.235
+ $X2=9.065 $Y2=2.08
r106 9 35 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=9.065 $Y=0.835
+ $X2=9.065 $Y2=1.75
r107 2 39 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=2.605 $X2=8.42 $Y2=3.265
r108 1 17 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.575 $X2=8.42 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFNR_1%Q 1 2 9 13 16 19 22 25
r20 25 27 6.68493 $w=2.19e-07 $l=1.2e-07 $layer=LI1_cond $X=9.275 $Y=2.807
+ $X2=9.395 $Y2=2.807
r21 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=2.85
+ $X2=9.275 $Y2=2.85
r22 17 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=1.035
+ $X2=9.395 $Y2=1.035
r23 16 27 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.395 $Y=2.68
+ $X2=9.395 $Y2=2.807
r24 15 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.12
+ $X2=9.395 $Y2=1.035
r25 15 16 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=9.395 $Y=1.12
+ $X2=9.395 $Y2=2.68
r26 11 25 2.22295 $w=1.7e-07 $l=1.30476e-07 $layer=LI1_cond $X=9.28 $Y=2.935
+ $X2=9.275 $Y2=2.807
r27 11 13 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.28 $Y=2.935
+ $X2=9.28 $Y2=3.265
r28 7 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=0.95 $X2=9.28
+ $Y2=1.035
r29 7 9 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.28 $Y=0.95 $X2=9.28
+ $Y2=0.74
r30 2 13 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=2.605 $X2=9.28 $Y2=3.265
r31 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.575 $X2=9.28 $Y2=0.74
.ends

