magic
tech sky130A
magscale 1 2
timestamp 1606864600
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 374 1341
<< nmos >>
rect 80 115 110 263
rect 152 115 182 263
rect 252 115 282 263
<< pmos >>
rect 80 817 110 1217
rect 166 817 196 1217
rect 252 817 282 1217
<< ndiff >>
rect 27 199 80 263
rect 27 131 35 199
rect 69 131 80 199
rect 27 115 80 131
rect 110 115 152 263
rect 182 199 252 263
rect 182 131 193 199
rect 227 131 252 199
rect 182 115 252 131
rect 282 199 335 263
rect 282 131 293 199
rect 327 131 335 199
rect 282 115 335 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 861 35 1201
rect 69 861 80 1201
rect 27 817 80 861
rect 110 1201 166 1217
rect 110 861 121 1201
rect 155 861 166 1201
rect 110 817 166 861
rect 196 1201 252 1217
rect 196 861 207 1201
rect 241 861 252 1201
rect 196 817 252 861
rect 282 1201 335 1217
rect 282 861 293 1201
rect 327 861 335 1201
rect 282 817 335 861
<< ndiffc >>
rect 35 131 69 199
rect 193 131 227 199
rect 293 131 327 199
<< pdiffc >>
rect 35 861 69 1201
rect 121 861 155 1201
rect 207 861 241 1201
rect 293 861 327 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 80 586 110 817
rect 27 570 110 586
rect 27 536 37 570
rect 71 536 110 570
rect 27 520 110 536
rect 80 263 110 520
rect 166 518 196 817
rect 252 592 282 817
rect 252 562 289 592
rect 152 502 217 518
rect 152 468 173 502
rect 207 468 217 502
rect 152 452 217 468
rect 152 263 182 452
rect 259 420 289 562
rect 259 404 313 420
rect 259 384 269 404
rect 252 370 269 384
rect 303 370 313 404
rect 252 354 313 370
rect 252 263 282 354
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
<< polycont >>
rect 37 536 71 570
rect 173 468 207 502
rect 269 370 303 404
<< locali >>
rect 0 1311 374 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 374 1311
rect 35 1201 69 1271
rect 121 1201 155 1217
rect 35 845 69 861
rect 105 861 121 879
rect 105 845 155 861
rect 207 1201 241 1271
rect 207 845 241 861
rect 293 1201 327 1217
rect 37 570 71 649
rect 37 520 71 536
rect 105 404 139 845
rect 173 502 207 575
rect 293 535 327 861
rect 173 452 207 468
rect 35 370 269 404
rect 303 370 319 404
rect 35 199 69 370
rect 35 115 69 131
rect 193 199 227 215
rect 193 61 227 131
rect 293 199 327 279
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 37 649 71 683
rect 173 575 207 609
rect 293 501 327 535
rect 293 279 327 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 374 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 374 1311
rect 0 1271 374 1277
rect 25 683 83 689
rect 25 649 37 683
rect 71 649 105 683
rect 25 643 83 649
rect 161 609 219 615
rect 140 575 173 609
rect 207 575 219 609
rect 161 569 219 575
rect 281 535 339 541
rect 281 501 293 535
rect 327 501 339 535
rect 281 495 339 501
rect 293 319 327 495
rect 281 313 339 319
rect 281 279 293 313
rect 327 279 339 313
rect 281 273 339 279
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 311 444 311 444 1 Y
port 1 n
rlabel metal1 55 666 55 666 1 A
port 2 n
rlabel metal1 191 592 191 592 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
