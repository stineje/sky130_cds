* File: sky130_osu_sc_18T_ls__addf_1.spice
* Created: Thu Oct 29 17:33:13 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ls__addf_1.pex.spice"
.subckt sky130_osu_sc_18T_ls__addf_1  GND VDD A B CI CON S CO
* 
* CO	CO
* S	S
* CON	CON
* CI	CI
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1011 N_GND_M1011_d N_A_M1011_g N_A_27_115#_M1011_s N_GND_M1011_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1000 N_A_27_115#_M1000_d N_B_M1000_g N_GND_M1011_d N_GND_M1011_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1001 N_CON_M1001_d N_CI_M1001_g N_A_27_115#_M1000_d N_GND_M1011_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1021 A_368_115# N_B_M1021_g N_CON_M1001_d N_GND_M1011_b NSHORT L=0.15 W=1
+ AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1025 N_GND_M1025_d N_A_M1025_g A_368_115# N_GND_M1011_b NSHORT L=0.15 W=1
+ AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.8
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1018 N_A_526_115#_M1018_d N_A_M1018_g N_GND_M1025_d N_GND_M1011_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75003.2 A=0.15 P=2.3 MULT=1
MM1020 N_GND_M1020_d N_B_M1020_g N_A_526_115#_M1018_d N_GND_M1011_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1013 N_A_526_115#_M1013_d N_CI_M1013_g N_GND_M1020_d N_GND_M1011_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.1 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1014 N_A_784_115#_M1014_d N_CON_M1014_g N_A_526_115#_M1013_d N_GND_M1011_b
+ NSHORT L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 A_870_115# N_B_M1015_g N_A_784_115#_M1014_d N_GND_M1011_b NSHORT L=0.15
+ W=1 AD=0.13 AS=0.14 PD=1.26 PS=1.28 NRD=8.988 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 A_952_115# N_CI_M1005_g A_870_115# N_GND_M1011_b NSHORT L=0.15 W=1
+ AD=0.13 AS=0.13 PD=1.26 PS=1.26 NRD=8.988 NRS=8.988 M=1 R=6.66667 SA=75004.4
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g A_952_115# N_GND_M1011_b NSHORT L=0.15 W=1
+ AD=0.17 AS=0.13 PD=1.34 PS=1.26 NRD=0 NRS=8.988 M=1 R=6.66667 SA=75004.8
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1016 N_S_M1016_d N_A_784_115#_M1016_g N_GND_M1002_d N_GND_M1011_b NSHORT
+ L=0.15 W=1 AD=0.265 AS=0.17 PD=2.53 PS=1.34 NRD=0 NRS=7.188 M=1 R=6.66667
+ SA=75005.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1019 N_CO_M1019_d N_CON_M1019_g N_GND_M1019_s N_GND_M1011_b NSHORT L=0.15 W=1
+ AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_VDD_M1009_d N_A_M1009_g N_A_27_617#_M1009_s N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75005.3 A=0.45 P=6.3 MULT=1
MM1022 N_A_27_617#_M1022_d N_B_M1022_g N_VDD_M1009_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75004.9 A=0.45 P=6.3 MULT=1
MM1012 N_CON_M1012_d N_CI_M1012_g N_A_27_617#_M1022_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001
+ SB=75004.4 A=0.45 P=6.3 MULT=1
MM1004 A_368_617# N_B_M1004_g N_CON_M1012_d N_VDD_M1009_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75001.5 SB=75004
+ A=0.45 P=6.3 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g A_368_617# N_VDD_M1009_b PHIGHVT L=0.15 W=3
+ AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.8
+ SB=75003.6 A=0.45 P=6.3 MULT=1
MM1010 N_A_526_617#_M1010_d N_A_M1010_g N_VDD_M1003_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.3
+ SB=75003.2 A=0.45 P=6.3 MULT=1
MM1027 N_VDD_M1027_d N_B_M1027_g N_A_526_617#_M1010_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.7
+ SB=75002.8 A=0.45 P=6.3 MULT=1
MM1017 N_A_526_617#_M1017_d N_CI_M1017_g N_VDD_M1027_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.1
+ SB=75002.4 A=0.45 P=6.3 MULT=1
MM1008 N_A_784_115#_M1008_d N_CON_M1008_g N_A_526_617#_M1017_d N_VDD_M1009_b
+ PHIGHVT L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20
+ SA=75003.6 SB=75001.9 A=0.45 P=6.3 MULT=1
MM1023 A_870_617# N_B_M1023_g N_A_784_115#_M1008_d N_VDD_M1009_b PHIGHVT L=0.15
+ W=3 AD=0.39 AS=0.42 PD=3.26 PS=3.28 NRD=4.9053 NRS=0 M=1 R=20 SA=75004
+ SB=75001.5 A=0.45 P=6.3 MULT=1
MM1026 A_952_617# N_CI_M1026_g A_870_617# N_VDD_M1009_b PHIGHVT L=0.15 W=3
+ AD=0.39 AS=0.39 PD=3.26 PS=3.26 NRD=4.9053 NRS=4.9053 M=1 R=20 SA=75004.4
+ SB=75001.1 A=0.45 P=6.3 MULT=1
MM1024 N_VDD_M1024_d N_A_M1024_g A_952_617# N_VDD_M1009_b PHIGHVT L=0.15 W=3
+ AD=0.51 AS=0.39 PD=3.34 PS=3.26 NRD=0 NRS=4.9053 M=1 R=20 SA=75004.8
+ SB=75000.7 A=0.45 P=6.3 MULT=1
MM1006 N_S_M1006_d N_A_784_115#_M1006_g N_VDD_M1024_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.51 PD=6.53 PS=3.34 NRD=0 NRS=3.9203 M=1 R=20
+ SA=75005.3 SB=75000.2 A=0.45 P=6.3 MULT=1
MM1007 N_CO_M1007_d N_CON_M1007_g N_VDD_M1007_s N_VDD_M1009_b PHIGHVT L=0.15 W=3
+ AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX28_noxref N_GND_M1011_b N_VDD_M1009_b NWDIODE A=27.436 P=22.04
pX29_noxref noxref_20 A A PROBETYPE=1
pX30_noxref noxref_21 B B PROBETYPE=1
pX31_noxref noxref_22 CI CI PROBETYPE=1
pX32_noxref noxref_23 S S PROBETYPE=1
pX33_noxref noxref_24 CON CON PROBETYPE=1
pX34_noxref noxref_25 CO CO PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__addf_1.pxi.spice"
*
.ends
*
*
