* File: sky130_osu_sc_15T_ms__addf_1.pex.spice
* Created: Fri Nov 12 14:39:29 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%GND 1 2 3 4 5 81 83 91 93 103 105 112
+ 114 127 129 136 153 155
r182 153 155 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r183 138 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=0.152
+ $X2=6.32 $Y2=0.152
r184 134 149 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.152
r185 134 136 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.74
r186 130 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.152
+ $X2=5.31 $Y2=0.152
r187 129 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.152
+ $X2=6.32 $Y2=0.152
r188 125 148 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.152
r189 125 127 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.74
r190 115 147 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0.152
+ $X2=3.2 $Y2=0.152
r191 114 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=0.152
+ $X2=5.31 $Y2=0.152
r192 110 147 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.152
r193 110 112 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.74
r194 105 147 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.152
+ $X2=3.2 $Y2=0.152
r195 101 103 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.34 $Y=0.305
+ $X2=2.34 $Y2=0.74
r196 94 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r197 89 143 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r198 89 91 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r199 83 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r200 81 155 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r201 81 153 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r202 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.34 $Y2=0.305
r203 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.255 $Y2=0.152
r204 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.425 $Y2=0.152
r205 81 138 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.46 $Y=0.152
+ $X2=6.405 $Y2=0.152
r206 81 129 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.235 $Y2=0.152
r207 81 130 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.395 $Y2=0.152
r208 81 114 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=0.152
+ $X2=5.225 $Y2=0.152
r209 81 115 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.285 $Y2=0.152
r210 81 105 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.115 $Y2=0.152
r211 81 106 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.425 $Y2=0.152
r212 81 93 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.255 $Y2=0.152
r213 81 94 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r214 81 83 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r215 5 136 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.195
+ $Y=0.575 $X2=6.32 $Y2=0.74
r216 4 127 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=5.17
+ $Y=0.575 $X2=5.31 $Y2=0.74
r217 3 112 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.575 $X2=3.2 $Y2=0.74
r218 2 103 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.2
+ $Y=0.575 $X2=2.34 $Y2=0.74
r219 1 91 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%VDD 1 2 3 4 5 61 63 70 74 82 86 92 96
+ 106 110 116 122 131 135
r110 131 135 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=6.46 $Y2=5.397
r111 122 135 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=5.36
+ $X2=6.46 $Y2=5.36
r112 120 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=5.397
+ $X2=6.32 $Y2=5.397
r113 120 122 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.405 $Y=5.397
+ $X2=6.46 $Y2=5.397
r114 116 119 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.32 $Y=3.215
+ $X2=6.32 $Y2=4.575
r115 114 129 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.32 $Y=5.245
+ $X2=6.32 $Y2=5.397
r116 114 119 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.32 $Y=5.245
+ $X2=6.32 $Y2=4.575
r117 111 128 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=5.397
+ $X2=5.31 $Y2=5.397
r118 111 113 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.395 $Y=5.397
+ $X2=5.78 $Y2=5.397
r119 110 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=5.397
+ $X2=6.32 $Y2=5.397
r120 110 113 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=6.235 $Y=5.397
+ $X2=5.78 $Y2=5.397
r121 106 109 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.31 $Y=3.895
+ $X2=5.31 $Y2=4.575
r122 104 128 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.31 $Y=5.245
+ $X2=5.31 $Y2=5.397
r123 104 109 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.31 $Y=5.245
+ $X2=5.31 $Y2=4.575
r124 101 103 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=4.42 $Y=5.397
+ $X2=5.1 $Y2=5.397
r125 99 101 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.74 $Y=5.397
+ $X2=4.42 $Y2=5.397
r126 97 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=5.397
+ $X2=3.2 $Y2=5.397
r127 97 99 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.285 $Y=5.397
+ $X2=3.74 $Y2=5.397
r128 96 128 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=5.397
+ $X2=5.31 $Y2=5.397
r129 96 103 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.225 $Y=5.397
+ $X2=5.1 $Y2=5.397
r130 92 95 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.2 $Y=3.895
+ $X2=3.2 $Y2=4.575
r131 90 127 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.2 $Y=5.245
+ $X2=3.2 $Y2=5.397
r132 90 95 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.2 $Y=5.245
+ $X2=3.2 $Y2=4.575
r133 87 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=5.397
+ $X2=2.34 $Y2=5.397
r134 87 89 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=2.425 $Y=5.397
+ $X2=3.06 $Y2=5.397
r135 86 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=5.397
+ $X2=3.2 $Y2=5.397
r136 86 89 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.115 $Y=5.397
+ $X2=3.06 $Y2=5.397
r137 82 85 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.34 $Y=3.555
+ $X2=2.34 $Y2=4.575
r138 80 126 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.34 $Y=5.245
+ $X2=2.34 $Y2=5.397
r139 80 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.34 $Y=5.245
+ $X2=2.34 $Y2=4.575
r140 77 79 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=5.397
+ $X2=1.7 $Y2=5.397
r141 75 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r142 75 77 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r143 74 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=5.397
+ $X2=2.34 $Y2=5.397
r144 74 79 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=2.255 $Y=5.397
+ $X2=1.7 $Y2=5.397
r145 70 73 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=3.895
+ $X2=0.69 $Y2=4.575
r146 68 124 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r147 68 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.575
r148 65 131 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r149 63 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r150 63 65 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r151 61 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=5.245 $X2=6.46 $Y2=5.33
r152 61 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=5.245 $X2=5.78 $Y2=5.33
r153 61 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=5.245 $X2=5.1 $Y2=5.33
r154 61 101 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=5.245 $X2=4.42 $Y2=5.33
r155 61 99 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r156 61 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r157 61 126 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r158 61 79 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r159 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r160 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r161 5 119 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=6.195
+ $Y=2.825 $X2=6.32 $Y2=4.575
r162 5 116 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=6.195
+ $Y=2.825 $X2=6.32 $Y2=3.215
r163 4 109 400 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=2.825 $X2=5.31 $Y2=4.575
r164 4 106 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=2.825 $X2=5.31 $Y2=3.895
r165 3 95 400 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=2.825 $X2=3.2 $Y2=4.575
r166 3 92 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=2.825 $X2=3.2 $Y2=3.895
r167 2 85 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.2
+ $Y=2.825 $X2=2.34 $Y2=4.575
r168 2 82 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=2.2
+ $Y=2.825 $X2=2.34 $Y2=3.555
r169 1 73 400 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.575
r170 1 70 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%A 3 6 8 10 11 13 14 15 16 17 19 22 23 25
+ 28 31 36 37 39 40 45 48 49 51 52 54 59 64 68 69 70 71 73 80
c208 71 0 6.92007e-20 $X=2.64 $Y=1.59
c209 69 0 1.32295e-19 $X=0.63 $Y=1.59
c210 68 0 1.77566e-19 $X=2.35 $Y=1.59
c211 52 0 2.67871e-19 $X=5.13 $Y=2.665
c212 40 0 3.73323e-20 $X=2.495 $Y=1.425
c213 31 0 1.32911e-19 $X=5.095 $Y=3.825
c214 19 0 1.74961e-19 $X=2.435 $Y=2.55
c215 14 0 9.53445e-20 $X=2.36 $Y=1.5
r216 71 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.64 $Y=1.59
+ $X2=2.495 $Y2=1.59
r217 70 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.01 $Y=1.59
+ $X2=5.155 $Y2=1.59
r218 70 71 2.28203 $w=1.7e-07 $l=2.37e-06 $layer=MET1_cond $X=5.01 $Y=1.59
+ $X2=2.64 $Y2=1.59
r219 69 73 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=1.59
+ $X2=0.485 $Y2=1.59
r220 68 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.35 $Y=1.59
+ $X2=2.495 $Y2=1.59
r221 68 69 1.65616 $w=1.7e-07 $l=1.72e-06 $layer=MET1_cond $X=2.35 $Y=1.59
+ $X2=0.63 $Y2=1.59
r222 64 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.155 $Y=1.59
+ $X2=5.155 $Y2=1.59
r223 59 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.495 $Y=1.59
+ $X2=2.495 $Y2=1.59
r224 54 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=1.59
+ $X2=0.485 $Y2=1.59
r225 51 52 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=5.13 $Y=2.515
+ $X2=5.13 $Y2=2.665
r226 50 51 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.165 $Y=1.755
+ $X2=5.165 $Y2=2.515
r227 48 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.59 $X2=5.155 $Y2=1.59
r228 48 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.59
+ $X2=5.155 $Y2=1.755
r229 48 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.59
+ $X2=5.155 $Y2=1.425
r230 44 45 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.435 $Y=2.625
+ $X2=2.555 $Y2=2.625
r231 42 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.59 $X2=2.495 $Y2=1.59
r232 42 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.59
+ $X2=2.495 $Y2=1.755
r233 39 42 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.495 $Y=1.5
+ $X2=2.495 $Y2=1.59
r234 39 40 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.495 $Y=1.5
+ $X2=2.495 $Y2=1.425
r235 36 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.59 $X2=0.485 $Y2=1.59
r236 36 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.59
+ $X2=0.485 $Y2=1.755
r237 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.59
+ $X2=0.485 $Y2=1.425
r238 31 52 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=5.095 $Y=3.825
+ $X2=5.095 $Y2=2.665
r239 28 49 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.095 $Y=0.945
+ $X2=5.095 $Y2=1.425
r240 23 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.555 $Y=2.7
+ $X2=2.555 $Y2=2.625
r241 23 25 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.555 $Y=2.7
+ $X2=2.555 $Y2=3.825
r242 22 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.555 $Y=0.945
+ $X2=2.555 $Y2=1.425
r243 19 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=2.55
+ $X2=2.435 $Y2=2.625
r244 19 43 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.435 $Y=2.55
+ $X2=2.435 $Y2=1.755
r245 16 44 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=2.625
+ $X2=2.435 $Y2=2.625
r246 16 17 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=2.625
+ $X2=2.2 $Y2=2.625
r247 14 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.36 $Y=1.5
+ $X2=2.495 $Y2=1.5
r248 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=1.5 $X2=2.2
+ $Y2=1.5
r249 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=2.7
+ $X2=2.2 $Y2=2.625
r250 11 13 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.125 $Y=2.7
+ $X2=2.125 $Y2=3.825
r251 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=1.425
+ $X2=2.2 $Y2=1.5
r252 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.125 $Y=1.425
+ $X2=2.125 $Y2=0.945
r253 6 38 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=1.755
r254 3 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=1.425
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%B 3 7 11 15 19 23 27 31 34 40 43 47 52
+ 56 59 65 70 75 79 80 82 84 85 86 87
c228 87 0 6.46001e-20 $X=3.67 $Y=2.332
c229 70 0 1.26882e-19 $X=0.485 $Y=2.33
c230 56 0 9.53445e-20 $X=2.305 $Y=2.33
c231 19 0 1.06533e-19 $X=2.985 $Y=0.945
c232 3 0 3.73323e-20 $X=0.905 $Y=0.945
r233 87 94 0.459737 $w=1.9e-07 $l=6.95999e-07 $layer=MET1_cond $X=3.67 $Y=2.332
+ $X2=2.975 $Y2=2.33
r234 86 96 0.124897 $w=2.19e-07 $l=2.05998e-07 $layer=MET1_cond $X=4.06 $Y=2.332
+ $X2=4.265 $Y2=2.33
r235 86 87 0.386904 $w=1.65e-07 $l=3.9e-07 $layer=MET1_cond $X=4.06 $Y=2.332
+ $X2=3.67 $Y2=2.332
r236 85 92 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.45 $Y=2.33
+ $X2=2.305 $Y2=2.33
r237 84 94 0.0970649 $w=1.9e-07 $l=1.45e-07 $layer=MET1_cond $X=2.83 $Y=2.33
+ $X2=2.975 $Y2=2.33
r238 84 85 0.365895 $w=1.7e-07 $l=3.8e-07 $layer=MET1_cond $X=2.83 $Y=2.33
+ $X2=2.45 $Y2=2.33
r239 80 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=2.33
+ $X2=0.485 $Y2=2.33
r240 80 82 0.0144432 $w=1.7e-07 $l=1.5e-08 $layer=MET1_cond $X=0.63 $Y=2.33
+ $X2=0.645 $Y2=2.33
r241 79 92 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.16 $Y=2.33
+ $X2=2.305 $Y2=2.33
r242 79 82 1.45877 $w=1.7e-07 $l=1.515e-06 $layer=MET1_cond $X=2.16 $Y=2.33
+ $X2=0.645 $Y2=2.33
r243 75 77 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.015 $Y=2.17
+ $X2=2.015 $Y2=2.33
r244 70 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=2.33
+ $X2=0.485 $Y2=2.33
r245 70 72 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.485 $Y=2.33
+ $X2=0.485 $Y2=2.5
r246 65 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.265 $Y=2.33
+ $X2=4.265 $Y2=2.33
r247 62 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=2.33
+ $X2=2.975 $Y2=2.33
r248 59 62 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.975 $Y=1.645
+ $X2=2.975 $Y2=2.33
r249 56 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.305 $Y=2.33
+ $X2=2.305 $Y2=2.33
r250 54 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.33
+ $X2=2.015 $Y2=2.33
r251 54 56 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.1 $Y=2.33
+ $X2=2.305 $Y2=2.33
r252 50 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=2.5
+ $X2=0.485 $Y2=2.5
r253 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.57 $Y=2.5
+ $X2=0.895 $Y2=2.5
r254 47 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=2.33 $X2=4.265 $Y2=2.33
r255 47 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.33
+ $X2=4.265 $Y2=2.495
r256 47 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.33
+ $X2=4.265 $Y2=2.165
r257 43 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.645 $X2=2.975 $Y2=1.645
r258 43 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.645
+ $X2=2.975 $Y2=1.81
r259 43 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.645
+ $X2=2.975 $Y2=1.48
r260 40 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=2.17 $X2=2.015 $Y2=2.17
r261 37 40 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.765 $Y=2.17
+ $X2=2.015 $Y2=2.17
r262 34 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=2.5 $X2=0.895 $Y2=2.5
r263 34 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.5
+ $X2=0.895 $Y2=2.665
r264 34 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.5
+ $X2=0.895 $Y2=2.335
r265 31 49 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=4.275 $Y=3.825
+ $X2=4.275 $Y2=2.495
r266 27 48 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=4.275 $Y=0.945
+ $X2=4.275 $Y2=2.165
r267 23 45 1033.22 $w=1.5e-07 $l=2.015e-06 $layer=POLY_cond $X=2.985 $Y=3.825
+ $X2=2.985 $Y2=1.81
r268 19 44 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.985 $Y=0.945
+ $X2=2.985 $Y2=1.48
r269 13 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.335
+ $X2=1.765 $Y2=2.17
r270 13 15 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=1.765 $Y=2.335
+ $X2=1.765 $Y2=3.825
r271 9 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.005
+ $X2=1.765 $Y2=2.17
r272 9 11 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.765 $Y=2.005
+ $X2=1.765 $Y2=0.945
r273 7 36 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.665
r274 3 35 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=2.335
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%CI 3 7 11 15 19 23 26 30 32 36 42 45 51
+ 55 56 57 58 60 66
c183 56 0 3.15979e-20 $X=1.47 $Y=1.96
c184 11 0 1.8492e-19 $X=3.415 $Y=0.945
c185 7 0 1.26882e-19 $X=1.335 $Y=3.825
c186 3 0 3.73323e-20 $X=1.335 $Y=0.945
r187 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.56 $Y=1.96
+ $X2=3.415 $Y2=1.96
r188 57 66 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.6 $Y=1.96
+ $X2=4.745 $Y2=1.96
r189 57 58 1.0014 $w=1.7e-07 $l=1.04e-06 $layer=MET1_cond $X=4.6 $Y=1.96
+ $X2=3.56 $Y2=1.96
r190 56 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.47 $Y=1.96
+ $X2=1.325 $Y2=1.96
r191 55 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.27 $Y=1.96
+ $X2=3.415 $Y2=1.96
r192 55 56 1.73319 $w=1.7e-07 $l=1.8e-06 $layer=MET1_cond $X=3.27 $Y=1.96
+ $X2=1.47 $Y2=1.96
r193 45 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.745 $Y=1.96
+ $X2=4.745 $Y2=1.96
r194 45 48 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.745 $Y=1.96
+ $X2=4.745 $Y2=2.14
r195 42 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.415 $Y=1.96
+ $X2=3.415 $Y2=1.96
r196 40 51 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=2.245
+ $X2=3.415 $Y2=2.33
r197 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.415 $Y=2.245
+ $X2=3.415 $Y2=1.96
r198 36 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.325 $Y=1.96
+ $X2=1.325 $Y2=1.96
r199 32 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=2.14 $X2=4.745 $Y2=2.14
r200 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=2.14
+ $X2=4.745 $Y2=2.305
r201 32 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=2.14
+ $X2=4.745 $Y2=1.975
r202 30 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=2.33 $X2=3.415 $Y2=2.33
r203 26 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.96 $X2=1.325 $Y2=1.96
r204 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.96
+ $X2=1.325 $Y2=2.125
r205 26 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.96
+ $X2=1.325 $Y2=1.795
r206 23 34 779.404 $w=1.5e-07 $l=1.52e-06 $layer=POLY_cond $X=4.685 $Y=3.825
+ $X2=4.685 $Y2=2.305
r207 19 33 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=4.685 $Y=0.945
+ $X2=4.685 $Y2=1.975
r208 13 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.495
+ $X2=3.415 $Y2=2.33
r209 13 15 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.415 $Y=2.495
+ $X2=3.415 $Y2=3.825
r210 9 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.165
+ $X2=3.415 $Y2=2.33
r211 9 11 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=3.415 $Y=2.165
+ $X2=3.415 $Y2=0.945
r212 7 28 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=1.335 $Y=3.825
+ $X2=1.335 $Y2=2.125
r213 3 27 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.335 $Y=0.945
+ $X2=1.335 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%CON 1 3 9 11 14 18 22 25 27 32 38 43 46
+ 50 54 58 63 68 70 71 72 73 80
c189 73 0 1.47588e-19 $X=4.115 $Y=1.22
c190 63 0 2.18019e-20 $X=3.97 $Y=1.59
c191 54 0 3.15979e-20 $X=1.665 $Y=1.505
c192 43 0 1.74961e-19 $X=1.665 $Y=2.765
c193 32 0 1.77566e-19 $X=1.55 $Y=0.74
c194 27 0 1.71092e-19 $X=6.41 $Y=2.48
c195 25 0 1.3267e-19 $X=3.845 $Y=1.59
c196 9 0 7.46754e-20 $X=3.845 $Y=1.425
r197 73 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.115 $Y=1.22
+ $X2=3.97 $Y2=1.22
r198 72 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.995 $Y=1.22
+ $X2=6.14 $Y2=1.22
r199 72 73 1.81022 $w=1.7e-07 $l=1.88e-06 $layer=MET1_cond $X=5.995 $Y=1.22
+ $X2=4.115 $Y2=1.22
r200 71 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r201 70 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.825 $Y=1.22
+ $X2=3.97 $Y2=1.22
r202 70 71 2.05094 $w=1.7e-07 $l=2.13e-06 $layer=MET1_cond $X=3.825 $Y=1.22
+ $X2=1.695 $Y2=1.22
r203 66 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.14 $Y=1.22
+ $X2=6.14 $Y2=1.22
r204 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.14 $Y=1.22
+ $X2=6.41 $Y2=1.22
r205 61 63 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.59
+ $X2=3.97 $Y2=1.59
r206 56 58 6.89435 $w=1.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=2.857
+ $X2=1.665 $Y2=2.857
r207 52 54 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=1.505
+ $X2=1.665 $Y2=1.505
r208 48 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.305
+ $X2=6.41 $Y2=1.22
r209 48 50 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.41 $Y=1.305
+ $X2=6.41 $Y2=2.48
r210 46 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.97 $Y=1.22
+ $X2=3.97 $Y2=1.22
r211 44 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=1.505
+ $X2=3.97 $Y2=1.59
r212 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.97 $Y=1.505
+ $X2=3.97 $Y2=1.22
r213 43 58 1.22693 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=1.665 $Y=2.765
+ $X2=1.665 $Y2=2.857
r214 42 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.59
+ $X2=1.665 $Y2=1.505
r215 42 43 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.665 $Y=1.59
+ $X2=1.665 $Y2=2.765
r216 38 40 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.55 $Y=3.555
+ $X2=1.55 $Y2=4.575
r217 36 56 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.55 $Y=2.95
+ $X2=1.55 $Y2=2.857
r218 36 38 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.55 $Y=2.95
+ $X2=1.55 $Y2=3.555
r219 35 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r220 32 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.22
r221 30 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.42
+ $X2=1.55 $Y2=1.505
r222 30 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.55 $Y=1.42 $X2=1.55
+ $Y2=1.22
r223 27 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=2.48 $X2=6.41 $Y2=2.48
r224 27 29 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.48
+ $X2=6.442 $Y2=2.645
r225 27 28 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.48
+ $X2=6.442 $Y2=2.315
r226 25 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.59 $X2=3.845 $Y2=1.59
r227 22 29 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=6.535 $Y=3.825
+ $X2=6.535 $Y2=2.645
r228 18 28 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=6.535 $Y=0.945
+ $X2=6.535 $Y2=2.315
r229 12 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.755
+ $X2=3.845 $Y2=1.59
r230 12 14 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=3.845 $Y=1.755
+ $X2=3.845 $Y2=3.825
r231 9 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.425
+ $X2=3.845 $Y2=1.59
r232 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.845 $Y=1.425
+ $X2=3.845 $Y2=0.945
r233 3 40 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.575
r234 3 38 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.555
r235 1 32 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%A_784_115# 1 3 11 15 18 20 21 22 23 25
+ 29 32 34 37 39
c121 37 0 7.55579e-20 $X=4.06 $Y=0.74
c122 34 0 9.63581e-20 $X=5.415 $Y=2.99
c123 20 0 6.46001e-20 $X=3.845 $Y=2.77
c124 18 0 3.07391e-19 $X=5.585 $Y=2.495
c125 15 0 1.71513e-19 $X=5.585 $Y=3.825
c126 11 0 1.71092e-19 $X=5.585 $Y=0.945
r127 39 41 7.30282 $w=2.84e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=2.495
+ $X2=5.585 $Y2=2.495
r128 37 38 10.7394 $w=2.84e-07 $l=2.5e-07 $layer=LI1_cond $X=4.06 $Y=0.737
+ $X2=4.31 $Y2=0.737
r129 33 39 3.73949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=2.66
+ $X2=5.415 $Y2=2.495
r130 33 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.415 $Y=2.66
+ $X2=5.415 $Y2=2.99
r131 31 38 3.73949 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.31 $Y=0.905
+ $X2=4.31 $Y2=0.737
r132 31 32 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.31 $Y=0.905
+ $X2=4.31 $Y2=1.875
r133 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.33 $Y=3.075
+ $X2=5.415 $Y2=2.99
r134 29 30 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=5.33 $Y=3.075
+ $X2=4.145 $Y2=3.075
r135 25 27 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.06 $Y=3.555
+ $X2=4.06 $Y2=4.575
r136 23 30 5.48216 $w=2.66e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=3.16
+ $X2=4.145 $Y2=3.075
r137 23 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.06 $Y=3.16
+ $X2=4.06 $Y2=3.555
r138 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.225 $Y=1.96
+ $X2=4.31 $Y2=1.875
r139 21 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.225 $Y=1.96
+ $X2=3.93 $Y2=1.96
r140 20 30 15.5724 $w=2.66e-07 $l=4.29564e-07 $layer=LI1_cond $X=3.845 $Y=2.77
+ $X2=4.145 $Y2=3.075
r141 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=2.045
+ $X2=3.93 $Y2=1.96
r142 19 20 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.845 $Y=2.045
+ $X2=3.845 $Y2=2.77
r143 18 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.585
+ $Y=2.495 $X2=5.585 $Y2=2.495
r144 13 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.66
+ $X2=5.585 $Y2=2.495
r145 13 15 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=5.585 $Y=2.66
+ $X2=5.585 $Y2=3.825
r146 9 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.33
+ $X2=5.585 $Y2=2.495
r147 9 11 710.181 $w=1.5e-07 $l=1.385e-06 $layer=POLY_cond $X=5.585 $Y=2.33
+ $X2=5.585 $Y2=0.945
r148 3 27 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.92
+ $Y=2.825 $X2=4.06 $Y2=4.575
r149 3 25 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=3.92
+ $Y=2.825 $X2=4.06 $Y2=3.555
r150 1 37 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.575 $X2=4.06 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%A_27_565# 1 2 11 15 19
r13 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=3.555
+ $X2=1.12 $Y2=4.575
r14 17 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.12 $Y=3.285
+ $X2=1.12 $Y2=3.555
r15 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.2
+ $X2=1.12 $Y2=3.285
r16 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.2
+ $X2=0.345 $Y2=3.2
r17 11 13 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=3.555
+ $X2=0.26 $Y2=4.575
r18 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.285
+ $X2=0.345 $Y2=3.2
r19 9 11 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.26 $Y=3.285 $X2=0.26
+ $Y2=3.555
r20 2 21 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r21 2 19 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.555
r22 1 13 300 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r23 1 11 300 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.555
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%A_526_565# 1 2 11 15 19
r12 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.63 $Y=3.555
+ $X2=3.63 $Y2=4.575
r13 17 19 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.63 $Y=3.28
+ $X2=3.63 $Y2=3.555
r14 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=3.195
+ $X2=3.63 $Y2=3.28
r15 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=3.195
+ $X2=2.855 $Y2=3.195
r16 11 13 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.77 $Y=3.555
+ $X2=2.77 $Y2=4.575
r17 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=3.28
+ $X2=2.855 $Y2=3.195
r18 9 11 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.77 $Y=3.28
+ $X2=2.77 $Y2=3.555
r19 2 21 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=2.825 $X2=3.63 $Y2=4.575
r20 2 19 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=2.825 $X2=3.63 $Y2=3.555
r21 1 13 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=2.825 $X2=2.77 $Y2=4.575
r22 1 11 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=2.825 $X2=2.77 $Y2=3.555
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%S 1 3 11 17 22 25 29 32
c49 32 0 1.32911e-19 $X=5.8 $Y=3.075
c50 29 0 1.41304e-19 $X=5.925 $Y=2.99
c51 25 0 1.66087e-19 $X=5.925 $Y=1.96
r52 27 29 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=2.99
+ $X2=5.925 $Y2=2.99
r53 23 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=1.96
+ $X2=5.925 $Y2=1.96
r54 22 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=2.905
+ $X2=5.925 $Y2=2.99
r55 21 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=2.045
+ $X2=5.925 $Y2=1.96
r56 21 22 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.925 $Y=2.045
+ $X2=5.925 $Y2=2.905
r57 17 19 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=5.8 $Y=3.555
+ $X2=5.8 $Y2=4.575
r58 15 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.8 $Y=3.075 $X2=5.8
+ $Y2=3.075
r59 15 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=3.075 $X2=5.8
+ $Y2=2.99
r60 15 17 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.8 $Y=3.075 $X2=5.8
+ $Y2=3.555
r61 9 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=1.875 $X2=5.8
+ $Y2=1.96
r62 9 11 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=5.8 $Y=1.875
+ $X2=5.8 $Y2=0.74
r63 3 19 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=5.66
+ $Y=2.825 $X2=5.8 $Y2=4.575
r64 3 17 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=5.66
+ $Y=2.825 $X2=5.8 $Y2=3.555
r65 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.66
+ $Y=0.575 $X2=5.8 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%CO 1 3 10 20
r15 15 17 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.75 $Y=3.215
+ $X2=6.75 $Y2=4.575
r16 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.75 $Y=2.7 $X2=6.75
+ $Y2=2.7
r17 13 15 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.75 $Y=2.7
+ $X2=6.75 $Y2=3.215
r18 10 13 127.872 $w=1.68e-07 $l=1.96e-06 $layer=LI1_cond $X=6.75 $Y=0.74
+ $X2=6.75 $Y2=2.7
r19 3 17 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=6.61
+ $Y=2.825 $X2=6.75 $Y2=4.575
r20 3 15 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=6.61
+ $Y=2.825 $X2=6.75 $Y2=3.215
r21 1 10 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=6.61
+ $Y=0.575 $X2=6.75 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%A_27_115# 1 2 11 13 14 17
c19 17 0 7.46645e-20 $X=1.12 $Y=0.74
c20 14 0 1.32295e-19 $X=0.345 $Y=1.175
r21 15 17 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.12 $Y=1.09
+ $X2=1.12 $Y2=0.74
r22 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.175
+ $X2=1.12 $Y2=1.09
r23 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.175
+ $X2=0.345 $Y2=1.175
r24 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.09
+ $X2=0.345 $Y2=1.175
r25 9 11 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.26 $Y=1.09 $X2=0.26
+ $Y2=0.74
r26 2 17 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.74
r27 1 11 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__ADDF_1%A_526_115# 1 2 11 13 14 17
c28 17 0 7.46093e-20 $X=3.63 $Y=0.74
c29 13 0 1.16312e-19 $X=3.545 $Y=1.175
c30 11 0 7.46645e-20 $X=2.77 $Y=0.74
r31 15 17 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.63 $Y=1.09
+ $X2=3.63 $Y2=0.74
r32 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=1.175
+ $X2=3.63 $Y2=1.09
r33 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=1.175
+ $X2=2.855 $Y2=1.175
r34 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.09
+ $X2=2.855 $Y2=1.175
r35 9 11 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.77 $Y=1.09 $X2=2.77
+ $Y2=0.74
r36 2 17 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.49
+ $Y=0.575 $X2=3.63 $Y2=0.74
r37 1 11 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.63
+ $Y=0.575 $X2=2.77 $Y2=0.74
.ends

