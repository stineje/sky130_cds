* File: sky130_osu_sc_15T_ls__dffs_l.pxi.spice
* Created: Fri Nov 12 14:56:16 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%GND N_GND_M1001_d N_GND_M1002_s N_GND_M1021_d
+ N_GND_M1009_d N_GND_M1026_d N_GND_M1010_d N_GND_M1013_b N_GND_c_2_p
+ N_GND_c_20_p N_GND_c_21_p N_GND_c_42_p N_GND_c_22_p N_GND_c_61_p N_GND_c_23_p
+ N_GND_c_6_p N_GND_c_7_p N_GND_c_141_p N_GND_c_142_p GND N_GND_c_3_p
+ PM_SKY130_OSU_SC_15T_LS__DFFS_L%GND
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%VDD N_VDD_M1012_s N_VDD_M1022_d N_VDD_M1025_s
+ N_VDD_M1005_d N_VDD_M1017_d N_VDD_M1027_s N_VDD_M1016_d N_VDD_M1029_d
+ N_VDD_M1012_b N_VDD_c_199_p N_VDD_c_200_p N_VDD_c_208_p N_VDD_c_209_p
+ N_VDD_c_217_p N_VDD_c_243_p N_VDD_c_227_p N_VDD_c_231_p N_VDD_c_232_p
+ N_VDD_c_233_p N_VDD_c_203_p N_VDD_c_204_p N_VDD_c_273_p N_VDD_c_274_p
+ N_VDD_c_290_p VDD N_VDD_c_201_p PM_SKY130_OSU_SC_15T_LS__DFFS_L%VDD
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%SN N_SN_M1013_g N_SN_M1012_g N_SN_c_307_n
+ N_SN_M1026_g N_SN_M1016_g N_SN_c_312_n N_SN_c_313_n N_SN_c_315_n N_SN_c_316_n
+ N_SN_c_318_n N_SN_c_326_n SN N_SN_c_327_n PM_SKY130_OSU_SC_15T_LS__DFFS_L%SN
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_152_89# N_A_152_89#_M1023_d
+ N_A_152_89#_M1000_d N_A_152_89#_M1001_g N_A_152_89#_M1022_g
+ N_A_152_89#_c_440_n N_A_152_89#_c_441_n N_A_152_89#_c_442_n
+ N_A_152_89#_c_445_n N_A_152_89#_c_457_n N_A_152_89#_c_460_n
+ N_A_152_89#_c_447_n N_A_152_89#_c_448_n N_A_152_89#_c_461_n
+ N_A_152_89#_c_473_n PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_152_89#
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%D N_D_M1002_g N_D_M1025_g N_D_c_525_n
+ N_D_c_526_n D PM_SKY130_OSU_SC_15T_LS__DFFS_L%D
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%CK N_CK_M1000_g N_CK_M1018_g N_CK_M1011_g
+ N_CK_M1019_g N_CK_M1004_g N_CK_c_561_n N_CK_M1008_g N_CK_c_562_n N_CK_c_563_n
+ N_CK_c_564_n N_CK_c_565_n N_CK_c_568_n N_CK_c_569_n N_CK_c_572_n N_CK_c_573_n
+ N_CK_c_577_n N_CK_c_578_n N_CK_c_579_n N_CK_c_580_n N_CK_c_581_n N_CK_c_582_n
+ N_CK_c_583_n N_CK_c_584_n N_CK_c_585_n N_CK_c_586_n N_CK_c_587_n N_CK_c_588_n
+ N_CK_c_589_n CK PM_SKY130_OSU_SC_15T_LS__DFFS_L%CK
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_27_115# N_A_27_115#_M1013_s
+ N_A_27_115#_M1012_d N_A_27_115#_M1021_g N_A_27_115#_M1005_g
+ N_A_27_115#_c_783_n N_A_27_115#_c_785_n N_A_27_115#_c_786_n
+ N_A_27_115#_c_787_n N_A_27_115#_M1014_g N_A_27_115#_M1024_g
+ N_A_27_115#_c_792_n N_A_27_115#_c_794_n N_A_27_115#_c_795_n
+ N_A_27_115#_c_796_n N_A_27_115#_c_799_n N_A_27_115#_c_801_n
+ N_A_27_115#_c_802_n N_A_27_115#_c_836_n
+ PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_27_115#
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_428_89# N_A_428_89#_M1004_d
+ N_A_428_89#_M1008_d N_A_428_89#_c_908_n N_A_428_89#_M1023_g
+ N_A_428_89#_c_911_n N_A_428_89#_c_912_n N_A_428_89#_c_913_n
+ N_A_428_89#_M1007_g N_A_428_89#_c_915_n N_A_428_89#_M1015_g
+ N_A_428_89#_c_917_n N_A_428_89#_c_918_n N_A_428_89#_M1003_g
+ N_A_428_89#_c_919_n N_A_428_89#_c_920_n N_A_428_89#_c_921_n
+ N_A_428_89#_c_922_n N_A_428_89#_c_923_n N_A_428_89#_c_926_n
+ N_A_428_89#_c_928_n N_A_428_89#_c_932_n N_A_428_89#_c_942_n
+ N_A_428_89#_c_933_n N_A_428_89#_c_934_n N_A_428_89#_c_935_n
+ N_A_428_89#_c_947_n PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_428_89#
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_970_89# N_A_970_89#_M1006_s
+ N_A_970_89#_M1027_d N_A_970_89#_M1009_g N_A_970_89#_M1017_g
+ N_A_970_89#_M1010_g N_A_970_89#_M1029_g N_A_970_89#_c_1105_n
+ N_A_970_89#_c_1106_n N_A_970_89#_c_1107_n N_A_970_89#_c_1108_n
+ N_A_970_89#_c_1109_n N_A_970_89#_c_1110_n N_A_970_89#_c_1111_n
+ N_A_970_89#_c_1112_n N_A_970_89#_c_1114_n N_A_970_89#_c_1115_n
+ N_A_970_89#_c_1116_n N_A_970_89#_c_1117_n N_A_970_89#_c_1120_n
+ N_A_970_89#_c_1121_n N_A_970_89#_c_1122_n N_A_970_89#_c_1123_n
+ PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_970_89#
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_808_115# N_A_808_115#_M1011_d
+ N_A_808_115#_M1015_d N_A_808_115#_M1006_g N_A_808_115#_M1027_g
+ N_A_808_115#_c_1266_n N_A_808_115#_c_1267_n N_A_808_115#_c_1291_n
+ N_A_808_115#_c_1292_n N_A_808_115#_c_1308_n N_A_808_115#_c_1336_n
+ N_A_808_115#_c_1268_n N_A_808_115#_c_1281_n N_A_808_115#_c_1271_n
+ N_A_808_115#_c_1272_n N_A_808_115#_c_1274_n N_A_808_115#_c_1275_n
+ PM_SKY130_OSU_SC_15T_LS__DFFS_L%A_808_115#
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%QN N_QN_M1010_s N_QN_M1029_s N_QN_M1028_g
+ N_QN_M1020_g N_QN_c_1394_n N_QN_c_1395_n N_QN_c_1399_n N_QN_c_1400_n
+ N_QN_c_1402_n N_QN_c_1403_n N_QN_c_1404_n N_QN_c_1405_n QN
+ PM_SKY130_OSU_SC_15T_LS__DFFS_L%QN
x_PM_SKY130_OSU_SC_15T_LS__DFFS_L%Q N_Q_M1028_d N_Q_M1020_d N_Q_c_1479_n
+ N_Q_c_1483_n N_Q_c_1481_n N_Q_c_1482_n N_Q_c_1487_n Q
+ PM_SKY130_OSU_SC_15T_LS__DFFS_L%Q
cc_1 N_GND_M1013_b N_SN_M1013_g 0.0335226f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_SN_M1013_g 0.00450746f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_SN_M1013_g 0.00468827f $X=7.815 $Y=0.19 $X2=0.475 $Y2=0.835
cc_4 N_GND_M1013_b N_SN_M1012_g 0.0715368f $X=-0.05 $Y=0 $X2=0.475 $Y2=4.195
cc_5 N_GND_M1013_b N_SN_c_307_n 0.0173166f $X=-0.05 $Y=0 $X2=6.665 $Y2=1.205
cc_6 N_GND_c_6_p N_SN_c_307_n 0.00591263f $X=6.795 $Y=0.152 $X2=6.665 $Y2=1.205
cc_7 N_GND_c_7_p N_SN_c_307_n 0.00502587f $X=6.88 $Y=0.74 $X2=6.665 $Y2=1.205
cc_8 N_GND_c_3_p N_SN_c_307_n 0.00468827f $X=7.815 $Y=0.19 $X2=6.665 $Y2=1.205
cc_9 N_GND_M1013_b N_SN_M1016_g 0.0764955f $X=-0.05 $Y=0 $X2=6.735 $Y2=4.195
cc_10 N_GND_M1013_b N_SN_c_312_n 0.0474126f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.59
cc_11 N_GND_M1013_b N_SN_c_313_n 0.0416576f $X=-0.05 $Y=0 $X2=6.735 $Y2=1.37
cc_12 N_GND_c_7_p N_SN_c_313_n 0.00161904f $X=6.88 $Y=0.74 $X2=6.735 $Y2=1.37
cc_13 N_GND_M1013_b N_SN_c_315_n 0.012812f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.22
cc_14 N_GND_M1013_b N_SN_c_316_n 0.00299613f $X=-0.05 $Y=0 $X2=6.86 $Y2=1.22
cc_15 N_GND_c_7_p N_SN_c_316_n 0.00785456f $X=6.88 $Y=0.74 $X2=6.86 $Y2=1.22
cc_16 N_GND_M1002_s N_SN_c_318_n 0.00506021f $X=1.515 $Y=0.575 $X2=6.715
+ $Y2=1.22
cc_17 N_GND_M1021_d N_SN_c_318_n 0.0107322f $X=3.25 $Y=0.575 $X2=6.715 $Y2=1.22
cc_18 N_GND_M1009_d N_SN_c_318_n 0.00557645f $X=5 $Y=0.575 $X2=6.715 $Y2=1.22
cc_19 N_GND_M1013_b N_SN_c_318_n 0.0394257f $X=-0.05 $Y=0 $X2=6.715 $Y2=1.22
cc_20 N_GND_c_20_p N_SN_c_318_n 0.00518821f $X=1.05 $Y=0.74 $X2=6.715 $Y2=1.22
cc_21 N_GND_c_21_p N_SN_c_318_n 0.0120854f $X=1.64 $Y=0.865 $X2=6.715 $Y2=1.22
cc_22 N_GND_c_22_p N_SN_c_318_n 0.00602612f $X=3.39 $Y=0.74 $X2=6.715 $Y2=1.22
cc_23 N_GND_c_23_p N_SN_c_318_n 0.0119903f $X=5.14 $Y=0.865 $X2=6.715 $Y2=1.22
cc_24 N_GND_M1013_b N_SN_c_326_n 0.0118483f $X=-0.05 $Y=0 $X2=0.465 $Y2=1.22
cc_25 N_GND_M1013_b N_SN_c_327_n 0.00723018f $X=-0.05 $Y=0 $X2=6.86 $Y2=1.22
cc_26 N_GND_c_7_p N_SN_c_327_n 0.00529633f $X=6.88 $Y=0.74 $X2=6.86 $Y2=1.22
cc_27 N_GND_M1013_b N_A_152_89#_M1001_g 0.0555613f $X=-0.05 $Y=0 $X2=0.835
+ $Y2=0.835
cc_28 N_GND_c_2_p N_A_152_89#_M1001_g 0.00590889f $X=0.965 $Y=0.152 $X2=0.835
+ $Y2=0.835
cc_29 N_GND_c_20_p N_A_152_89#_M1001_g 0.00502587f $X=1.05 $Y=0.74 $X2=0.835
+ $Y2=0.835
cc_30 N_GND_c_21_p N_A_152_89#_M1001_g 0.00573513f $X=1.64 $Y=0.865 $X2=0.835
+ $Y2=0.835
cc_31 N_GND_c_3_p N_A_152_89#_M1001_g 0.00468827f $X=7.815 $Y=0.19 $X2=0.835
+ $Y2=0.835
cc_32 N_GND_M1013_b N_A_152_89#_M1022_g 0.0275072f $X=-0.05 $Y=0 $X2=0.905
+ $Y2=4.195
cc_33 N_GND_M1013_b N_A_152_89#_c_440_n 0.0440769f $X=-0.05 $Y=0 $X2=1.03
+ $Y2=2.045
cc_34 N_GND_M1013_b N_A_152_89#_c_441_n 0.0125993f $X=-0.05 $Y=0 $X2=1.03
+ $Y2=2.045
cc_35 N_GND_M1013_b N_A_152_89#_c_442_n 0.0257731f $X=-0.05 $Y=0 $X2=2.33
+ $Y2=1.505
cc_36 N_GND_c_20_p N_A_152_89#_c_442_n 2.96796e-19 $X=1.05 $Y=0.74 $X2=2.33
+ $Y2=1.505
cc_37 N_GND_c_21_p N_A_152_89#_c_442_n 0.00673409f $X=1.64 $Y=0.865 $X2=2.33
+ $Y2=1.505
cc_38 N_GND_M1013_b N_A_152_89#_c_445_n 0.00367876f $X=-0.05 $Y=0 $X2=1.115
+ $Y2=1.505
cc_39 N_GND_c_20_p N_A_152_89#_c_445_n 0.00263009f $X=1.05 $Y=0.74 $X2=1.115
+ $Y2=1.505
cc_40 N_GND_M1013_b N_A_152_89#_c_447_n 0.00198494f $X=-0.05 $Y=0 $X2=2.415
+ $Y2=1.42
cc_41 N_GND_M1013_b N_A_152_89#_c_448_n 0.00313474f $X=-0.05 $Y=0 $X2=2.515
+ $Y2=0.865
cc_42 N_GND_c_42_p N_A_152_89#_c_448_n 0.0148509f $X=3.305 $Y=0.152 $X2=2.515
+ $Y2=0.865
cc_43 N_GND_c_3_p N_A_152_89#_c_448_n 0.00955491f $X=7.815 $Y=0.19 $X2=2.515
+ $Y2=0.865
cc_44 N_GND_M1013_b N_D_M1002_g 0.0421748f $X=-0.05 $Y=0 $X2=1.855 $Y2=0.945
cc_45 N_GND_c_21_p N_D_M1002_g 0.0086813f $X=1.64 $Y=0.865 $X2=1.855 $Y2=0.945
cc_46 N_GND_c_42_p N_D_M1002_g 0.00606474f $X=3.305 $Y=0.152 $X2=1.855 $Y2=0.945
cc_47 N_GND_c_3_p N_D_M1002_g 0.00468827f $X=7.815 $Y=0.19 $X2=1.855 $Y2=0.945
cc_48 N_GND_M1013_b N_D_M1025_g 0.0367665f $X=-0.05 $Y=0 $X2=1.855 $Y2=3.825
cc_49 N_GND_M1013_b N_D_c_525_n 0.0305253f $X=-0.05 $Y=0 $X2=1.915 $Y2=1.96
cc_50 N_GND_M1013_b N_D_c_526_n 0.00311208f $X=-0.05 $Y=0 $X2=1.915 $Y2=1.96
cc_51 N_GND_M1013_b D 0.01184f $X=-0.05 $Y=0 $X2=1.915 $Y2=1.96
cc_52 N_GND_M1013_b N_CK_c_561_n 0.0311248f $X=-0.05 $Y=0 $X2=5.355 $Y2=2.67
cc_53 N_GND_M1013_b N_CK_c_562_n 0.0444827f $X=-0.05 $Y=0 $X2=5.41 $Y2=2.34
cc_54 N_GND_M1013_b N_CK_c_563_n 0.0244095f $X=-0.05 $Y=0 $X2=2.275 $Y2=2.505
cc_55 N_GND_M1013_b N_CK_c_564_n 0.0254608f $X=-0.05 $Y=0 $X2=2.755 $Y2=1.59
cc_56 N_GND_M1013_b N_CK_c_565_n 0.0173906f $X=-0.05 $Y=0 $X2=2.755 $Y2=1.425
cc_57 N_GND_c_42_p N_CK_c_565_n 0.00606474f $X=3.305 $Y=0.152 $X2=2.755
+ $Y2=1.425
cc_58 N_GND_c_3_p N_CK_c_565_n 0.00468827f $X=7.815 $Y=0.19 $X2=2.755 $Y2=1.425
cc_59 N_GND_M1013_b N_CK_c_568_n 0.0252285f $X=-0.05 $Y=0 $X2=4.025 $Y2=1.59
cc_60 N_GND_M1013_b N_CK_c_569_n 0.0175305f $X=-0.05 $Y=0 $X2=4.025 $Y2=1.425
cc_61 N_GND_c_61_p N_CK_c_569_n 0.00606474f $X=5.055 $Y=0.152 $X2=4.025
+ $Y2=1.425
cc_62 N_GND_c_3_p N_CK_c_569_n 0.00468827f $X=7.815 $Y=0.19 $X2=4.025 $Y2=1.425
cc_63 N_GND_M1013_b N_CK_c_572_n 0.0233827f $X=-0.05 $Y=0 $X2=4.505 $Y2=2.505
cc_64 N_GND_M1013_b N_CK_c_573_n 0.0206446f $X=-0.05 $Y=0 $X2=5.382 $Y2=1.425
cc_65 N_GND_c_23_p N_CK_c_573_n 0.00390533f $X=5.14 $Y=0.865 $X2=5.382 $Y2=1.425
cc_66 N_GND_c_6_p N_CK_c_573_n 0.00606474f $X=6.795 $Y=0.152 $X2=5.382 $Y2=1.425
cc_67 N_GND_c_3_p N_CK_c_573_n 0.00468827f $X=7.815 $Y=0.19 $X2=5.382 $Y2=1.425
cc_68 N_GND_M1013_b N_CK_c_577_n 0.0128304f $X=-0.05 $Y=0 $X2=5.382 $Y2=1.575
cc_69 N_GND_M1013_b N_CK_c_578_n 0.00609317f $X=-0.05 $Y=0 $X2=2.67 $Y2=2.33
cc_70 N_GND_M1013_b N_CK_c_579_n 0.00921066f $X=-0.05 $Y=0 $X2=2.755 $Y2=1.59
cc_71 N_GND_M1013_b N_CK_c_580_n 0.00838835f $X=-0.05 $Y=0 $X2=4.025 $Y2=1.59
cc_72 N_GND_M1013_b N_CK_c_581_n 0.00543853f $X=-0.05 $Y=0 $X2=4.42 $Y2=2.33
cc_73 N_GND_M1013_b N_CK_c_582_n 5.00459e-19 $X=-0.05 $Y=0 $X2=4.11 $Y2=2.33
cc_74 N_GND_M1013_b N_CK_c_583_n 6.58573e-19 $X=-0.05 $Y=0 $X2=5.5 $Y2=2.33
cc_75 N_GND_M1013_b N_CK_c_584_n 0.00276905f $X=-0.05 $Y=0 $X2=2.275 $Y2=2.33
cc_76 N_GND_M1013_b N_CK_c_585_n 0.00265612f $X=-0.05 $Y=0 $X2=4.505 $Y2=2.33
cc_77 N_GND_M1013_b N_CK_c_586_n 0.0345662f $X=-0.05 $Y=0 $X2=4.36 $Y2=2.33
cc_78 N_GND_M1013_b N_CK_c_587_n 0.00714094f $X=-0.05 $Y=0 $X2=2.42 $Y2=2.33
cc_79 N_GND_M1013_b N_CK_c_588_n 0.0181831f $X=-0.05 $Y=0 $X2=5.355 $Y2=2.33
cc_80 N_GND_M1013_b N_CK_c_589_n 0.0041728f $X=-0.05 $Y=0 $X2=4.65 $Y2=2.33
cc_81 N_GND_M1013_b CK 0.00236135f $X=-0.05 $Y=0 $X2=5.5 $Y2=2.33
cc_82 N_GND_M1013_b N_A_27_115#_M1021_g 0.0171814f $X=-0.05 $Y=0 $X2=3.175
+ $Y2=0.945
cc_83 N_GND_c_42_p N_A_27_115#_M1021_g 0.00606474f $X=3.305 $Y=0.152 $X2=3.175
+ $Y2=0.945
cc_84 N_GND_c_22_p N_A_27_115#_M1021_g 0.00308284f $X=3.39 $Y=0.74 $X2=3.175
+ $Y2=0.945
cc_85 N_GND_c_3_p N_A_27_115#_M1021_g 0.00468827f $X=7.815 $Y=0.19 $X2=3.175
+ $Y2=0.945
cc_86 N_GND_M1013_b N_A_27_115#_c_783_n 0.024077f $X=-0.05 $Y=0 $X2=3.53
+ $Y2=1.59
cc_87 N_GND_c_22_p N_A_27_115#_c_783_n 8.60298e-19 $X=3.39 $Y=0.74 $X2=3.53
+ $Y2=1.59
cc_88 N_GND_M1013_b N_A_27_115#_c_785_n 0.0105855f $X=-0.05 $Y=0 $X2=3.25
+ $Y2=1.59
cc_89 N_GND_M1013_b N_A_27_115#_c_786_n 0.0232417f $X=-0.05 $Y=0 $X2=3.53
+ $Y2=2.505
cc_90 N_GND_M1013_b N_A_27_115#_c_787_n 0.0105265f $X=-0.05 $Y=0 $X2=3.25
+ $Y2=2.505
cc_91 N_GND_M1013_b N_A_27_115#_M1014_g 0.0163216f $X=-0.05 $Y=0 $X2=3.605
+ $Y2=0.945
cc_92 N_GND_c_22_p N_A_27_115#_M1014_g 0.00308284f $X=3.39 $Y=0.74 $X2=3.605
+ $Y2=0.945
cc_93 N_GND_c_61_p N_A_27_115#_M1014_g 0.00606474f $X=5.055 $Y=0.152 $X2=3.605
+ $Y2=0.945
cc_94 N_GND_c_3_p N_A_27_115#_M1014_g 0.00468827f $X=7.815 $Y=0.19 $X2=3.605
+ $Y2=0.945
cc_95 N_GND_c_2_p N_A_27_115#_c_792_n 0.00735989f $X=0.965 $Y=0.152 $X2=0.605
+ $Y2=0.88
cc_96 N_GND_c_3_p N_A_27_115#_c_792_n 0.0101399f $X=7.815 $Y=0.19 $X2=0.605
+ $Y2=0.88
cc_97 N_GND_M1013_b N_A_27_115#_c_794_n 0.0151571f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=1.59
cc_98 N_GND_M1013_b N_A_27_115#_c_795_n 0.00871176f $X=-0.05 $Y=0 $X2=3.345
+ $Y2=2.505
cc_99 N_GND_M1013_b N_A_27_115#_c_796_n 0.00154463f $X=-0.05 $Y=0 $X2=0.26
+ $Y2=0.74
cc_100 N_GND_c_2_p N_A_27_115#_c_796_n 0.00706731f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_101 N_GND_c_3_p N_A_27_115#_c_796_n 0.00467951f $X=7.815 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_102 N_GND_M1013_b N_A_27_115#_c_799_n 0.00236783f $X=-0.05 $Y=0 $X2=3.345
+ $Y2=1.59
cc_103 N_GND_c_22_p N_A_27_115#_c_799_n 0.00215957f $X=3.39 $Y=0.74 $X2=3.345
+ $Y2=1.59
cc_104 N_GND_M1013_b N_A_27_115#_c_801_n 0.0341069f $X=-0.05 $Y=0 $X2=3.11
+ $Y2=1.59
cc_105 N_GND_M1013_b N_A_27_115#_c_802_n 0.00235788f $X=-0.05 $Y=0 $X2=0.835
+ $Y2=1.59
cc_106 N_GND_M1013_b N_A_428_89#_c_908_n 0.0173059f $X=-0.05 $Y=0 $X2=2.215
+ $Y2=1.425
cc_107 N_GND_c_42_p N_A_428_89#_c_908_n 0.00606474f $X=3.305 $Y=0.152 $X2=2.215
+ $Y2=1.425
cc_108 N_GND_c_3_p N_A_428_89#_c_908_n 0.00468827f $X=7.815 $Y=0.19 $X2=2.215
+ $Y2=1.425
cc_109 N_GND_M1013_b N_A_428_89#_c_911_n 0.0203057f $X=-0.05 $Y=0 $X2=2.335
+ $Y2=1.965
cc_110 N_GND_M1013_b N_A_428_89#_c_912_n 0.0187566f $X=-0.05 $Y=0 $X2=2.74
+ $Y2=2.04
cc_111 N_GND_M1013_b N_A_428_89#_c_913_n 0.00755029f $X=-0.05 $Y=0 $X2=2.41
+ $Y2=2.04
cc_112 N_GND_M1013_b N_A_428_89#_M1007_g 0.032457f $X=-0.05 $Y=0 $X2=2.815
+ $Y2=3.825
cc_113 N_GND_M1013_b N_A_428_89#_c_915_n 0.0559794f $X=-0.05 $Y=0 $X2=3.89
+ $Y2=2.04
cc_114 N_GND_M1013_b N_A_428_89#_M1015_g 0.0319667f $X=-0.05 $Y=0 $X2=3.965
+ $Y2=3.825
cc_115 N_GND_M1013_b N_A_428_89#_c_917_n 0.0270462f $X=-0.05 $Y=0 $X2=4.37
+ $Y2=2.04
cc_116 N_GND_M1013_b N_A_428_89#_c_918_n 0.0125754f $X=-0.05 $Y=0 $X2=4.445
+ $Y2=1.965
cc_117 N_GND_M1013_b N_A_428_89#_c_919_n 0.0141451f $X=-0.05 $Y=0 $X2=2.335
+ $Y2=1.5
cc_118 N_GND_M1013_b N_A_428_89#_c_920_n 0.00426512f $X=-0.05 $Y=0 $X2=2.815
+ $Y2=2.04
cc_119 N_GND_M1013_b N_A_428_89#_c_921_n 0.00426512f $X=-0.05 $Y=0 $X2=3.965
+ $Y2=2.04
cc_120 N_GND_M1013_b N_A_428_89#_c_922_n 0.0256431f $X=-0.05 $Y=0 $X2=4.505
+ $Y2=1.59
cc_121 N_GND_M1013_b N_A_428_89#_c_923_n 0.01755f $X=-0.05 $Y=0 $X2=4.505
+ $Y2=1.425
cc_122 N_GND_c_61_p N_A_428_89#_c_923_n 0.00606474f $X=5.055 $Y=0.152 $X2=4.505
+ $Y2=1.425
cc_123 N_GND_c_3_p N_A_428_89#_c_923_n 0.00468827f $X=7.815 $Y=0.19 $X2=4.505
+ $Y2=1.425
cc_124 N_GND_M1013_b N_A_428_89#_c_926_n 0.0116005f $X=-0.05 $Y=0 $X2=5.485
+ $Y2=1.59
cc_125 N_GND_c_23_p N_A_428_89#_c_926_n 0.00564434f $X=5.14 $Y=0.865 $X2=5.485
+ $Y2=1.59
cc_126 N_GND_M1013_b N_A_428_89#_c_928_n 0.00549177f $X=-0.05 $Y=0 $X2=5.57
+ $Y2=0.865
cc_127 N_GND_c_23_p N_A_428_89#_c_928_n 4.65312e-19 $X=5.14 $Y=0.865 $X2=5.57
+ $Y2=0.865
cc_128 N_GND_c_6_p N_A_428_89#_c_928_n 0.00747016f $X=6.795 $Y=0.152 $X2=5.57
+ $Y2=0.865
cc_129 N_GND_c_3_p N_A_428_89#_c_928_n 0.00476261f $X=7.815 $Y=0.19 $X2=5.57
+ $Y2=0.865
cc_130 N_GND_M1013_b N_A_428_89#_c_932_n 0.0046852f $X=-0.05 $Y=0 $X2=5.57
+ $Y2=1.905
cc_131 N_GND_M1013_b N_A_428_89#_c_933_n 0.0131399f $X=-0.05 $Y=0 $X2=5.845
+ $Y2=2.84
cc_132 N_GND_M1013_b N_A_428_89#_c_934_n 8.79856e-19 $X=-0.05 $Y=0 $X2=5.57
+ $Y2=1.59
cc_133 N_GND_M1013_b N_A_428_89#_c_935_n 0.0128476f $X=-0.05 $Y=0 $X2=5.845
+ $Y2=1.99
cc_134 N_GND_M1013_b N_A_970_89#_M1009_g 0.0319752f $X=-0.05 $Y=0 $X2=4.925
+ $Y2=0.945
cc_135 N_GND_c_61_p N_A_970_89#_M1009_g 0.00606474f $X=5.055 $Y=0.152 $X2=4.925
+ $Y2=0.945
cc_136 N_GND_c_23_p N_A_970_89#_M1009_g 0.00394143f $X=5.14 $Y=0.865 $X2=4.925
+ $Y2=0.945
cc_137 N_GND_c_3_p N_A_970_89#_M1009_g 0.00468827f $X=7.815 $Y=0.19 $X2=4.925
+ $Y2=0.945
cc_138 N_GND_M1013_b N_A_970_89#_M1017_g 0.0330331f $X=-0.05 $Y=0 $X2=4.925
+ $Y2=3.825
cc_139 N_GND_M1013_b N_A_970_89#_M1010_g 0.0301453f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=0.835
cc_140 N_GND_c_7_p N_A_970_89#_M1010_g 0.00343503f $X=6.88 $Y=0.74 $X2=7.685
+ $Y2=0.835
cc_141 N_GND_c_141_p N_A_970_89#_M1010_g 0.00606474f $X=7.815 $Y=0.152 $X2=7.685
+ $Y2=0.835
cc_142 N_GND_c_142_p N_A_970_89#_M1010_g 0.00308284f $X=7.9 $Y=0.74 $X2=7.685
+ $Y2=0.835
cc_143 N_GND_c_3_p N_A_970_89#_M1010_g 0.00468827f $X=7.815 $Y=0.19 $X2=7.685
+ $Y2=0.835
cc_144 N_GND_M1013_b N_A_970_89#_c_1105_n 0.0263191f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=1.93
cc_145 N_GND_M1013_b N_A_970_89#_c_1106_n 0.0292185f $X=-0.05 $Y=0 $X2=7.57
+ $Y2=1.93
cc_146 N_GND_M1013_b N_A_970_89#_c_1107_n 0.0154776f $X=-0.05 $Y=0 $X2=7.572
+ $Y2=1.765
cc_147 N_GND_M1013_b N_A_970_89#_c_1108_n 0.0139483f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=1.54
cc_148 N_GND_M1013_b N_A_970_89#_c_1109_n 0.0365245f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=2.595
cc_149 N_GND_M1013_b N_A_970_89#_c_1110_n 0.00495925f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=2.745
cc_150 N_GND_M1013_b N_A_970_89#_c_1111_n 0.00396219f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=1.93
cc_151 N_GND_c_6_p N_A_970_89#_c_1112_n 0.00658268f $X=6.795 $Y=0.152 $X2=6.435
+ $Y2=0.91
cc_152 N_GND_c_3_p N_A_970_89#_c_1112_n 0.0099265f $X=7.815 $Y=0.19 $X2=6.435
+ $Y2=0.91
cc_153 N_GND_M1013_b N_A_970_89#_c_1114_n 0.0104445f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=1.845
cc_154 N_GND_M1013_b N_A_970_89#_c_1115_n 0.0140059f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=4.565
cc_155 N_GND_M1013_b N_A_970_89#_c_1116_n 0.0188943f $X=-0.05 $Y=0 $X2=7.57
+ $Y2=1.93
cc_156 N_GND_M1013_b N_A_970_89#_c_1117_n 0.00154674f $X=-0.05 $Y=0 $X2=6.09
+ $Y2=0.74
cc_157 N_GND_c_6_p N_A_970_89#_c_1117_n 0.00732079f $X=6.795 $Y=0.152 $X2=6.09
+ $Y2=0.74
cc_158 N_GND_c_3_p N_A_970_89#_c_1117_n 0.00469007f $X=7.815 $Y=0.19 $X2=6.09
+ $Y2=0.74
cc_159 N_GND_M1013_b N_A_970_89#_c_1120_n 0.00193448f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=1.93
cc_160 N_GND_M1013_b N_A_970_89#_c_1121_n 0.0581356f $X=-0.05 $Y=0 $X2=7.425
+ $Y2=1.93
cc_161 N_GND_M1013_b N_A_970_89#_c_1122_n 0.0017195f $X=-0.05 $Y=0 $X2=5.13
+ $Y2=1.93
cc_162 N_GND_M1013_b N_A_970_89#_c_1123_n 0.00173636f $X=-0.05 $Y=0 $X2=7.57
+ $Y2=1.93
cc_163 N_GND_M1013_b N_A_808_115#_M1006_g 0.0343172f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=0.835
cc_164 N_GND_c_6_p N_A_808_115#_M1006_g 0.00454486f $X=6.795 $Y=0.152 $X2=6.305
+ $Y2=0.835
cc_165 N_GND_c_3_p N_A_808_115#_M1006_g 0.00468827f $X=7.815 $Y=0.19 $X2=6.305
+ $Y2=0.835
cc_166 N_GND_M1013_b N_A_808_115#_M1027_g 0.0548413f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=4.195
cc_167 N_GND_M1013_b N_A_808_115#_c_1266_n 0.0455464f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=1.59
cc_168 N_GND_M1013_b N_A_808_115#_c_1267_n 0.0112983f $X=-0.05 $Y=0 $X2=3.685
+ $Y2=1.59
cc_169 N_GND_M1013_b N_A_808_115#_c_1268_n 0.00313975f $X=-0.05 $Y=0 $X2=4.265
+ $Y2=0.865
cc_170 N_GND_c_61_p N_A_808_115#_c_1268_n 0.014959f $X=5.055 $Y=0.152 $X2=4.265
+ $Y2=0.865
cc_171 N_GND_c_3_p N_A_808_115#_c_1268_n 0.00958198f $X=7.815 $Y=0.19 $X2=4.265
+ $Y2=0.865
cc_172 N_GND_M1013_b N_A_808_115#_c_1271_n 0.00161958f $X=-0.05 $Y=0 $X2=6.1
+ $Y2=1.59
cc_173 N_GND_M1013_b N_A_808_115#_c_1272_n 0.0204013f $X=-0.05 $Y=0 $X2=5.955
+ $Y2=1.59
cc_174 N_GND_c_23_p N_A_808_115#_c_1272_n 5.03331e-19 $X=5.14 $Y=0.865 $X2=5.955
+ $Y2=1.59
cc_175 N_GND_M1013_b N_A_808_115#_c_1274_n 0.00120467f $X=-0.05 $Y=0 $X2=3.83
+ $Y2=1.59
cc_176 N_GND_M1013_b N_A_808_115#_c_1275_n 6.71961e-19 $X=-0.05 $Y=0 $X2=6.1
+ $Y2=1.59
cc_177 N_GND_M1013_b N_QN_M1028_g 0.0685226f $X=-0.05 $Y=0 $X2=8.115 $Y2=0.835
cc_178 N_GND_c_142_p N_QN_M1028_g 0.00308284f $X=7.9 $Y=0.74 $X2=8.115 $Y2=0.835
cc_179 N_GND_c_3_p N_QN_M1028_g 0.00468827f $X=7.815 $Y=0.19 $X2=8.115 $Y2=0.835
cc_180 N_GND_M1013_b N_QN_M1020_g 0.0186095f $X=-0.05 $Y=0 $X2=8.115 $Y2=4.195
cc_181 N_GND_M1013_b N_QN_c_1394_n 0.0291912f $X=-0.05 $Y=0 $X2=8.055 $Y2=2.135
cc_182 N_GND_M1013_b N_QN_c_1395_n 0.0103449f $X=-0.05 $Y=0 $X2=7.47 $Y2=0.74
cc_183 N_GND_c_7_p N_QN_c_1395_n 0.0123103f $X=6.88 $Y=0.74 $X2=7.47 $Y2=0.74
cc_184 N_GND_c_141_p N_QN_c_1395_n 0.00757793f $X=7.815 $Y=0.152 $X2=7.47
+ $Y2=0.74
cc_185 N_GND_c_3_p N_QN_c_1395_n 0.00476261f $X=7.815 $Y=0.19 $X2=7.47 $Y2=0.74
cc_186 N_GND_M1013_b N_QN_c_1399_n 0.00138285f $X=-0.05 $Y=0 $X2=7.47 $Y2=2.7
cc_187 N_GND_M1013_b N_QN_c_1400_n 0.0139574f $X=-0.05 $Y=0 $X2=7.97 $Y2=1.59
cc_188 N_GND_c_142_p N_QN_c_1400_n 0.00556529f $X=7.9 $Y=0.74 $X2=7.97 $Y2=1.59
cc_189 N_GND_M1013_b N_QN_c_1402_n 0.00351986f $X=-0.05 $Y=0 $X2=7.555 $Y2=1.59
cc_190 N_GND_M1013_b N_QN_c_1403_n 0.0176115f $X=-0.05 $Y=0 $X2=7.97 $Y2=2.505
cc_191 N_GND_M1013_b N_QN_c_1404_n 0.00426693f $X=-0.05 $Y=0 $X2=7.555 $Y2=2.505
cc_192 N_GND_M1013_b N_QN_c_1405_n 0.0034889f $X=-0.05 $Y=0 $X2=8.055 $Y2=2.135
cc_193 N_GND_M1013_b QN 0.0029781f $X=-0.05 $Y=0 $X2=7.475 $Y2=2.7
cc_194 N_GND_M1013_b N_Q_c_1479_n 0.0132557f $X=-0.05 $Y=0 $X2=8.33 $Y2=0.74
cc_195 N_GND_c_3_p N_Q_c_1479_n 0.00474182f $X=7.815 $Y=0.19 $X2=8.33 $Y2=0.74
cc_196 N_GND_M1013_b N_Q_c_1481_n 0.0625704f $X=-0.05 $Y=0 $X2=8.445 $Y2=2.9
cc_197 N_GND_M1013_b N_Q_c_1482_n 0.0184431f $X=-0.05 $Y=0 $X2=8.445 $Y2=1.255
cc_198 N_VDD_M1012_b N_SN_M1012_g 0.0868572f $X=-0.05 $Y=2.645 $X2=0.475
+ $Y2=4.195
cc_199 N_VDD_c_199_p N_SN_M1012_g 0.00751602f $X=0.26 $Y=4.565 $X2=0.475
+ $Y2=4.195
cc_200 N_VDD_c_200_p N_SN_M1012_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475
+ $Y2=4.195
cc_201 N_VDD_c_201_p N_SN_M1012_g 0.00429146f $X=7.815 $Y=5.36 $X2=0.475
+ $Y2=4.195
cc_202 N_VDD_M1012_b N_SN_M1016_g 0.070867f $X=-0.05 $Y=2.645 $X2=6.735
+ $Y2=4.195
cc_203 N_VDD_c_203_p N_SN_M1016_g 0.00496961f $X=6.865 $Y=5.397 $X2=6.735
+ $Y2=4.195
cc_204 N_VDD_c_204_p N_SN_M1016_g 0.00751602f $X=6.95 $Y=4.565 $X2=6.735
+ $Y2=4.195
cc_205 N_VDD_c_201_p N_SN_M1016_g 0.00429146f $X=7.815 $Y=5.36 $X2=6.735
+ $Y2=4.195
cc_206 N_VDD_M1012_b N_A_152_89#_M1022_g 0.0752288f $X=-0.05 $Y=2.645 $X2=0.905
+ $Y2=4.195
cc_207 N_VDD_c_200_p N_A_152_89#_M1022_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905
+ $Y2=4.195
cc_208 N_VDD_c_208_p N_A_152_89#_M1022_g 0.00751602f $X=1.12 $Y=4.565 $X2=0.905
+ $Y2=4.195
cc_209 N_VDD_c_209_p N_A_152_89#_M1022_g 0.0242413f $X=1.64 $Y=3.545 $X2=0.905
+ $Y2=4.195
cc_210 N_VDD_c_201_p N_A_152_89#_M1022_g 0.00429146f $X=7.815 $Y=5.36 $X2=0.905
+ $Y2=4.195
cc_211 N_VDD_M1012_b N_A_152_89#_c_441_n 0.00286294f $X=-0.05 $Y=2.645 $X2=1.03
+ $Y2=2.045
cc_212 N_VDD_M1025_s N_A_152_89#_c_457_n 0.0125004f $X=1.515 $Y=2.825 $X2=2.345
+ $Y2=2.925
cc_213 N_VDD_M1012_b N_A_152_89#_c_457_n 0.0286398f $X=-0.05 $Y=2.645 $X2=2.345
+ $Y2=2.925
cc_214 N_VDD_c_209_p N_A_152_89#_c_457_n 0.00952036f $X=1.64 $Y=3.545 $X2=2.345
+ $Y2=2.925
cc_215 N_VDD_M1012_b N_A_152_89#_c_460_n 0.00545748f $X=-0.05 $Y=2.645 $X2=1.115
+ $Y2=2.925
cc_216 N_VDD_M1012_b N_A_152_89#_c_461_n 0.00402069f $X=-0.05 $Y=2.645 $X2=2.515
+ $Y2=3.205
cc_217 N_VDD_c_217_p N_A_152_89#_c_461_n 0.00925832f $X=3.305 $Y=5.397 $X2=2.515
+ $Y2=3.205
cc_218 N_VDD_c_201_p N_A_152_89#_c_461_n 0.00876183f $X=7.815 $Y=5.36 $X2=2.515
+ $Y2=3.205
cc_219 N_VDD_M1012_b N_D_M1025_g 0.022678f $X=-0.05 $Y=2.645 $X2=1.855 $Y2=3.825
cc_220 N_VDD_c_209_p N_D_M1025_g 0.00751602f $X=1.64 $Y=3.545 $X2=1.855
+ $Y2=3.825
cc_221 N_VDD_c_217_p N_D_M1025_g 0.00496961f $X=3.305 $Y=5.397 $X2=1.855
+ $Y2=3.825
cc_222 N_VDD_c_201_p N_D_M1025_g 0.00429146f $X=7.815 $Y=5.36 $X2=1.855
+ $Y2=3.825
cc_223 N_VDD_M1012_b N_CK_M1000_g 0.0205191f $X=-0.05 $Y=2.645 $X2=2.215
+ $Y2=3.825
cc_224 N_VDD_c_217_p N_CK_M1000_g 0.00496961f $X=3.305 $Y=5.397 $X2=2.215
+ $Y2=3.825
cc_225 N_VDD_c_201_p N_CK_M1000_g 0.00429146f $X=7.815 $Y=5.36 $X2=2.215
+ $Y2=3.825
cc_226 N_VDD_M1012_b N_CK_M1019_g 0.0205191f $X=-0.05 $Y=2.645 $X2=4.565
+ $Y2=3.825
cc_227 N_VDD_c_227_p N_CK_M1019_g 0.00496961f $X=5.055 $Y=5.397 $X2=4.565
+ $Y2=3.825
cc_228 N_VDD_c_201_p N_CK_M1019_g 0.00429146f $X=7.815 $Y=5.36 $X2=4.565
+ $Y2=3.825
cc_229 N_VDD_M1012_b N_CK_c_561_n 0.00774555f $X=-0.05 $Y=2.645 $X2=5.355
+ $Y2=2.67
cc_230 N_VDD_M1012_b N_CK_M1008_g 0.0218559f $X=-0.05 $Y=2.645 $X2=5.355
+ $Y2=3.825
cc_231 N_VDD_c_231_p N_CK_M1008_g 0.00362996f $X=5.14 $Y=3.205 $X2=5.355
+ $Y2=3.825
cc_232 N_VDD_c_232_p N_CK_M1008_g 0.00496961f $X=6.005 $Y=5.397 $X2=5.355
+ $Y2=3.825
cc_233 N_VDD_c_233_p N_CK_M1008_g 0.0039843f $X=6.09 $Y=4.565 $X2=5.355
+ $Y2=3.825
cc_234 N_VDD_c_201_p N_CK_M1008_g 0.00429146f $X=7.815 $Y=5.36 $X2=5.355
+ $Y2=3.825
cc_235 N_VDD_M1012_b N_CK_c_563_n 0.00487135f $X=-0.05 $Y=2.645 $X2=2.275
+ $Y2=2.505
cc_236 N_VDD_M1012_b N_CK_c_572_n 0.00487051f $X=-0.05 $Y=2.645 $X2=4.505
+ $Y2=2.505
cc_237 N_VDD_M1012_b N_CK_c_583_n 0.00302835f $X=-0.05 $Y=2.645 $X2=5.5 $Y2=2.33
cc_238 N_VDD_M1012_b N_CK_c_584_n 6.42499e-19 $X=-0.05 $Y=2.645 $X2=2.275
+ $Y2=2.33
cc_239 N_VDD_M1012_b N_CK_c_585_n 0.0022456f $X=-0.05 $Y=2.645 $X2=4.505
+ $Y2=2.33
cc_240 N_VDD_c_231_p N_CK_c_588_n 0.00634153f $X=5.14 $Y=3.205 $X2=5.355
+ $Y2=2.33
cc_241 N_VDD_M1012_b N_A_27_115#_M1005_g 0.019613f $X=-0.05 $Y=2.645 $X2=3.175
+ $Y2=3.825
cc_242 N_VDD_c_217_p N_A_27_115#_M1005_g 0.00496961f $X=3.305 $Y=5.397 $X2=3.175
+ $Y2=3.825
cc_243 N_VDD_c_243_p N_A_27_115#_M1005_g 0.00362996f $X=3.39 $Y=3.545 $X2=3.175
+ $Y2=3.825
cc_244 N_VDD_c_201_p N_A_27_115#_M1005_g 0.00429146f $X=7.815 $Y=5.36 $X2=3.175
+ $Y2=3.825
cc_245 N_VDD_c_243_p N_A_27_115#_c_786_n 8.24975e-19 $X=3.39 $Y=3.545 $X2=3.53
+ $Y2=2.505
cc_246 N_VDD_M1012_b N_A_27_115#_M1024_g 0.0185009f $X=-0.05 $Y=2.645 $X2=3.605
+ $Y2=3.825
cc_247 N_VDD_c_243_p N_A_27_115#_M1024_g 0.00362996f $X=3.39 $Y=3.545 $X2=3.605
+ $Y2=3.825
cc_248 N_VDD_c_227_p N_A_27_115#_M1024_g 0.00496961f $X=5.055 $Y=5.397 $X2=3.605
+ $Y2=3.825
cc_249 N_VDD_c_201_p N_A_27_115#_M1024_g 0.00429146f $X=7.815 $Y=5.36 $X2=3.605
+ $Y2=3.825
cc_250 N_VDD_M1012_b N_A_27_115#_c_794_n 0.0230106f $X=-0.05 $Y=2.645 $X2=0.69
+ $Y2=1.59
cc_251 N_VDD_c_200_p N_A_27_115#_c_794_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69
+ $Y2=1.59
cc_252 N_VDD_c_201_p N_A_27_115#_c_794_n 0.00434939f $X=7.815 $Y=5.36 $X2=0.69
+ $Y2=1.59
cc_253 N_VDD_M1012_b N_A_27_115#_c_795_n 0.00424346f $X=-0.05 $Y=2.645 $X2=3.345
+ $Y2=2.505
cc_254 N_VDD_c_243_p N_A_27_115#_c_795_n 0.004428f $X=3.39 $Y=3.545 $X2=3.345
+ $Y2=2.505
cc_255 N_VDD_M1012_b N_A_428_89#_M1007_g 0.0219042f $X=-0.05 $Y=2.645 $X2=2.815
+ $Y2=3.825
cc_256 N_VDD_c_217_p N_A_428_89#_M1007_g 0.00496961f $X=3.305 $Y=5.397 $X2=2.815
+ $Y2=3.825
cc_257 N_VDD_c_201_p N_A_428_89#_M1007_g 0.00429146f $X=7.815 $Y=5.36 $X2=2.815
+ $Y2=3.825
cc_258 N_VDD_M1012_b N_A_428_89#_M1015_g 0.0218732f $X=-0.05 $Y=2.645 $X2=3.965
+ $Y2=3.825
cc_259 N_VDD_c_227_p N_A_428_89#_M1015_g 0.00496961f $X=5.055 $Y=5.397 $X2=3.965
+ $Y2=3.825
cc_260 N_VDD_c_201_p N_A_428_89#_M1015_g 0.00429146f $X=7.815 $Y=5.36 $X2=3.965
+ $Y2=3.825
cc_261 N_VDD_M1012_b N_A_428_89#_c_942_n 0.00199838f $X=-0.05 $Y=2.645 $X2=5.57
+ $Y2=3.205
cc_262 N_VDD_c_232_p N_A_428_89#_c_942_n 0.00464846f $X=6.005 $Y=5.397 $X2=5.57
+ $Y2=3.205
cc_263 N_VDD_c_233_p N_A_428_89#_c_942_n 0.0222136f $X=6.09 $Y=4.565 $X2=5.57
+ $Y2=3.205
cc_264 N_VDD_c_201_p N_A_428_89#_c_942_n 0.00435496f $X=7.815 $Y=5.36 $X2=5.57
+ $Y2=3.205
cc_265 N_VDD_M1012_b N_A_428_89#_c_933_n 0.00560125f $X=-0.05 $Y=2.645 $X2=5.845
+ $Y2=2.84
cc_266 N_VDD_M1012_b N_A_428_89#_c_947_n 0.0139078f $X=-0.05 $Y=2.645 $X2=5.845
+ $Y2=2.925
cc_267 N_VDD_M1012_b N_A_970_89#_M1017_g 0.0201557f $X=-0.05 $Y=2.645 $X2=4.925
+ $Y2=3.825
cc_268 N_VDD_c_227_p N_A_970_89#_M1017_g 0.00496961f $X=5.055 $Y=5.397 $X2=4.925
+ $Y2=3.825
cc_269 N_VDD_c_231_p N_A_970_89#_M1017_g 0.00362996f $X=5.14 $Y=3.205 $X2=4.925
+ $Y2=3.825
cc_270 N_VDD_c_201_p N_A_970_89#_M1017_g 0.00429146f $X=7.815 $Y=5.36 $X2=4.925
+ $Y2=3.825
cc_271 N_VDD_M1012_b N_A_970_89#_M1029_g 0.0596222f $X=-0.05 $Y=2.645 $X2=7.685
+ $Y2=4.195
cc_272 N_VDD_c_204_p N_A_970_89#_M1029_g 0.0039843f $X=6.95 $Y=4.565 $X2=7.685
+ $Y2=4.195
cc_273 N_VDD_c_273_p N_A_970_89#_M1029_g 0.00496961f $X=7.815 $Y=5.397 $X2=7.685
+ $Y2=4.195
cc_274 N_VDD_c_274_p N_A_970_89#_M1029_g 0.00362996f $X=7.9 $Y=4.225 $X2=7.685
+ $Y2=4.195
cc_275 N_VDD_c_201_p N_A_970_89#_M1029_g 0.00429146f $X=7.815 $Y=5.36 $X2=7.685
+ $Y2=4.195
cc_276 N_VDD_M1012_b N_A_970_89#_c_1110_n 0.00913729f $X=-0.05 $Y=2.645 $X2=7.66
+ $Y2=2.745
cc_277 N_VDD_M1012_b N_A_970_89#_c_1115_n 0.023545f $X=-0.05 $Y=2.645 $X2=6.52
+ $Y2=4.565
cc_278 N_VDD_c_203_p N_A_970_89#_c_1115_n 0.0045126f $X=6.865 $Y=5.397 $X2=6.52
+ $Y2=4.565
cc_279 N_VDD_c_201_p N_A_970_89#_c_1115_n 0.00434939f $X=7.815 $Y=5.36 $X2=6.52
+ $Y2=4.565
cc_280 N_VDD_M1012_b N_A_808_115#_M1027_g 0.0689232f $X=-0.05 $Y=2.645 $X2=6.305
+ $Y2=4.195
cc_281 N_VDD_c_233_p N_A_808_115#_M1027_g 0.00751602f $X=6.09 $Y=4.565 $X2=6.305
+ $Y2=4.195
cc_282 N_VDD_c_203_p N_A_808_115#_M1027_g 0.00496961f $X=6.865 $Y=5.397
+ $X2=6.305 $Y2=4.195
cc_283 N_VDD_c_201_p N_A_808_115#_M1027_g 0.00429146f $X=7.815 $Y=5.36 $X2=6.305
+ $Y2=4.195
cc_284 N_VDD_M1012_b N_A_808_115#_c_1267_n 0.00168314f $X=-0.05 $Y=2.645
+ $X2=3.685 $Y2=1.59
cc_285 N_VDD_M1012_b N_A_808_115#_c_1281_n 0.00402069f $X=-0.05 $Y=2.645
+ $X2=4.265 $Y2=3.545
cc_286 N_VDD_c_227_p N_A_808_115#_c_1281_n 0.0092728f $X=5.055 $Y=5.397
+ $X2=4.265 $Y2=3.545
cc_287 N_VDD_c_201_p N_A_808_115#_c_1281_n 0.00876183f $X=7.815 $Y=5.36
+ $X2=4.265 $Y2=3.545
cc_288 N_VDD_M1012_b N_QN_M1020_g 0.0698409f $X=-0.05 $Y=2.645 $X2=8.115
+ $Y2=4.195
cc_289 N_VDD_c_274_p N_QN_M1020_g 0.00362996f $X=7.9 $Y=4.225 $X2=8.115
+ $Y2=4.195
cc_290 N_VDD_c_290_p N_QN_M1020_g 0.00496961f $X=7.815 $Y=5.36 $X2=8.115
+ $Y2=4.195
cc_291 N_VDD_c_201_p N_QN_M1020_g 0.00429146f $X=7.815 $Y=5.36 $X2=8.115
+ $Y2=4.195
cc_292 N_VDD_M1012_b N_QN_c_1399_n 0.0275535f $X=-0.05 $Y=2.645 $X2=7.47 $Y2=2.7
cc_293 N_VDD_c_204_p N_QN_c_1399_n 0.0222136f $X=6.95 $Y=4.565 $X2=7.47 $Y2=2.7
cc_294 N_VDD_c_273_p N_QN_c_1399_n 0.00477009f $X=7.815 $Y=5.397 $X2=7.47
+ $Y2=2.7
cc_295 N_VDD_c_201_p N_QN_c_1399_n 0.00435496f $X=7.815 $Y=5.36 $X2=7.47 $Y2=2.7
cc_296 N_VDD_M1012_b QN 0.0110667f $X=-0.05 $Y=2.645 $X2=7.475 $Y2=2.7
cc_297 N_VDD_M1012_b N_Q_c_1483_n 0.0217788f $X=-0.05 $Y=2.645 $X2=8.33
+ $Y2=4.225
cc_298 N_VDD_c_290_p N_Q_c_1483_n 0.00477009f $X=7.815 $Y=5.36 $X2=8.33
+ $Y2=4.225
cc_299 N_VDD_c_201_p N_Q_c_1483_n 0.00435496f $X=7.815 $Y=5.36 $X2=8.33
+ $Y2=4.225
cc_300 N_VDD_M1012_b N_Q_c_1481_n 0.0127419f $X=-0.05 $Y=2.645 $X2=8.445 $Y2=2.9
cc_301 N_VDD_M1012_b N_Q_c_1487_n 0.0207082f $X=-0.05 $Y=2.645 $X2=8.33
+ $Y2=3.027
cc_302 N_VDD_M1012_b Q 0.0106945f $X=-0.05 $Y=2.645 $X2=8.325 $Y2=3.07
cc_303 N_SN_c_318_n N_A_152_89#_M1023_d 0.00558831f $X=6.715 $Y=1.22 $X2=2.29
+ $Y2=0.575
cc_304 N_SN_M1013_g N_A_152_89#_M1001_g 0.0541587f $X=0.475 $Y=0.835 $X2=0.835
+ $Y2=0.835
cc_305 N_SN_c_315_n N_A_152_89#_M1001_g 5.71653e-19 $X=0.32 $Y=1.22 $X2=0.835
+ $Y2=0.835
cc_306 N_SN_c_318_n N_A_152_89#_M1001_g 0.0100323f $X=6.715 $Y=1.22 $X2=0.835
+ $Y2=0.835
cc_307 N_SN_M1012_g N_A_152_89#_M1022_g 0.0832006f $X=0.475 $Y=4.195 $X2=0.905
+ $Y2=4.195
cc_308 N_SN_c_312_n N_A_152_89#_c_440_n 0.0541587f $X=0.32 $Y=1.59 $X2=1.03
+ $Y2=2.045
cc_309 N_SN_c_318_n N_A_152_89#_c_442_n 0.0293129f $X=6.715 $Y=1.22 $X2=2.33
+ $Y2=1.505
cc_310 N_SN_c_318_n N_A_152_89#_c_445_n 0.00298029f $X=6.715 $Y=1.22 $X2=1.115
+ $Y2=1.505
cc_311 N_SN_c_318_n N_A_152_89#_c_447_n 0.0151351f $X=6.715 $Y=1.22 $X2=2.415
+ $Y2=1.42
cc_312 N_SN_c_318_n N_A_152_89#_c_473_n 0.0253593f $X=6.715 $Y=1.22 $X2=2.507
+ $Y2=1.155
cc_313 N_SN_c_318_n N_D_M1002_g 0.0116357f $X=6.715 $Y=1.22 $X2=1.855 $Y2=0.945
cc_314 N_SN_c_318_n N_CK_c_564_n 8.06574e-19 $X=6.715 $Y=1.22 $X2=2.755 $Y2=1.59
cc_315 N_SN_c_318_n N_CK_c_565_n 0.0106495f $X=6.715 $Y=1.22 $X2=2.755 $Y2=1.425
cc_316 N_SN_c_318_n N_CK_c_568_n 8.06574e-19 $X=6.715 $Y=1.22 $X2=4.025 $Y2=1.59
cc_317 N_SN_c_318_n N_CK_c_569_n 0.00177838f $X=6.715 $Y=1.22 $X2=4.025
+ $Y2=1.425
cc_318 N_SN_c_318_n N_CK_c_573_n 0.01159f $X=6.715 $Y=1.22 $X2=5.382 $Y2=1.425
cc_319 N_SN_c_318_n N_CK_c_577_n 0.00107886f $X=6.715 $Y=1.22 $X2=5.382
+ $Y2=1.575
cc_320 N_SN_c_318_n N_CK_c_579_n 0.00496158f $X=6.715 $Y=1.22 $X2=2.755 $Y2=1.59
cc_321 N_SN_c_318_n N_CK_c_580_n 0.00118606f $X=6.715 $Y=1.22 $X2=4.025 $Y2=1.59
cc_322 N_SN_c_318_n N_A_27_115#_M1021_g 0.0104272f $X=6.715 $Y=1.22 $X2=3.175
+ $Y2=0.945
cc_323 N_SN_c_318_n N_A_27_115#_c_783_n 2.42482e-19 $X=6.715 $Y=1.22 $X2=3.53
+ $Y2=1.59
cc_324 N_SN_c_318_n N_A_27_115#_M1014_g 0.00491871f $X=6.715 $Y=1.22 $X2=3.605
+ $Y2=0.945
cc_325 N_SN_M1013_g N_A_27_115#_c_792_n 0.00956945f $X=0.475 $Y=0.835 $X2=0.605
+ $Y2=0.88
cc_326 N_SN_c_315_n N_A_27_115#_c_792_n 0.00227392f $X=0.32 $Y=1.22 $X2=0.605
+ $Y2=0.88
cc_327 N_SN_c_318_n N_A_27_115#_c_792_n 0.00579965f $X=6.715 $Y=1.22 $X2=0.605
+ $Y2=0.88
cc_328 N_SN_c_326_n N_A_27_115#_c_792_n 0.00419291f $X=0.465 $Y=1.22 $X2=0.605
+ $Y2=0.88
cc_329 N_SN_M1013_g N_A_27_115#_c_794_n 0.051502f $X=0.475 $Y=0.835 $X2=0.69
+ $Y2=1.59
cc_330 N_SN_c_315_n N_A_27_115#_c_794_n 0.0352919f $X=0.32 $Y=1.22 $X2=0.69
+ $Y2=1.59
cc_331 N_SN_c_318_n N_A_27_115#_c_794_n 0.0201876f $X=6.715 $Y=1.22 $X2=0.69
+ $Y2=1.59
cc_332 N_SN_c_326_n N_A_27_115#_c_794_n 0.00217814f $X=0.465 $Y=1.22 $X2=0.69
+ $Y2=1.59
cc_333 N_SN_c_312_n N_A_27_115#_c_796_n 0.00198052f $X=0.32 $Y=1.59 $X2=0.26
+ $Y2=0.74
cc_334 N_SN_c_315_n N_A_27_115#_c_796_n 0.00758432f $X=0.32 $Y=1.22 $X2=0.26
+ $Y2=0.74
cc_335 N_SN_c_326_n N_A_27_115#_c_796_n 0.00633086f $X=0.465 $Y=1.22 $X2=0.26
+ $Y2=0.74
cc_336 N_SN_c_318_n N_A_27_115#_c_799_n 0.00527975f $X=6.715 $Y=1.22 $X2=3.345
+ $Y2=1.59
cc_337 N_SN_c_318_n N_A_27_115#_c_801_n 0.183238f $X=6.715 $Y=1.22 $X2=3.11
+ $Y2=1.59
cc_338 N_SN_c_312_n N_A_27_115#_c_802_n 0.00336326f $X=0.32 $Y=1.59 $X2=0.835
+ $Y2=1.59
cc_339 N_SN_c_315_n N_A_27_115#_c_802_n 0.00667526f $X=0.32 $Y=1.22 $X2=0.835
+ $Y2=1.59
cc_340 N_SN_c_318_n N_A_27_115#_c_802_n 0.0252695f $X=6.715 $Y=1.22 $X2=0.835
+ $Y2=1.59
cc_341 N_SN_c_318_n N_A_27_115#_c_836_n 0.0259207f $X=6.715 $Y=1.22 $X2=3.255
+ $Y2=1.59
cc_342 N_SN_c_318_n N_A_428_89#_M1004_d 0.0042281f $X=6.715 $Y=1.22 $X2=5.43
+ $Y2=0.575
cc_343 N_SN_c_318_n N_A_428_89#_c_908_n 0.0102209f $X=6.715 $Y=1.22 $X2=2.215
+ $Y2=1.425
cc_344 N_SN_c_318_n N_A_428_89#_c_922_n 0.00232964f $X=6.715 $Y=1.22 $X2=4.505
+ $Y2=1.59
cc_345 N_SN_c_318_n N_A_428_89#_c_923_n 0.0103799f $X=6.715 $Y=1.22 $X2=4.505
+ $Y2=1.425
cc_346 N_SN_c_318_n N_A_428_89#_c_926_n 0.0115848f $X=6.715 $Y=1.22 $X2=5.485
+ $Y2=1.59
cc_347 N_SN_c_318_n N_A_428_89#_c_928_n 0.0255624f $X=6.715 $Y=1.22 $X2=5.57
+ $Y2=0.865
cc_348 N_SN_c_318_n N_A_428_89#_c_935_n 4.57217e-19 $X=6.715 $Y=1.22 $X2=5.845
+ $Y2=1.99
cc_349 N_SN_c_318_n N_A_970_89#_M1009_g 0.0100216f $X=6.715 $Y=1.22 $X2=4.925
+ $Y2=0.945
cc_350 N_SN_c_313_n N_A_970_89#_M1010_g 0.00257345f $X=6.735 $Y=1.37 $X2=7.685
+ $Y2=0.835
cc_351 N_SN_M1016_g N_A_970_89#_c_1106_n 0.00575596f $X=6.735 $Y=4.195 $X2=7.57
+ $Y2=1.93
cc_352 N_SN_c_313_n N_A_970_89#_c_1108_n 0.00211346f $X=6.735 $Y=1.37 $X2=7.66
+ $Y2=1.54
cc_353 N_SN_c_307_n N_A_970_89#_c_1112_n 0.00658297f $X=6.665 $Y=1.205 $X2=6.435
+ $Y2=0.91
cc_354 N_SN_c_318_n N_A_970_89#_c_1112_n 0.00992087f $X=6.715 $Y=1.22 $X2=6.435
+ $Y2=0.91
cc_355 N_SN_c_307_n N_A_970_89#_c_1114_n 0.00637042f $X=6.665 $Y=1.205 $X2=6.52
+ $Y2=1.845
cc_356 N_SN_c_313_n N_A_970_89#_c_1114_n 0.0123936f $X=6.735 $Y=1.37 $X2=6.52
+ $Y2=1.845
cc_357 N_SN_c_316_n N_A_970_89#_c_1114_n 0.026885f $X=6.86 $Y=1.22 $X2=6.52
+ $Y2=1.845
cc_358 N_SN_c_318_n N_A_970_89#_c_1114_n 0.0233408f $X=6.715 $Y=1.22 $X2=6.52
+ $Y2=1.845
cc_359 N_SN_c_327_n N_A_970_89#_c_1114_n 0.00211162f $X=6.86 $Y=1.22 $X2=6.52
+ $Y2=1.845
cc_360 N_SN_M1016_g N_A_970_89#_c_1115_n 0.0406135f $X=6.735 $Y=4.195 $X2=6.52
+ $Y2=4.565
cc_361 N_SN_M1016_g N_A_970_89#_c_1116_n 0.0140209f $X=6.735 $Y=4.195 $X2=7.57
+ $Y2=1.93
cc_362 N_SN_c_313_n N_A_970_89#_c_1116_n 0.00362913f $X=6.735 $Y=1.37 $X2=7.57
+ $Y2=1.93
cc_363 N_SN_c_316_n N_A_970_89#_c_1116_n 0.00587817f $X=6.86 $Y=1.22 $X2=7.57
+ $Y2=1.93
cc_364 N_SN_c_318_n N_A_970_89#_c_1116_n 9.00052e-19 $X=6.715 $Y=1.22 $X2=7.57
+ $Y2=1.93
cc_365 N_SN_c_327_n N_A_970_89#_c_1116_n 0.00125279f $X=6.86 $Y=1.22 $X2=7.57
+ $Y2=1.93
cc_366 N_SN_c_318_n N_A_970_89#_c_1117_n 0.00562997f $X=6.715 $Y=1.22 $X2=6.09
+ $Y2=0.74
cc_367 N_SN_M1016_g N_A_970_89#_c_1121_n 0.00850956f $X=6.735 $Y=4.195 $X2=7.425
+ $Y2=1.93
cc_368 N_SN_c_313_n N_A_970_89#_c_1121_n 0.00178318f $X=6.735 $Y=1.37 $X2=7.425
+ $Y2=1.93
cc_369 N_SN_c_316_n N_A_970_89#_c_1121_n 0.00162152f $X=6.86 $Y=1.22 $X2=7.425
+ $Y2=1.93
cc_370 N_SN_c_318_n N_A_970_89#_c_1121_n 0.0209725f $X=6.715 $Y=1.22 $X2=7.425
+ $Y2=1.93
cc_371 N_SN_c_327_n N_A_970_89#_c_1121_n 0.0140445f $X=6.86 $Y=1.22 $X2=7.425
+ $Y2=1.93
cc_372 N_SN_M1016_g N_A_970_89#_c_1123_n 7.50694e-19 $X=6.735 $Y=4.195 $X2=7.57
+ $Y2=1.93
cc_373 N_SN_c_318_n N_A_808_115#_M1011_d 0.0051762f $X=6.715 $Y=1.22 $X2=4.04
+ $Y2=0.575
cc_374 N_SN_c_307_n N_A_808_115#_M1006_g 0.0595025f $X=6.665 $Y=1.205 $X2=6.305
+ $Y2=0.835
cc_375 N_SN_c_313_n N_A_808_115#_M1006_g 0.0571754f $X=6.735 $Y=1.37 $X2=6.305
+ $Y2=0.835
cc_376 N_SN_c_318_n N_A_808_115#_M1006_g 0.00789198f $X=6.715 $Y=1.22 $X2=6.305
+ $Y2=0.835
cc_377 N_SN_M1016_g N_A_808_115#_c_1266_n 0.0571754f $X=6.735 $Y=4.195 $X2=6.305
+ $Y2=1.59
cc_378 N_SN_c_318_n N_A_808_115#_c_1266_n 0.00412631f $X=6.715 $Y=1.22 $X2=6.305
+ $Y2=1.59
cc_379 N_SN_c_318_n N_A_808_115#_c_1267_n 0.00616681f $X=6.715 $Y=1.22 $X2=3.685
+ $Y2=1.59
cc_380 N_SN_c_318_n N_A_808_115#_c_1291_n 0.0536303f $X=6.715 $Y=1.22 $X2=4.095
+ $Y2=1.17
cc_381 N_SN_c_318_n N_A_808_115#_c_1292_n 0.0129425f $X=6.715 $Y=1.22 $X2=3.77
+ $Y2=1.17
cc_382 N_SN_c_318_n N_A_808_115#_c_1271_n 0.00261991f $X=6.715 $Y=1.22 $X2=6.1
+ $Y2=1.59
cc_383 N_SN_c_318_n N_A_808_115#_c_1272_n 0.176894f $X=6.715 $Y=1.22 $X2=5.955
+ $Y2=1.59
cc_384 N_SN_c_318_n N_A_808_115#_c_1274_n 0.0252354f $X=6.715 $Y=1.22 $X2=3.83
+ $Y2=1.59
cc_385 N_SN_c_318_n N_A_808_115#_c_1275_n 0.0267298f $X=6.715 $Y=1.22 $X2=6.1
+ $Y2=1.59
cc_386 N_SN_c_307_n N_QN_c_1395_n 0.00524207f $X=6.665 $Y=1.205 $X2=7.47
+ $Y2=0.74
cc_387 N_SN_c_313_n N_QN_c_1395_n 0.00233719f $X=6.735 $Y=1.37 $X2=7.47 $Y2=0.74
cc_388 N_SN_c_316_n N_QN_c_1395_n 0.0104081f $X=6.86 $Y=1.22 $X2=7.47 $Y2=0.74
cc_389 N_SN_c_327_n N_QN_c_1395_n 0.00696569f $X=6.86 $Y=1.22 $X2=7.47 $Y2=0.74
cc_390 N_SN_M1016_g N_QN_c_1399_n 0.0385239f $X=6.735 $Y=4.195 $X2=7.47 $Y2=2.7
cc_391 N_SN_M1016_g N_QN_c_1402_n 0.00376438f $X=6.735 $Y=4.195 $X2=7.555
+ $Y2=1.59
cc_392 N_SN_c_313_n N_QN_c_1402_n 2.90827e-19 $X=6.735 $Y=1.37 $X2=7.555
+ $Y2=1.59
cc_393 N_SN_c_316_n N_QN_c_1402_n 0.00119452f $X=6.86 $Y=1.22 $X2=7.555 $Y2=1.59
cc_394 N_SN_M1016_g N_QN_c_1404_n 0.00454519f $X=6.735 $Y=4.195 $X2=7.555
+ $Y2=2.505
cc_395 N_SN_M1016_g QN 0.00491824f $X=6.735 $Y=4.195 $X2=7.475 $Y2=2.7
cc_396 N_SN_c_318_n A_386_115# 0.00911585f $X=6.715 $Y=1.22 $X2=1.93 $Y2=0.575
cc_397 N_SN_c_318_n A_578_115# 0.0100396f $X=6.715 $Y=1.22 $X2=2.89 $Y2=0.575
cc_398 N_SN_c_318_n A_736_115# 0.00106636f $X=6.715 $Y=1.22 $X2=3.68 $Y2=0.575
cc_399 N_SN_c_318_n A_928_115# 0.00917995f $X=6.715 $Y=1.22 $X2=4.64 $Y2=0.575
cc_400 N_A_152_89#_c_441_n N_D_M1002_g 0.00508967f $X=1.03 $Y=2.045 $X2=1.855
+ $Y2=0.945
cc_401 N_A_152_89#_c_442_n N_D_M1002_g 0.0123125f $X=2.33 $Y=1.505 $X2=1.855
+ $Y2=0.945
cc_402 N_A_152_89#_c_441_n N_D_M1025_g 0.0129373f $X=1.03 $Y=2.045 $X2=1.855
+ $Y2=3.825
cc_403 N_A_152_89#_c_457_n N_D_M1025_g 0.0211938f $X=2.345 $Y=2.925 $X2=1.855
+ $Y2=3.825
cc_404 N_A_152_89#_c_440_n N_D_c_525_n 0.00628944f $X=1.03 $Y=2.045 $X2=1.915
+ $Y2=1.96
cc_405 N_A_152_89#_c_441_n N_D_c_525_n 0.00131071f $X=1.03 $Y=2.045 $X2=1.915
+ $Y2=1.96
cc_406 N_A_152_89#_c_442_n N_D_c_525_n 0.00207628f $X=2.33 $Y=1.505 $X2=1.915
+ $Y2=1.96
cc_407 N_A_152_89#_c_440_n N_D_c_526_n 0.00168445f $X=1.03 $Y=2.045 $X2=1.915
+ $Y2=1.96
cc_408 N_A_152_89#_c_442_n N_D_c_526_n 0.0086486f $X=2.33 $Y=1.505 $X2=1.915
+ $Y2=1.96
cc_409 N_A_152_89#_c_440_n D 0.00279288f $X=1.03 $Y=2.045 $X2=1.915 $Y2=1.96
cc_410 N_A_152_89#_c_442_n D 0.00200799f $X=2.33 $Y=1.505 $X2=1.915 $Y2=1.96
cc_411 N_A_152_89#_c_457_n N_CK_M1000_g 0.0153421f $X=2.345 $Y=2.925 $X2=2.215
+ $Y2=3.825
cc_412 N_A_152_89#_c_457_n N_CK_c_563_n 0.00150627f $X=2.345 $Y=2.925 $X2=2.275
+ $Y2=2.505
cc_413 N_A_152_89#_c_442_n N_CK_c_564_n 9.45214e-19 $X=2.33 $Y=1.505 $X2=2.755
+ $Y2=1.59
cc_414 N_A_152_89#_c_473_n N_CK_c_564_n 0.00168646f $X=2.507 $Y=1.155 $X2=2.755
+ $Y2=1.59
cc_415 N_A_152_89#_c_447_n N_CK_c_565_n 0.00464203f $X=2.415 $Y=1.42 $X2=2.755
+ $Y2=1.425
cc_416 N_A_152_89#_c_473_n N_CK_c_565_n 0.00381867f $X=2.507 $Y=1.155 $X2=2.755
+ $Y2=1.425
cc_417 N_A_152_89#_c_442_n N_CK_c_578_n 0.0019742f $X=2.33 $Y=1.505 $X2=2.67
+ $Y2=2.33
cc_418 N_A_152_89#_c_457_n N_CK_c_578_n 0.00883015f $X=2.345 $Y=2.925 $X2=2.67
+ $Y2=2.33
cc_419 N_A_152_89#_c_442_n N_CK_c_579_n 0.012316f $X=2.33 $Y=1.505 $X2=2.755
+ $Y2=1.59
cc_420 N_A_152_89#_c_473_n N_CK_c_579_n 5.27251e-19 $X=2.507 $Y=1.155 $X2=2.755
+ $Y2=1.59
cc_421 N_A_152_89#_c_442_n N_CK_c_584_n 0.00224444f $X=2.33 $Y=1.505 $X2=2.275
+ $Y2=2.33
cc_422 N_A_152_89#_c_457_n N_CK_c_584_n 0.0101098f $X=2.345 $Y=2.925 $X2=2.275
+ $Y2=2.33
cc_423 N_A_152_89#_c_457_n N_CK_c_586_n 0.00601583f $X=2.345 $Y=2.925 $X2=4.36
+ $Y2=2.33
cc_424 N_A_152_89#_c_457_n N_CK_c_587_n 0.00409373f $X=2.345 $Y=2.925 $X2=2.42
+ $Y2=2.33
cc_425 N_A_152_89#_M1001_g N_A_27_115#_c_792_n 0.00556511f $X=0.835 $Y=0.835
+ $X2=0.605 $Y2=0.88
cc_426 N_A_152_89#_M1001_g N_A_27_115#_c_794_n 0.0237748f $X=0.835 $Y=0.835
+ $X2=0.69 $Y2=1.59
cc_427 N_A_152_89#_M1022_g N_A_27_115#_c_794_n 0.0224702f $X=0.905 $Y=4.195
+ $X2=0.69 $Y2=1.59
cc_428 N_A_152_89#_c_440_n N_A_27_115#_c_794_n 0.00720273f $X=1.03 $Y=2.045
+ $X2=0.69 $Y2=1.59
cc_429 N_A_152_89#_c_441_n N_A_27_115#_c_794_n 0.0874214f $X=1.03 $Y=2.045
+ $X2=0.69 $Y2=1.59
cc_430 N_A_152_89#_c_445_n N_A_27_115#_c_794_n 0.0124515f $X=1.115 $Y=1.505
+ $X2=0.69 $Y2=1.59
cc_431 N_A_152_89#_c_460_n N_A_27_115#_c_794_n 0.013584f $X=1.115 $Y=2.925
+ $X2=0.69 $Y2=1.59
cc_432 N_A_152_89#_M1001_g N_A_27_115#_c_801_n 0.0065801f $X=0.835 $Y=0.835
+ $X2=3.11 $Y2=1.59
cc_433 N_A_152_89#_c_440_n N_A_27_115#_c_801_n 0.00224331f $X=1.03 $Y=2.045
+ $X2=3.11 $Y2=1.59
cc_434 N_A_152_89#_c_441_n N_A_27_115#_c_801_n 0.00977499f $X=1.03 $Y=2.045
+ $X2=3.11 $Y2=1.59
cc_435 N_A_152_89#_c_442_n N_A_27_115#_c_801_n 0.0532017f $X=2.33 $Y=1.505
+ $X2=3.11 $Y2=1.59
cc_436 N_A_152_89#_c_445_n N_A_27_115#_c_801_n 0.00400514f $X=1.115 $Y=1.505
+ $X2=3.11 $Y2=1.59
cc_437 N_A_152_89#_c_473_n N_A_27_115#_c_801_n 8.67164e-19 $X=2.507 $Y=1.155
+ $X2=3.11 $Y2=1.59
cc_438 N_A_152_89#_M1001_g N_A_27_115#_c_802_n 0.00343239f $X=0.835 $Y=0.835
+ $X2=0.835 $Y2=1.59
cc_439 N_A_152_89#_c_441_n N_A_27_115#_c_802_n 8.0088e-19 $X=1.03 $Y=2.045
+ $X2=0.835 $Y2=1.59
cc_440 N_A_152_89#_c_445_n N_A_27_115#_c_802_n 8.3209e-19 $X=1.115 $Y=1.505
+ $X2=0.835 $Y2=1.59
cc_441 N_A_152_89#_c_442_n N_A_428_89#_c_908_n 0.0022787f $X=2.33 $Y=1.505
+ $X2=2.215 $Y2=1.425
cc_442 N_A_152_89#_c_473_n N_A_428_89#_c_908_n 0.0060945f $X=2.507 $Y=1.155
+ $X2=2.215 $Y2=1.425
cc_443 N_A_152_89#_c_442_n N_A_428_89#_c_911_n 0.00324141f $X=2.33 $Y=1.505
+ $X2=2.335 $Y2=1.965
cc_444 N_A_152_89#_c_442_n N_A_428_89#_c_919_n 0.00993431f $X=2.33 $Y=1.505
+ $X2=2.335 $Y2=1.5
cc_445 N_A_152_89#_c_457_n A_386_565# 0.00732587f $X=2.345 $Y=2.925 $X2=1.93
+ $Y2=2.825
cc_446 N_D_M1025_g N_CK_c_563_n 0.157821f $X=1.855 $Y=3.825 $X2=2.275 $Y2=2.505
cc_447 N_D_c_525_n N_CK_c_579_n 2.89615e-19 $X=1.915 $Y=1.96 $X2=2.755 $Y2=1.59
cc_448 N_D_c_526_n N_CK_c_579_n 0.00478177f $X=1.915 $Y=1.96 $X2=2.755 $Y2=1.59
cc_449 D N_CK_c_579_n 0.00551577f $X=1.915 $Y=1.96 $X2=2.755 $Y2=1.59
cc_450 N_D_M1025_g N_CK_c_584_n 0.00494364f $X=1.855 $Y=3.825 $X2=2.275 $Y2=2.33
cc_451 N_D_M1025_g N_CK_c_587_n 0.00515433f $X=1.855 $Y=3.825 $X2=2.42 $Y2=2.33
cc_452 D N_CK_c_587_n 0.00375733f $X=1.915 $Y=1.96 $X2=2.42 $Y2=2.33
cc_453 N_D_M1002_g N_A_27_115#_c_801_n 0.0030176f $X=1.855 $Y=0.945 $X2=3.11
+ $Y2=1.59
cc_454 N_D_c_525_n N_A_27_115#_c_801_n 7.9412e-19 $X=1.915 $Y=1.96 $X2=3.11
+ $Y2=1.59
cc_455 N_D_c_526_n N_A_27_115#_c_801_n 0.00111625f $X=1.915 $Y=1.96 $X2=3.11
+ $Y2=1.59
cc_456 D N_A_27_115#_c_801_n 0.0353362f $X=1.915 $Y=1.96 $X2=3.11 $Y2=1.59
cc_457 N_D_M1002_g N_A_428_89#_c_908_n 0.0695166f $X=1.855 $Y=0.945 $X2=2.215
+ $Y2=1.425
cc_458 N_D_M1002_g N_A_428_89#_c_911_n 0.00932846f $X=1.855 $Y=0.945 $X2=2.335
+ $Y2=1.965
cc_459 N_D_c_525_n N_A_428_89#_c_911_n 0.0210215f $X=1.915 $Y=1.96 $X2=2.335
+ $Y2=1.965
cc_460 N_D_c_526_n N_A_428_89#_c_911_n 0.00164409f $X=1.915 $Y=1.96 $X2=2.335
+ $Y2=1.965
cc_461 D N_A_428_89#_c_911_n 0.00342011f $X=1.915 $Y=1.96 $X2=2.335 $Y2=1.965
cc_462 D N_A_428_89#_c_913_n 4.62757e-19 $X=1.915 $Y=1.96 $X2=2.41 $Y2=2.04
cc_463 N_CK_c_565_n N_A_27_115#_M1021_g 0.0406519f $X=2.755 $Y=1.425 $X2=3.175
+ $Y2=0.945
cc_464 N_CK_c_579_n N_A_27_115#_M1021_g 0.00109079f $X=2.755 $Y=1.59 $X2=3.175
+ $Y2=0.945
cc_465 N_CK_c_568_n N_A_27_115#_c_783_n 0.0396058f $X=4.025 $Y=1.59 $X2=3.53
+ $Y2=1.59
cc_466 N_CK_c_564_n N_A_27_115#_c_785_n 0.0406519f $X=2.755 $Y=1.59 $X2=3.25
+ $Y2=1.59
cc_467 N_CK_c_586_n N_A_27_115#_c_786_n 0.00772879f $X=4.36 $Y=2.33 $X2=3.53
+ $Y2=2.505
cc_468 N_CK_c_586_n N_A_27_115#_c_787_n 0.00679967f $X=4.36 $Y=2.33 $X2=3.25
+ $Y2=2.505
cc_469 N_CK_c_569_n N_A_27_115#_M1014_g 0.0396058f $X=4.025 $Y=1.425 $X2=3.605
+ $Y2=0.945
cc_470 N_CK_c_580_n N_A_27_115#_M1014_g 3.67139e-19 $X=4.025 $Y=1.59 $X2=3.605
+ $Y2=0.945
cc_471 N_CK_c_564_n N_A_27_115#_c_795_n 7.30049e-19 $X=2.755 $Y=1.59 $X2=3.345
+ $Y2=2.505
cc_472 N_CK_c_578_n N_A_27_115#_c_795_n 0.00401809f $X=2.67 $Y=2.33 $X2=3.345
+ $Y2=2.505
cc_473 N_CK_c_579_n N_A_27_115#_c_795_n 0.0203851f $X=2.755 $Y=1.59 $X2=3.345
+ $Y2=2.505
cc_474 N_CK_c_586_n N_A_27_115#_c_795_n 0.0206884f $X=4.36 $Y=2.33 $X2=3.345
+ $Y2=2.505
cc_475 N_CK_c_564_n N_A_27_115#_c_799_n 7.18106e-19 $X=2.755 $Y=1.59 $X2=3.345
+ $Y2=1.59
cc_476 N_CK_c_579_n N_A_27_115#_c_799_n 0.00742068f $X=2.755 $Y=1.59 $X2=3.345
+ $Y2=1.59
cc_477 N_CK_c_586_n N_A_27_115#_c_799_n 0.00102309f $X=4.36 $Y=2.33 $X2=3.345
+ $Y2=1.59
cc_478 N_CK_c_564_n N_A_27_115#_c_801_n 0.00383172f $X=2.755 $Y=1.59 $X2=3.11
+ $Y2=1.59
cc_479 N_CK_c_578_n N_A_27_115#_c_801_n 0.00443421f $X=2.67 $Y=2.33 $X2=3.11
+ $Y2=1.59
cc_480 N_CK_c_579_n N_A_27_115#_c_801_n 0.0149977f $X=2.755 $Y=1.59 $X2=3.11
+ $Y2=1.59
cc_481 N_CK_c_584_n N_A_27_115#_c_801_n 7.12046e-19 $X=2.275 $Y=2.33 $X2=3.11
+ $Y2=1.59
cc_482 N_CK_c_587_n N_A_27_115#_c_801_n 0.0126164f $X=2.42 $Y=2.33 $X2=3.11
+ $Y2=1.59
cc_483 N_CK_c_564_n N_A_27_115#_c_836_n 3.3031e-19 $X=2.755 $Y=1.59 $X2=3.255
+ $Y2=1.59
cc_484 N_CK_c_579_n N_A_27_115#_c_836_n 0.00143592f $X=2.755 $Y=1.59 $X2=3.255
+ $Y2=1.59
cc_485 N_CK_c_586_n N_A_27_115#_c_836_n 0.0129652f $X=4.36 $Y=2.33 $X2=3.255
+ $Y2=1.59
cc_486 N_CK_c_565_n N_A_428_89#_c_908_n 0.020867f $X=2.755 $Y=1.425 $X2=2.215
+ $Y2=1.425
cc_487 N_CK_c_579_n N_A_428_89#_c_911_n 0.00613747f $X=2.755 $Y=1.59 $X2=2.335
+ $Y2=1.965
cc_488 N_CK_c_564_n N_A_428_89#_c_912_n 0.0183603f $X=2.755 $Y=1.59 $X2=2.74
+ $Y2=2.04
cc_489 N_CK_c_579_n N_A_428_89#_c_912_n 0.00630484f $X=2.755 $Y=1.59 $X2=2.74
+ $Y2=2.04
cc_490 N_CK_c_586_n N_A_428_89#_c_912_n 0.00613485f $X=4.36 $Y=2.33 $X2=2.74
+ $Y2=2.04
cc_491 N_CK_c_563_n N_A_428_89#_c_913_n 0.00904036f $X=2.275 $Y=2.505 $X2=2.41
+ $Y2=2.04
cc_492 N_CK_c_578_n N_A_428_89#_c_913_n 0.00878348f $X=2.67 $Y=2.33 $X2=2.41
+ $Y2=2.04
cc_493 N_CK_c_584_n N_A_428_89#_c_913_n 0.00109468f $X=2.275 $Y=2.33 $X2=2.41
+ $Y2=2.04
cc_494 N_CK_c_587_n N_A_428_89#_c_913_n 0.00137501f $X=2.42 $Y=2.33 $X2=2.41
+ $Y2=2.04
cc_495 N_CK_M1000_g N_A_428_89#_M1007_g 0.0441985f $X=2.215 $Y=3.825 $X2=2.815
+ $Y2=3.825
cc_496 N_CK_c_563_n N_A_428_89#_M1007_g 0.0128384f $X=2.275 $Y=2.505 $X2=2.815
+ $Y2=3.825
cc_497 N_CK_c_578_n N_A_428_89#_M1007_g 0.0081071f $X=2.67 $Y=2.33 $X2=2.815
+ $Y2=3.825
cc_498 N_CK_c_579_n N_A_428_89#_M1007_g 0.00478024f $X=2.755 $Y=1.59 $X2=2.815
+ $Y2=3.825
cc_499 N_CK_c_584_n N_A_428_89#_M1007_g 0.00184124f $X=2.275 $Y=2.33 $X2=2.815
+ $Y2=3.825
cc_500 N_CK_c_586_n N_A_428_89#_M1007_g 0.00938974f $X=4.36 $Y=2.33 $X2=2.815
+ $Y2=3.825
cc_501 N_CK_c_587_n N_A_428_89#_M1007_g 4.2e-19 $X=2.42 $Y=2.33 $X2=2.815
+ $Y2=3.825
cc_502 N_CK_c_586_n N_A_428_89#_c_915_n 0.00607908f $X=4.36 $Y=2.33 $X2=3.89
+ $Y2=2.04
cc_503 N_CK_M1019_g N_A_428_89#_M1015_g 0.0441985f $X=4.565 $Y=3.825 $X2=3.965
+ $Y2=3.825
cc_504 N_CK_c_572_n N_A_428_89#_M1015_g 0.0118393f $X=4.505 $Y=2.505 $X2=3.965
+ $Y2=3.825
cc_505 N_CK_c_580_n N_A_428_89#_M1015_g 0.00399495f $X=4.025 $Y=1.59 $X2=3.965
+ $Y2=3.825
cc_506 N_CK_c_582_n N_A_428_89#_M1015_g 0.00654233f $X=4.11 $Y=2.33 $X2=3.965
+ $Y2=3.825
cc_507 N_CK_c_585_n N_A_428_89#_M1015_g 0.00128351f $X=4.505 $Y=2.33 $X2=3.965
+ $Y2=3.825
cc_508 N_CK_c_586_n N_A_428_89#_M1015_g 0.00497421f $X=4.36 $Y=2.33 $X2=3.965
+ $Y2=3.825
cc_509 N_CK_c_589_n N_A_428_89#_M1015_g 4.2e-19 $X=4.65 $Y=2.33 $X2=3.965
+ $Y2=3.825
cc_510 N_CK_c_572_n N_A_428_89#_c_917_n 0.00904036f $X=4.505 $Y=2.505 $X2=4.37
+ $Y2=2.04
cc_511 N_CK_c_580_n N_A_428_89#_c_917_n 0.00909647f $X=4.025 $Y=1.59 $X2=4.37
+ $Y2=2.04
cc_512 N_CK_c_581_n N_A_428_89#_c_917_n 0.00924811f $X=4.42 $Y=2.33 $X2=4.37
+ $Y2=2.04
cc_513 N_CK_c_585_n N_A_428_89#_c_917_n 0.00102633f $X=4.505 $Y=2.33 $X2=4.37
+ $Y2=2.04
cc_514 N_CK_c_586_n N_A_428_89#_c_917_n 0.00613485f $X=4.36 $Y=2.33 $X2=4.37
+ $Y2=2.04
cc_515 N_CK_c_589_n N_A_428_89#_c_917_n 0.00137501f $X=4.65 $Y=2.33 $X2=4.37
+ $Y2=2.04
cc_516 N_CK_c_580_n N_A_428_89#_c_918_n 0.00649764f $X=4.025 $Y=1.59 $X2=4.445
+ $Y2=1.965
cc_517 N_CK_c_564_n N_A_428_89#_c_919_n 0.0216263f $X=2.755 $Y=1.59 $X2=2.335
+ $Y2=1.5
cc_518 N_CK_c_584_n N_A_428_89#_c_919_n 2.45465e-19 $X=2.275 $Y=2.33 $X2=2.335
+ $Y2=1.5
cc_519 N_CK_c_579_n N_A_428_89#_c_920_n 0.00568091f $X=2.755 $Y=1.59 $X2=2.815
+ $Y2=2.04
cc_520 N_CK_c_568_n N_A_428_89#_c_921_n 0.0183603f $X=4.025 $Y=1.59 $X2=3.965
+ $Y2=2.04
cc_521 N_CK_c_580_n N_A_428_89#_c_921_n 0.00436024f $X=4.025 $Y=1.59 $X2=3.965
+ $Y2=2.04
cc_522 N_CK_c_568_n N_A_428_89#_c_922_n 0.0220721f $X=4.025 $Y=1.59 $X2=4.505
+ $Y2=1.59
cc_523 N_CK_c_572_n N_A_428_89#_c_922_n 0.00227671f $X=4.505 $Y=2.505 $X2=4.505
+ $Y2=1.59
cc_524 N_CK_c_580_n N_A_428_89#_c_922_n 0.00131283f $X=4.025 $Y=1.59 $X2=4.505
+ $Y2=1.59
cc_525 N_CK_c_585_n N_A_428_89#_c_922_n 5.27321e-19 $X=4.505 $Y=2.33 $X2=4.505
+ $Y2=1.59
cc_526 N_CK_c_589_n N_A_428_89#_c_922_n 8.78837e-19 $X=4.65 $Y=2.33 $X2=4.505
+ $Y2=1.59
cc_527 N_CK_c_569_n N_A_428_89#_c_923_n 0.022472f $X=4.025 $Y=1.425 $X2=4.505
+ $Y2=1.425
cc_528 N_CK_c_562_n N_A_428_89#_c_926_n 0.00592387f $X=5.41 $Y=2.34 $X2=5.485
+ $Y2=1.59
cc_529 N_CK_c_568_n N_A_428_89#_c_926_n 8.05876e-19 $X=4.025 $Y=1.59 $X2=5.485
+ $Y2=1.59
cc_530 N_CK_c_572_n N_A_428_89#_c_926_n 5.56676e-19 $X=4.505 $Y=2.505 $X2=5.485
+ $Y2=1.59
cc_531 N_CK_c_577_n N_A_428_89#_c_926_n 0.00762848f $X=5.382 $Y=1.575 $X2=5.485
+ $Y2=1.59
cc_532 N_CK_c_580_n N_A_428_89#_c_926_n 0.00853323f $X=4.025 $Y=1.59 $X2=5.485
+ $Y2=1.59
cc_533 N_CK_c_581_n N_A_428_89#_c_926_n 0.00132011f $X=4.42 $Y=2.33 $X2=5.485
+ $Y2=1.59
cc_534 N_CK_c_583_n N_A_428_89#_c_926_n 8.24249e-19 $X=5.5 $Y=2.33 $X2=5.485
+ $Y2=1.59
cc_535 N_CK_c_585_n N_A_428_89#_c_926_n 0.00261697f $X=4.505 $Y=2.33 $X2=5.485
+ $Y2=1.59
cc_536 N_CK_c_586_n N_A_428_89#_c_926_n 3.12599e-19 $X=4.36 $Y=2.33 $X2=5.485
+ $Y2=1.59
cc_537 N_CK_c_588_n N_A_428_89#_c_926_n 0.00341454f $X=5.355 $Y=2.33 $X2=5.485
+ $Y2=1.59
cc_538 N_CK_c_589_n N_A_428_89#_c_926_n 0.00221563f $X=4.65 $Y=2.33 $X2=5.485
+ $Y2=1.59
cc_539 N_CK_c_573_n N_A_428_89#_c_928_n 0.0117675f $X=5.382 $Y=1.425 $X2=5.57
+ $Y2=0.865
cc_540 N_CK_c_577_n N_A_428_89#_c_928_n 0.0022869f $X=5.382 $Y=1.575 $X2=5.57
+ $Y2=0.865
cc_541 N_CK_c_562_n N_A_428_89#_c_932_n 0.00735778f $X=5.41 $Y=2.34 $X2=5.57
+ $Y2=1.905
cc_542 N_CK_c_561_n N_A_428_89#_c_933_n 0.00333903f $X=5.355 $Y=2.67 $X2=5.845
+ $Y2=2.84
cc_543 N_CK_M1008_g N_A_428_89#_c_933_n 0.00495264f $X=5.355 $Y=3.825 $X2=5.845
+ $Y2=2.84
cc_544 N_CK_c_562_n N_A_428_89#_c_933_n 0.00567067f $X=5.41 $Y=2.34 $X2=5.845
+ $Y2=2.84
cc_545 N_CK_c_583_n N_A_428_89#_c_933_n 0.0289277f $X=5.5 $Y=2.33 $X2=5.845
+ $Y2=2.84
cc_546 CK N_A_428_89#_c_933_n 0.00852929f $X=5.5 $Y=2.33 $X2=5.845 $Y2=2.84
cc_547 N_CK_c_562_n N_A_428_89#_c_934_n 0.00114916f $X=5.41 $Y=2.34 $X2=5.57
+ $Y2=1.59
cc_548 N_CK_c_577_n N_A_428_89#_c_934_n 8.09104e-19 $X=5.382 $Y=1.575 $X2=5.57
+ $Y2=1.59
cc_549 N_CK_c_561_n N_A_428_89#_c_935_n 0.00198338f $X=5.355 $Y=2.67 $X2=5.845
+ $Y2=1.99
cc_550 N_CK_c_562_n N_A_428_89#_c_935_n 0.00559872f $X=5.41 $Y=2.34 $X2=5.845
+ $Y2=1.99
cc_551 N_CK_c_583_n N_A_428_89#_c_935_n 0.00661696f $X=5.5 $Y=2.33 $X2=5.845
+ $Y2=1.99
cc_552 CK N_A_428_89#_c_935_n 0.00236431f $X=5.5 $Y=2.33 $X2=5.845 $Y2=1.99
cc_553 N_CK_c_561_n N_A_428_89#_c_947_n 0.00260941f $X=5.355 $Y=2.67 $X2=5.845
+ $Y2=2.925
cc_554 N_CK_c_583_n N_A_428_89#_c_947_n 0.00706443f $X=5.5 $Y=2.33 $X2=5.845
+ $Y2=2.925
cc_555 CK N_A_428_89#_c_947_n 0.00259785f $X=5.5 $Y=2.33 $X2=5.845 $Y2=2.925
cc_556 N_CK_c_562_n N_A_970_89#_M1009_g 0.00697006f $X=5.41 $Y=2.34 $X2=4.925
+ $Y2=0.945
cc_557 N_CK_c_573_n N_A_970_89#_M1009_g 0.0315481f $X=5.382 $Y=1.425 $X2=4.925
+ $Y2=0.945
cc_558 N_CK_c_561_n N_A_970_89#_M1017_g 0.0294691f $X=5.355 $Y=2.67 $X2=4.925
+ $Y2=3.825
cc_559 N_CK_c_562_n N_A_970_89#_M1017_g 0.0175925f $X=5.41 $Y=2.34 $X2=4.925
+ $Y2=3.825
cc_560 N_CK_c_572_n N_A_970_89#_M1017_g 0.156645f $X=4.505 $Y=2.505 $X2=4.925
+ $Y2=3.825
cc_561 N_CK_c_583_n N_A_970_89#_M1017_g 0.0026346f $X=5.5 $Y=2.33 $X2=4.925
+ $Y2=3.825
cc_562 N_CK_c_585_n N_A_970_89#_M1017_g 0.00453616f $X=4.505 $Y=2.33 $X2=4.925
+ $Y2=3.825
cc_563 N_CK_c_588_n N_A_970_89#_M1017_g 0.0114893f $X=5.355 $Y=2.33 $X2=4.925
+ $Y2=3.825
cc_564 N_CK_c_589_n N_A_970_89#_M1017_g 0.00113587f $X=4.65 $Y=2.33 $X2=4.925
+ $Y2=3.825
cc_565 CK N_A_970_89#_M1017_g 3.05655e-19 $X=5.5 $Y=2.33 $X2=4.925 $Y2=3.825
cc_566 N_CK_c_562_n N_A_970_89#_c_1105_n 0.0213116f $X=5.41 $Y=2.34 $X2=4.985
+ $Y2=1.93
cc_567 N_CK_c_588_n N_A_970_89#_c_1105_n 0.00185875f $X=5.355 $Y=2.33 $X2=4.985
+ $Y2=1.93
cc_568 N_CK_c_562_n N_A_970_89#_c_1111_n 9.0669e-19 $X=5.41 $Y=2.34 $X2=4.985
+ $Y2=1.93
cc_569 N_CK_c_588_n N_A_970_89#_c_1111_n 0.00488871f $X=5.355 $Y=2.33 $X2=4.985
+ $Y2=1.93
cc_570 N_CK_c_562_n N_A_970_89#_c_1121_n 0.00431553f $X=5.41 $Y=2.34 $X2=7.425
+ $Y2=1.93
cc_571 N_CK_c_583_n N_A_970_89#_c_1121_n 5.80133e-19 $X=5.5 $Y=2.33 $X2=7.425
+ $Y2=1.93
cc_572 N_CK_c_588_n N_A_970_89#_c_1121_n 0.0179446f $X=5.355 $Y=2.33 $X2=7.425
+ $Y2=1.93
cc_573 CK N_A_970_89#_c_1121_n 0.0240913f $X=5.5 $Y=2.33 $X2=7.425 $Y2=1.93
cc_574 N_CK_c_562_n N_A_970_89#_c_1122_n 8.66236e-19 $X=5.41 $Y=2.34 $X2=5.13
+ $Y2=1.93
cc_575 N_CK_c_588_n N_A_970_89#_c_1122_n 0.0247156f $X=5.355 $Y=2.33 $X2=5.13
+ $Y2=1.93
cc_576 N_CK_c_561_n N_A_808_115#_M1027_g 0.0044653f $X=5.355 $Y=2.67 $X2=6.305
+ $Y2=4.195
cc_577 N_CK_c_577_n N_A_808_115#_c_1266_n 0.00662135f $X=5.382 $Y=1.575
+ $X2=6.305 $Y2=1.59
cc_578 N_CK_c_569_n N_A_808_115#_c_1267_n 0.00554221f $X=4.025 $Y=1.425
+ $X2=3.685 $Y2=1.59
cc_579 N_CK_c_580_n N_A_808_115#_c_1267_n 0.057541f $X=4.025 $Y=1.59 $X2=3.685
+ $Y2=1.59
cc_580 N_CK_c_582_n N_A_808_115#_c_1267_n 0.0116326f $X=4.11 $Y=2.33 $X2=3.685
+ $Y2=1.59
cc_581 N_CK_c_585_n N_A_808_115#_c_1267_n 0.00613815f $X=4.505 $Y=2.33 $X2=3.685
+ $Y2=1.59
cc_582 N_CK_c_586_n N_A_808_115#_c_1267_n 0.020361f $X=4.36 $Y=2.33 $X2=3.685
+ $Y2=1.59
cc_583 N_CK_c_589_n N_A_808_115#_c_1267_n 6.61118e-19 $X=4.65 $Y=2.33 $X2=3.685
+ $Y2=1.59
cc_584 N_CK_c_568_n N_A_808_115#_c_1291_n 0.00227142f $X=4.025 $Y=1.59 $X2=4.095
+ $Y2=1.17
cc_585 N_CK_c_569_n N_A_808_115#_c_1291_n 0.0147334f $X=4.025 $Y=1.425 $X2=4.095
+ $Y2=1.17
cc_586 N_CK_c_580_n N_A_808_115#_c_1291_n 0.0103267f $X=4.025 $Y=1.59 $X2=4.095
+ $Y2=1.17
cc_587 N_CK_c_572_n N_A_808_115#_c_1308_n 0.00150627f $X=4.505 $Y=2.505
+ $X2=4.095 $Y2=2.925
cc_588 N_CK_c_581_n N_A_808_115#_c_1308_n 0.00843004f $X=4.42 $Y=2.33 $X2=4.095
+ $Y2=2.925
cc_589 N_CK_c_582_n N_A_808_115#_c_1308_n 0.00323798f $X=4.11 $Y=2.33 $X2=4.095
+ $Y2=2.925
cc_590 N_CK_c_585_n N_A_808_115#_c_1308_n 0.00103871f $X=4.505 $Y=2.33 $X2=4.095
+ $Y2=2.925
cc_591 N_CK_c_586_n N_A_808_115#_c_1308_n 0.012754f $X=4.36 $Y=2.33 $X2=4.095
+ $Y2=2.925
cc_592 N_CK_c_589_n N_A_808_115#_c_1308_n 0.00146098f $X=4.65 $Y=2.33 $X2=4.095
+ $Y2=2.925
cc_593 N_CK_c_577_n N_A_808_115#_c_1271_n 3.50905e-19 $X=5.382 $Y=1.575 $X2=6.1
+ $Y2=1.59
cc_594 N_CK_c_562_n N_A_808_115#_c_1272_n 0.00128484f $X=5.41 $Y=2.34 $X2=5.955
+ $Y2=1.59
cc_595 N_CK_c_568_n N_A_808_115#_c_1272_n 0.00362401f $X=4.025 $Y=1.59 $X2=5.955
+ $Y2=1.59
cc_596 N_CK_c_577_n N_A_808_115#_c_1272_n 0.00179204f $X=5.382 $Y=1.575
+ $X2=5.955 $Y2=1.59
cc_597 N_CK_c_580_n N_A_808_115#_c_1272_n 0.0127028f $X=4.025 $Y=1.59 $X2=5.955
+ $Y2=1.59
cc_598 N_CK_c_581_n N_A_808_115#_c_1272_n 0.00451177f $X=4.42 $Y=2.33 $X2=5.955
+ $Y2=1.59
cc_599 N_CK_c_585_n N_A_808_115#_c_1272_n 6.39375e-19 $X=4.505 $Y=2.33 $X2=5.955
+ $Y2=1.59
cc_600 N_CK_c_589_n N_A_808_115#_c_1272_n 0.0144351f $X=4.65 $Y=2.33 $X2=5.955
+ $Y2=1.59
cc_601 N_CK_c_568_n N_A_808_115#_c_1274_n 9.79344e-19 $X=4.025 $Y=1.59 $X2=3.83
+ $Y2=1.59
cc_602 N_CK_c_580_n N_A_808_115#_c_1274_n 0.00180575f $X=4.025 $Y=1.59 $X2=3.83
+ $Y2=1.59
cc_603 N_CK_c_586_n N_A_808_115#_c_1274_n 0.0128239f $X=4.36 $Y=2.33 $X2=3.83
+ $Y2=1.59
cc_604 N_A_27_115#_c_801_n N_A_428_89#_c_911_n 0.00253253f $X=3.11 $Y=1.59
+ $X2=2.335 $Y2=1.965
cc_605 N_A_27_115#_c_801_n N_A_428_89#_c_912_n 0.00296105f $X=3.11 $Y=1.59
+ $X2=2.74 $Y2=2.04
cc_606 N_A_27_115#_c_787_n N_A_428_89#_M1007_g 0.157117f $X=3.25 $Y=2.505
+ $X2=2.815 $Y2=3.825
cc_607 N_A_27_115#_c_795_n N_A_428_89#_M1007_g 0.00486364f $X=3.345 $Y=2.505
+ $X2=2.815 $Y2=3.825
cc_608 N_A_27_115#_c_785_n N_A_428_89#_c_915_n 0.0342351f $X=3.25 $Y=1.59
+ $X2=3.89 $Y2=2.04
cc_609 N_A_27_115#_c_787_n N_A_428_89#_c_915_n 0.0307748f $X=3.25 $Y=2.505
+ $X2=3.89 $Y2=2.04
cc_610 N_A_27_115#_c_795_n N_A_428_89#_c_915_n 0.0113171f $X=3.345 $Y=2.505
+ $X2=3.89 $Y2=2.04
cc_611 N_A_27_115#_c_799_n N_A_428_89#_c_915_n 8.69982e-19 $X=3.345 $Y=1.59
+ $X2=3.89 $Y2=2.04
cc_612 N_A_27_115#_c_801_n N_A_428_89#_c_915_n 0.00486036f $X=3.11 $Y=1.59
+ $X2=3.89 $Y2=2.04
cc_613 N_A_27_115#_c_836_n N_A_428_89#_c_915_n 4.12801e-19 $X=3.255 $Y=1.59
+ $X2=3.89 $Y2=2.04
cc_614 N_A_27_115#_c_786_n N_A_428_89#_M1015_g 0.153702f $X=3.53 $Y=2.505
+ $X2=3.965 $Y2=3.825
cc_615 N_A_27_115#_M1021_g N_A_808_115#_c_1267_n 0.001069f $X=3.175 $Y=0.945
+ $X2=3.685 $Y2=1.59
cc_616 N_A_27_115#_M1005_g N_A_808_115#_c_1267_n 9.36754e-19 $X=3.175 $Y=3.825
+ $X2=3.685 $Y2=1.59
cc_617 N_A_27_115#_c_783_n N_A_808_115#_c_1267_n 0.0061959f $X=3.53 $Y=1.59
+ $X2=3.685 $Y2=1.59
cc_618 N_A_27_115#_c_786_n N_A_808_115#_c_1267_n 0.00738718f $X=3.53 $Y=2.505
+ $X2=3.685 $Y2=1.59
cc_619 N_A_27_115#_M1014_g N_A_808_115#_c_1267_n 0.00502021f $X=3.605 $Y=0.945
+ $X2=3.685 $Y2=1.59
cc_620 N_A_27_115#_M1024_g N_A_808_115#_c_1267_n 0.00479454f $X=3.605 $Y=3.825
+ $X2=3.685 $Y2=1.59
cc_621 N_A_27_115#_c_795_n N_A_808_115#_c_1267_n 0.0702347f $X=3.345 $Y=2.505
+ $X2=3.685 $Y2=1.59
cc_622 N_A_27_115#_c_799_n N_A_808_115#_c_1267_n 0.0157315f $X=3.345 $Y=1.59
+ $X2=3.685 $Y2=1.59
cc_623 N_A_27_115#_c_836_n N_A_808_115#_c_1267_n 4.18442e-19 $X=3.255 $Y=1.59
+ $X2=3.685 $Y2=1.59
cc_624 N_A_27_115#_M1021_g N_A_808_115#_c_1292_n 0.00136315f $X=3.175 $Y=0.945
+ $X2=3.77 $Y2=1.17
cc_625 N_A_27_115#_M1014_g N_A_808_115#_c_1292_n 0.00979345f $X=3.605 $Y=0.945
+ $X2=3.77 $Y2=1.17
cc_626 N_A_27_115#_M1005_g N_A_808_115#_c_1336_n 9.13132e-19 $X=3.175 $Y=3.825
+ $X2=3.77 $Y2=2.925
cc_627 N_A_27_115#_M1024_g N_A_808_115#_c_1336_n 0.0096885f $X=3.605 $Y=3.825
+ $X2=3.77 $Y2=2.925
cc_628 N_A_27_115#_c_783_n N_A_808_115#_c_1274_n 0.00229064f $X=3.53 $Y=1.59
+ $X2=3.83 $Y2=1.59
cc_629 N_A_27_115#_c_799_n N_A_808_115#_c_1274_n 0.0012094f $X=3.345 $Y=1.59
+ $X2=3.83 $Y2=1.59
cc_630 N_A_27_115#_c_836_n N_A_808_115#_c_1274_n 0.0241863f $X=3.255 $Y=1.59
+ $X2=3.83 $Y2=1.59
cc_631 N_A_27_115#_c_792_n A_110_115# 0.00170398f $X=0.605 $Y=0.88 $X2=0.55
+ $Y2=0.575
cc_632 N_A_428_89#_c_918_n N_A_970_89#_M1009_g 0.0073696f $X=4.445 $Y=1.965
+ $X2=4.925 $Y2=0.945
cc_633 N_A_428_89#_c_923_n N_A_970_89#_M1009_g 0.0823485f $X=4.505 $Y=1.425
+ $X2=4.925 $Y2=0.945
cc_634 N_A_428_89#_c_926_n N_A_970_89#_M1009_g 0.0107575f $X=5.485 $Y=1.59
+ $X2=4.925 $Y2=0.945
cc_635 N_A_428_89#_c_917_n N_A_970_89#_c_1105_n 0.0073696f $X=4.37 $Y=2.04
+ $X2=4.985 $Y2=1.93
cc_636 N_A_428_89#_c_926_n N_A_970_89#_c_1105_n 0.00290516f $X=5.485 $Y=1.59
+ $X2=4.985 $Y2=1.93
cc_637 N_A_428_89#_c_935_n N_A_970_89#_c_1105_n 4.7338e-19 $X=5.845 $Y=1.99
+ $X2=4.985 $Y2=1.93
cc_638 N_A_428_89#_c_918_n N_A_970_89#_c_1111_n 0.0035305f $X=4.445 $Y=1.965
+ $X2=4.985 $Y2=1.93
cc_639 N_A_428_89#_c_926_n N_A_970_89#_c_1111_n 0.0219931f $X=5.485 $Y=1.59
+ $X2=4.985 $Y2=1.93
cc_640 N_A_428_89#_c_932_n N_A_970_89#_c_1111_n 0.00215086f $X=5.57 $Y=1.905
+ $X2=4.985 $Y2=1.93
cc_641 N_A_428_89#_c_935_n N_A_970_89#_c_1111_n 0.00359729f $X=5.845 $Y=1.99
+ $X2=4.985 $Y2=1.93
cc_642 N_A_428_89#_c_933_n N_A_970_89#_c_1115_n 0.0272317f $X=5.845 $Y=2.84
+ $X2=6.52 $Y2=4.565
cc_643 N_A_428_89#_c_935_n N_A_970_89#_c_1115_n 0.00224409f $X=5.845 $Y=1.99
+ $X2=6.52 $Y2=4.565
cc_644 N_A_428_89#_c_947_n N_A_970_89#_c_1115_n 0.00644034f $X=5.845 $Y=2.925
+ $X2=6.52 $Y2=4.565
cc_645 N_A_428_89#_c_928_n N_A_970_89#_c_1117_n 0.0179417f $X=5.57 $Y=0.865
+ $X2=6.09 $Y2=0.74
cc_646 N_A_428_89#_c_935_n N_A_970_89#_c_1120_n 0.00254232f $X=5.845 $Y=1.99
+ $X2=6.52 $Y2=1.93
cc_647 N_A_428_89#_c_926_n N_A_970_89#_c_1121_n 0.00314603f $X=5.485 $Y=1.59
+ $X2=7.425 $Y2=1.93
cc_648 N_A_428_89#_c_932_n N_A_970_89#_c_1121_n 0.00659876f $X=5.57 $Y=1.905
+ $X2=7.425 $Y2=1.93
cc_649 N_A_428_89#_c_933_n N_A_970_89#_c_1121_n 0.00167455f $X=5.845 $Y=2.84
+ $X2=7.425 $Y2=1.93
cc_650 N_A_428_89#_c_935_n N_A_970_89#_c_1121_n 0.0235843f $X=5.845 $Y=1.99
+ $X2=7.425 $Y2=1.93
cc_651 N_A_428_89#_c_918_n N_A_970_89#_c_1122_n 9.14174e-19 $X=4.445 $Y=1.965
+ $X2=5.13 $Y2=1.93
cc_652 N_A_428_89#_c_926_n N_A_970_89#_c_1122_n 0.0010261f $X=5.485 $Y=1.59
+ $X2=5.13 $Y2=1.93
cc_653 N_A_428_89#_c_932_n N_A_970_89#_c_1122_n 0.00122156f $X=5.57 $Y=1.905
+ $X2=5.13 $Y2=1.93
cc_654 N_A_428_89#_c_935_n N_A_970_89#_c_1122_n 0.00122726f $X=5.845 $Y=1.99
+ $X2=5.13 $Y2=1.93
cc_655 N_A_428_89#_c_928_n N_A_808_115#_M1006_g 0.00809903f $X=5.57 $Y=0.865
+ $X2=6.305 $Y2=0.835
cc_656 N_A_428_89#_c_932_n N_A_808_115#_M1027_g 0.00280704f $X=5.57 $Y=1.905
+ $X2=6.305 $Y2=4.195
cc_657 N_A_428_89#_c_942_n N_A_808_115#_M1027_g 0.0301523f $X=5.57 $Y=3.205
+ $X2=6.305 $Y2=4.195
cc_658 N_A_428_89#_c_933_n N_A_808_115#_M1027_g 0.0115825f $X=5.845 $Y=2.84
+ $X2=6.305 $Y2=4.195
cc_659 N_A_428_89#_c_935_n N_A_808_115#_M1027_g 0.00278359f $X=5.845 $Y=1.99
+ $X2=6.305 $Y2=4.195
cc_660 N_A_428_89#_c_947_n N_A_808_115#_M1027_g 0.00343288f $X=5.845 $Y=2.925
+ $X2=6.305 $Y2=4.195
cc_661 N_A_428_89#_c_928_n N_A_808_115#_c_1266_n 0.00153999f $X=5.57 $Y=0.865
+ $X2=6.305 $Y2=1.59
cc_662 N_A_428_89#_c_932_n N_A_808_115#_c_1266_n 0.00153999f $X=5.57 $Y=1.905
+ $X2=6.305 $Y2=1.59
cc_663 N_A_428_89#_c_934_n N_A_808_115#_c_1266_n 5.35151e-19 $X=5.57 $Y=1.59
+ $X2=6.305 $Y2=1.59
cc_664 N_A_428_89#_c_915_n N_A_808_115#_c_1267_n 0.0124213f $X=3.89 $Y=2.04
+ $X2=3.685 $Y2=1.59
cc_665 N_A_428_89#_M1015_g N_A_808_115#_c_1267_n 0.0111407f $X=3.965 $Y=3.825
+ $X2=3.685 $Y2=1.59
cc_666 N_A_428_89#_c_922_n N_A_808_115#_c_1291_n 0.00174653f $X=4.505 $Y=1.59
+ $X2=4.095 $Y2=1.17
cc_667 N_A_428_89#_c_923_n N_A_808_115#_c_1291_n 0.00205316f $X=4.505 $Y=1.425
+ $X2=4.095 $Y2=1.17
cc_668 N_A_428_89#_c_926_n N_A_808_115#_c_1291_n 0.00436807f $X=5.485 $Y=1.59
+ $X2=4.095 $Y2=1.17
cc_669 N_A_428_89#_M1015_g N_A_808_115#_c_1308_n 0.0162544f $X=3.965 $Y=3.825
+ $X2=4.095 $Y2=2.925
cc_670 N_A_428_89#_c_934_n N_A_808_115#_c_1271_n 0.00755683f $X=5.57 $Y=1.59
+ $X2=6.1 $Y2=1.59
cc_671 N_A_428_89#_c_915_n N_A_808_115#_c_1272_n 0.00156696f $X=3.89 $Y=2.04
+ $X2=5.955 $Y2=1.59
cc_672 N_A_428_89#_c_917_n N_A_808_115#_c_1272_n 0.00244106f $X=4.37 $Y=2.04
+ $X2=5.955 $Y2=1.59
cc_673 N_A_428_89#_c_921_n N_A_808_115#_c_1272_n 5.19983e-19 $X=3.965 $Y=2.04
+ $X2=5.955 $Y2=1.59
cc_674 N_A_428_89#_c_922_n N_A_808_115#_c_1272_n 0.00455939f $X=4.505 $Y=1.59
+ $X2=5.955 $Y2=1.59
cc_675 N_A_428_89#_c_926_n N_A_808_115#_c_1272_n 0.0492477f $X=5.485 $Y=1.59
+ $X2=5.955 $Y2=1.59
cc_676 N_A_428_89#_c_934_n N_A_808_115#_c_1272_n 0.0106815f $X=5.57 $Y=1.59
+ $X2=5.955 $Y2=1.59
cc_677 N_A_428_89#_c_935_n N_A_808_115#_c_1272_n 0.00191587f $X=5.845 $Y=1.99
+ $X2=5.955 $Y2=1.59
cc_678 N_A_428_89#_c_915_n N_A_808_115#_c_1274_n 0.00120486f $X=3.89 $Y=2.04
+ $X2=3.83 $Y2=1.59
cc_679 N_A_428_89#_c_928_n N_A_808_115#_c_1275_n 0.00126742f $X=5.57 $Y=0.865
+ $X2=6.1 $Y2=1.59
cc_680 N_A_428_89#_c_932_n N_A_808_115#_c_1275_n 0.00126742f $X=5.57 $Y=1.905
+ $X2=6.1 $Y2=1.59
cc_681 N_A_970_89#_c_1112_n N_A_808_115#_M1006_g 0.0104634f $X=6.435 $Y=0.91
+ $X2=6.305 $Y2=0.835
cc_682 N_A_970_89#_c_1114_n N_A_808_115#_M1006_g 0.014817f $X=6.52 $Y=1.845
+ $X2=6.305 $Y2=0.835
cc_683 N_A_970_89#_c_1115_n N_A_808_115#_M1027_g 0.0281253f $X=6.52 $Y=4.565
+ $X2=6.305 $Y2=4.195
cc_684 N_A_970_89#_c_1120_n N_A_808_115#_M1027_g 0.00261985f $X=6.52 $Y=1.93
+ $X2=6.305 $Y2=4.195
cc_685 N_A_970_89#_c_1121_n N_A_808_115#_M1027_g 0.0130428f $X=7.425 $Y=1.93
+ $X2=6.305 $Y2=4.195
cc_686 N_A_970_89#_c_1117_n N_A_808_115#_c_1266_n 0.00333003f $X=6.09 $Y=0.74
+ $X2=6.305 $Y2=1.59
cc_687 N_A_970_89#_c_1121_n N_A_808_115#_c_1266_n 0.0041429f $X=7.425 $Y=1.93
+ $X2=6.305 $Y2=1.59
cc_688 N_A_970_89#_c_1112_n N_A_808_115#_c_1271_n 8.45088e-19 $X=6.435 $Y=0.91
+ $X2=6.1 $Y2=1.59
cc_689 N_A_970_89#_c_1114_n N_A_808_115#_c_1271_n 0.0115453f $X=6.52 $Y=1.845
+ $X2=6.1 $Y2=1.59
cc_690 N_A_970_89#_c_1117_n N_A_808_115#_c_1271_n 0.00254346f $X=6.09 $Y=0.74
+ $X2=6.1 $Y2=1.59
cc_691 N_A_970_89#_c_1121_n N_A_808_115#_c_1271_n 0.00483015f $X=7.425 $Y=1.93
+ $X2=6.1 $Y2=1.59
cc_692 N_A_970_89#_M1009_g N_A_808_115#_c_1272_n 0.00231271f $X=4.925 $Y=0.945
+ $X2=5.955 $Y2=1.59
cc_693 N_A_970_89#_c_1105_n N_A_808_115#_c_1272_n 0.00187603f $X=4.985 $Y=1.93
+ $X2=5.955 $Y2=1.59
cc_694 N_A_970_89#_c_1111_n N_A_808_115#_c_1272_n 0.00166223f $X=4.985 $Y=1.93
+ $X2=5.955 $Y2=1.59
cc_695 N_A_970_89#_c_1121_n N_A_808_115#_c_1272_n 0.073586f $X=7.425 $Y=1.93
+ $X2=5.955 $Y2=1.59
cc_696 N_A_970_89#_c_1122_n N_A_808_115#_c_1272_n 0.0289631f $X=5.13 $Y=1.93
+ $X2=5.955 $Y2=1.59
cc_697 N_A_970_89#_c_1114_n N_A_808_115#_c_1275_n 0.00389142f $X=6.52 $Y=1.845
+ $X2=6.1 $Y2=1.59
cc_698 N_A_970_89#_c_1121_n N_A_808_115#_c_1275_n 0.0291144f $X=7.425 $Y=1.93
+ $X2=6.1 $Y2=1.59
cc_699 N_A_970_89#_M1010_g N_QN_M1028_g 0.0302686f $X=7.685 $Y=0.835 $X2=8.115
+ $Y2=0.835
cc_700 N_A_970_89#_c_1107_n N_QN_M1028_g 0.0153129f $X=7.572 $Y=1.765 $X2=8.115
+ $Y2=0.835
cc_701 N_A_970_89#_c_1116_n N_QN_M1028_g 4.79563e-19 $X=7.57 $Y=1.93 $X2=8.115
+ $Y2=0.835
cc_702 N_A_970_89#_c_1109_n N_QN_M1020_g 0.0102953f $X=7.66 $Y=2.595 $X2=8.115
+ $Y2=4.195
cc_703 N_A_970_89#_c_1110_n N_QN_M1020_g 0.0669165f $X=7.66 $Y=2.745 $X2=8.115
+ $Y2=4.195
cc_704 N_A_970_89#_c_1106_n N_QN_c_1394_n 0.021196f $X=7.57 $Y=1.93 $X2=8.055
+ $Y2=2.135
cc_705 N_A_970_89#_c_1116_n N_QN_c_1394_n 3.0115e-19 $X=7.57 $Y=1.93 $X2=8.055
+ $Y2=2.135
cc_706 N_A_970_89#_c_1123_n N_QN_c_1394_n 4.60229e-19 $X=7.57 $Y=1.93 $X2=8.055
+ $Y2=2.135
cc_707 N_A_970_89#_M1010_g N_QN_c_1395_n 0.0124316f $X=7.685 $Y=0.835 $X2=7.47
+ $Y2=0.74
cc_708 N_A_970_89#_c_1108_n N_QN_c_1395_n 0.00339046f $X=7.66 $Y=1.54 $X2=7.47
+ $Y2=0.74
cc_709 N_A_970_89#_M1029_g N_QN_c_1399_n 0.041548f $X=7.685 $Y=4.195 $X2=7.47
+ $Y2=2.7
cc_710 N_A_970_89#_c_1109_n N_QN_c_1399_n 0.00567875f $X=7.66 $Y=2.595 $X2=7.47
+ $Y2=2.7
cc_711 N_A_970_89#_c_1107_n N_QN_c_1400_n 0.00799433f $X=7.572 $Y=1.765 $X2=7.97
+ $Y2=1.59
cc_712 N_A_970_89#_c_1108_n N_QN_c_1400_n 0.0108908f $X=7.66 $Y=1.54 $X2=7.97
+ $Y2=1.59
cc_713 N_A_970_89#_c_1116_n N_QN_c_1400_n 0.0110498f $X=7.57 $Y=1.93 $X2=7.97
+ $Y2=1.59
cc_714 N_A_970_89#_c_1123_n N_QN_c_1400_n 0.00387586f $X=7.57 $Y=1.93 $X2=7.97
+ $Y2=1.59
cc_715 N_A_970_89#_c_1106_n N_QN_c_1402_n 0.00308111f $X=7.57 $Y=1.93 $X2=7.555
+ $Y2=1.59
cc_716 N_A_970_89#_c_1116_n N_QN_c_1402_n 0.0120703f $X=7.57 $Y=1.93 $X2=7.555
+ $Y2=1.59
cc_717 N_A_970_89#_c_1121_n N_QN_c_1402_n 0.0010572f $X=7.425 $Y=1.93 $X2=7.555
+ $Y2=1.59
cc_718 N_A_970_89#_c_1123_n N_QN_c_1402_n 0.00336135f $X=7.57 $Y=1.93 $X2=7.555
+ $Y2=1.59
cc_719 N_A_970_89#_c_1109_n N_QN_c_1403_n 0.016126f $X=7.66 $Y=2.595 $X2=7.97
+ $Y2=2.505
cc_720 N_A_970_89#_c_1110_n N_QN_c_1403_n 0.00248624f $X=7.66 $Y=2.745 $X2=7.97
+ $Y2=2.505
cc_721 N_A_970_89#_c_1116_n N_QN_c_1403_n 0.00426371f $X=7.57 $Y=1.93 $X2=7.97
+ $Y2=2.505
cc_722 N_A_970_89#_c_1123_n N_QN_c_1403_n 0.00253233f $X=7.57 $Y=1.93 $X2=7.97
+ $Y2=2.505
cc_723 N_A_970_89#_c_1106_n N_QN_c_1404_n 0.00265611f $X=7.57 $Y=1.93 $X2=7.555
+ $Y2=2.505
cc_724 N_A_970_89#_c_1116_n N_QN_c_1404_n 0.00471962f $X=7.57 $Y=1.93 $X2=7.555
+ $Y2=2.505
cc_725 N_A_970_89#_c_1121_n N_QN_c_1404_n 9.40773e-19 $X=7.425 $Y=1.93 $X2=7.555
+ $Y2=2.505
cc_726 N_A_970_89#_c_1123_n N_QN_c_1404_n 0.00140341f $X=7.57 $Y=1.93 $X2=7.555
+ $Y2=2.505
cc_727 N_A_970_89#_c_1106_n N_QN_c_1405_n 0.00216137f $X=7.57 $Y=1.93 $X2=8.055
+ $Y2=2.135
cc_728 N_A_970_89#_c_1107_n N_QN_c_1405_n 0.00323473f $X=7.572 $Y=1.765
+ $X2=8.055 $Y2=2.135
cc_729 N_A_970_89#_c_1109_n N_QN_c_1405_n 0.00226435f $X=7.66 $Y=2.595 $X2=8.055
+ $Y2=2.135
cc_730 N_A_970_89#_c_1116_n N_QN_c_1405_n 0.00987106f $X=7.57 $Y=1.93 $X2=8.055
+ $Y2=2.135
cc_731 N_A_970_89#_c_1123_n N_QN_c_1405_n 0.00377439f $X=7.57 $Y=1.93 $X2=8.055
+ $Y2=2.135
cc_732 N_A_970_89#_M1029_g QN 0.00233857f $X=7.685 $Y=4.195 $X2=7.475 $Y2=2.7
cc_733 N_A_970_89#_c_1110_n QN 0.00508004f $X=7.66 $Y=2.745 $X2=7.475 $Y2=2.7
cc_734 N_A_970_89#_c_1115_n QN 0.00570662f $X=6.52 $Y=4.565 $X2=7.475 $Y2=2.7
cc_735 N_A_970_89#_c_1116_n QN 0.00359685f $X=7.57 $Y=1.93 $X2=7.475 $Y2=2.7
cc_736 N_A_970_89#_c_1123_n QN 0.00842298f $X=7.57 $Y=1.93 $X2=7.475 $Y2=2.7
cc_737 N_A_970_89#_M1029_g Q 0.0011399f $X=7.685 $Y=4.195 $X2=8.325 $Y2=3.07
cc_738 N_A_970_89#_c_1112_n A_1276_115# 0.00176584f $X=6.435 $Y=0.91 $X2=6.38
+ $Y2=0.575
cc_739 N_A_808_115#_c_1308_n A_736_565# 0.00342591f $X=4.095 $Y=2.925 $X2=3.68
+ $Y2=2.825
cc_740 N_A_808_115#_c_1336_n A_736_565# 0.00144354f $X=3.77 $Y=2.925 $X2=3.68
+ $Y2=2.825
cc_741 N_A_808_115#_c_1267_n A_736_115# 9.4749e-19 $X=3.685 $Y=1.59 $X2=3.68
+ $Y2=0.575
cc_742 N_A_808_115#_c_1291_n A_736_115# 0.00337089f $X=4.095 $Y=1.17 $X2=3.68
+ $Y2=0.575
cc_743 N_A_808_115#_c_1292_n A_736_115# 0.00148865f $X=3.77 $Y=1.17 $X2=3.68
+ $Y2=0.575
cc_744 N_QN_M1028_g N_Q_c_1479_n 0.00595603f $X=8.115 $Y=0.835 $X2=8.33 $Y2=0.74
cc_745 N_QN_M1020_g N_Q_c_1483_n 0.0258599f $X=8.115 $Y=4.195 $X2=8.33 $Y2=4.225
cc_746 N_QN_M1028_g N_Q_c_1481_n 0.0383548f $X=8.115 $Y=0.835 $X2=8.445 $Y2=2.9
cc_747 N_QN_c_1400_n N_Q_c_1481_n 0.0111776f $X=7.97 $Y=1.59 $X2=8.445 $Y2=2.9
cc_748 N_QN_c_1403_n N_Q_c_1481_n 0.0111776f $X=7.97 $Y=2.505 $X2=8.445 $Y2=2.9
cc_749 N_QN_c_1405_n N_Q_c_1481_n 0.0438362f $X=8.055 $Y=2.135 $X2=8.445 $Y2=2.9
cc_750 N_QN_M1028_g N_Q_c_1482_n 0.00695117f $X=8.115 $Y=0.835 $X2=8.445
+ $Y2=1.255
cc_751 N_QN_M1020_g N_Q_c_1487_n 0.00911548f $X=8.115 $Y=4.195 $X2=8.33
+ $Y2=3.027
cc_752 N_QN_M1020_g Q 0.0145232f $X=8.115 $Y=4.195 $X2=8.325 $Y2=3.07
cc_753 N_QN_c_1399_n Q 0.00553023f $X=7.47 $Y=2.7 $X2=8.325 $Y2=3.07
cc_754 N_QN_c_1403_n Q 0.00245821f $X=7.97 $Y=2.505 $X2=8.325 $Y2=3.07
