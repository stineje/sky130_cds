* File: sky130_osu_sc_18T_hs__or2_2.pex.spice
* Created: Fri Nov 12 13:52:30 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__OR2_2%GND 1 2 3 31 35 37 44 46 54 64 66
r43 64 66 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r44 52 54 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r45 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r46 46 52 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.305
r47 42 60 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r48 42 44 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r49 37 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r50 33 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r51 31 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r52 31 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r53 31 33 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r54 31 38 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r55 31 46 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r56 31 47 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r57 31 37 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r58 31 38 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r59 3 54 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r60 2 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r61 1 35 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_2%VDD 1 2 21 23 32 36 43 49 53
r30 49 53 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r31 43 46 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r32 41 46 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r33 39 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.47 $X2=1.7
+ $Y2=6.47
r34 37 47 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r35 37 39 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r36 36 41 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.98 $Y2=6.355
r37 36 39 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r38 32 35 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=5.835
r39 30 47 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r40 30 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r41 25 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r42 25 29 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r43 23 47 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r44 23 29 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r45 21 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r46 21 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r47 21 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r48 2 46 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r49 2 43 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r50 1 35 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r51 1 32 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_2%B 3 7 12 15 21
r28 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.96
+ $X2=0.27 $Y2=2.96
r29 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.675
+ $X2=0.27 $Y2=2.96
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.675 $X2=0.27 $Y2=2.675
r31 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.675
+ $X2=0.475 $Y2=2.675
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.84
+ $X2=0.475 $Y2=2.675
r33 5 7 894.777 $w=1.5e-07 $l=1.745e-06 $layer=POLY_cond $X=0.475 $Y=2.84
+ $X2=0.475 $Y2=4.585
r34 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.51
+ $X2=0.475 $Y2=2.675
r35 1 3 735.819 $w=1.5e-07 $l=1.435e-06 $layer=POLY_cond $X=0.475 $Y=2.51
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_2%A 3 7 10 14 20
c44 7 0 1.37149e-19 $X=0.905 $Y=4.585
r45 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=3.33
+ $X2=0.95 $Y2=3.33
r46 14 17 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=3.33
r47 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.385 $X2=0.95 $Y2=2.385
r48 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=2.55
r49 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=2.22
r50 7 12 1043.48 $w=1.5e-07 $l=2.035e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.55
r51 3 11 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.22
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_2%A_27_617# 1 3 11 13 15 17 18 22 24 26 27
+ 31 35 39 40 42 45 49 51
r87 47 51 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.935
+ $X2=0.65 $Y2=1.935
r88 47 49 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.935
+ $X2=1.43 $Y2=1.935
r89 43 51 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.65 $Y2=1.935
r90 43 45 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=0.825
r91 41 51 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.65 $Y2=1.935
r92 41 42 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r93 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.63
+ $X2=0.61 $Y2=3.545
r94 39 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.63
+ $X2=0.345 $Y2=3.63
r95 35 37 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.26 $Y=3.795
+ $X2=0.26 $Y2=5.835
r96 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.715
+ $X2=0.345 $Y2=3.63
r97 33 35 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=3.715 $X2=0.26
+ $Y2=3.795
r98 31 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r99 29 31 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.935 $X2=1.43
+ $Y2=1.935
r100 28 29 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.935
+ $X2=1.37 $Y2=1.935
r101 24 26 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r102 20 31 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.43 $Y2=1.935
r103 20 22 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r104 19 27 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.885
+ $X2=1.352 $Y2=2.885
r105 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.96
r106 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.445 $Y2=2.885
r107 17 27 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.81
+ $X2=1.352 $Y2=2.885
r108 16 29 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=1.935
r109 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=2.81
r110 13 27 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.352 $Y2=2.885
r111 13 15 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r112 9 28 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.935
r113 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r114 3 37 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=0.135 $Y=3.085 $X2=0.26 $Y2=5.835
r115 3 35 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=0.135 $Y=3.085 $X2=0.26 $Y2=3.795
r116 1 45 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_2%Y 1 3 10 16 26 29 32
c41 16 0 1.37149e-19 $X=1.55 $Y=2.59
r42 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r43 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r44 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r45 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r46 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r47 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r48 16 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r49 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r50 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r51 3 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r52 3 19 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r53 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

