* File: sky130_osu_sc_12T_hs__and2_1.spice
* Created: Fri Nov 12 15:06:44 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__and2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_1  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_B_M1002_g A_110_115# N_GND_M1003_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.09625 PD=1.63 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_B_M1004_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_VDD_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9449 P=7.95
pX7_noxref noxref_8 A A PROBETYPE=1
pX8_noxref noxref_9 B B PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_1.pxi.spice"
*
.ends
*
*
