* File: sky130_osu_sc_18T_ms__tbufi_l.pex.spice
* Created: Fri Nov 12 14:06:52 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%GND 1 17 19 26 35 38
r35 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r36 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r37 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r38 24 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r39 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r40 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r41 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r42 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r43 1 26 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%VDD 1 13 15 21 27 31 34
r21 31 34 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r22 27 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r23 25 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r24 25 27 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507 $X2=1.02
+ $Y2=6.507
r25 21 24 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=4.475
+ $X2=0.69 $Y2=5.835
r26 19 29 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r27 19 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r28 15 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r29 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r30 13 27 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r31 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r32 1 24 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=5.835
r33 1 21 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%OE 2 5 9 13 17 22 25 32 35
c62 32 0 2.60266e-19 $X=0.69 $Y=1.85
r63 29 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.965
+ $X2=0.69 $Y2=1.85
r64 29 35 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=0.69 $Y=1.965
+ $X2=0.69 $Y2=2.845
r65 25 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=1.85
r66 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.85 $X2=0.69 $Y2=1.85
r67 15 17 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.935
+ $X2=0.475 $Y2=2.935
r68 11 22 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.905 $Y=1.65
+ $X2=0.69 $Y2=1.832
r69 11 13 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=1.65
+ $X2=0.905 $Y2=0.945
r70 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.475 $Y2=2.935
r71 7 9 1063.99 $w=1.5e-07 $l=2.075e-06 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.475 $Y2=5.085
r72 3 22 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.69 $Y2=1.832
r73 3 5 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=1.65 $X2=0.475
+ $Y2=0.945
r74 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.86 $X2=0.27
+ $Y2=2.935
r75 1 3 44.3094 $w=2.23e-07 $l=2.69768e-07 $layer=POLY_cond $X=0.27 $Y=1.8
+ $X2=0.475 $Y2=1.65
r76 1 2 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.8 $X2=0.27
+ $Y2=2.86
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%A_27_115# 1 3 11 16 20 24 28 30 33
r50 29 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.48
+ $X2=0.26 $Y2=2.48
r51 28 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.48
+ $X2=0.8 $Y2=2.48
r52 28 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=2.48
+ $X2=0.345 $Y2=2.48
r53 24 26 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=4.475
+ $X2=0.26 $Y2=5.835
r54 22 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.565
+ $X2=0.26 $Y2=2.48
r55 22 24 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=0.26 $Y=2.565
+ $X2=0.26 $Y2=4.475
r56 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.395
+ $X2=0.26 $Y2=2.48
r57 18 20 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=0.26 $Y=2.395
+ $X2=0.26 $Y2=0.825
r58 14 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=2.48 $X2=0.8 $Y2=2.48
r59 14 16 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.8 $Y=2.48
+ $X2=0.905 $Y2=2.48
r60 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.645
+ $X2=0.905 $Y2=2.48
r61 9 11 1251.15 $w=1.5e-07 $l=2.44e-06 $layer=POLY_cond $X=0.905 $Y=2.645
+ $X2=0.905 $Y2=5.085
r62 3 26 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=5.835
r63 3 24 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=4.475
r64 1 20 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%A 3 7 10 15 20 23
c46 10 0 1.90743e-19 $X=1.325 $Y=2.09
c47 3 0 6.95226e-20 $X=1.265 $Y=0.945
r48 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=2.09
+ $X2=1.325 $Y2=2.09
r49 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=3.33
+ $X2=1.14 $Y2=3.33
r50 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.175
+ $X2=1.14 $Y2=2.09
r51 13 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=2.175
+ $X2=1.14 $Y2=3.33
r52 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.09 $X2=1.325 $Y2=2.09
r53 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.09
+ $X2=1.325 $Y2=2.255
r54 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.09
+ $X2=1.325 $Y2=1.925
r55 7 12 1451.13 $w=1.5e-07 $l=2.83e-06 $layer=POLY_cond $X=1.265 $Y=5.085
+ $X2=1.265 $Y2=2.255
r56 3 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.265 $Y=0.945
+ $X2=1.265 $Y2=1.925
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__TBUFI_L%Y 1 3 10 16 26 29 32
r34 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.475
+ $X2=1.48 $Y2=2.59
r35 24 26 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.475
+ $X2=1.48 $Y2=1.82
r36 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.595
+ $X2=1.48 $Y2=1.48
r37 23 26 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.595
+ $X2=1.48 $Y2=1.82
r38 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.48 $Y=4.475
+ $X2=1.48 $Y2=5.835
r39 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.59
+ $X2=1.48 $Y2=2.59
r40 16 19 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=1.48 $Y=2.59
+ $X2=1.48 $Y2=4.475
r41 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.48
+ $X2=1.48 $Y2=1.48
r42 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.48 $Y=0.825
+ $X2=1.48 $Y2=1.48
r43 3 21 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=4.085 $X2=1.48 $Y2=5.835
r44 3 19 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=4.085 $X2=1.48 $Y2=4.475
r45 1 10 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.825
.ends

