* File: sky130_osu_sc_18T_ms__dffsr_1.pex.spice
* Created: Thu Oct 29 17:29:21 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%GND 1 2 3 4 5 6 7 8 9 88 92 94 101 103
+ 113 119 121 131 133 143 145 152 154 164 166 173 192 194
c248 152 0 1.63226e-19 $X=7.47 $Y=0.825
c249 143 0 1.67294e-19 $X=6.52 $Y=0.825
c250 119 0 3.07193e-19 $X=3.02 $Y=0.825
c251 113 0 2.98797e-19 $X=2.5 $Y=0.825
c252 101 0 1.90798e-19 $X=1.22 $Y=0.825
c253 88 0 1.91032e-19 $X=-0.05 $Y=0
r254 192 194 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.855 $Y2=0.152
r255 186 187 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=0.152
+ $X2=9.71 $Y2=0.152
r256 171 187 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.152
r257 171 173 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.825
r258 167 185 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.152
+ $X2=8.75 $Y2=0.152
r259 166 187 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=0.152
+ $X2=9.71 $Y2=0.152
r260 162 185 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.152
r261 162 164 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.825
r262 155 184 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.152
+ $X2=7.47 $Y2=0.152
r263 154 185 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.152
+ $X2=8.75 $Y2=0.152
r264 150 184 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.152
r265 150 152 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.825
r266 145 184 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=0.152
+ $X2=7.47 $Y2=0.152
r267 141 143 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.52 $Y=0.305
+ $X2=6.52 $Y2=0.825
r268 134 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.152
+ $X2=4.77 $Y2=0.152
r269 129 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.152
r270 129 131 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.825
r271 121 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.152
+ $X2=4.77 $Y2=0.152
r272 117 119 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.02 $Y=0.305
+ $X2=3.02 $Y2=0.825
r273 116 176 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.152
+ $X2=2.5 $Y2=0.152
r274 115 116 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=2.935 $Y=0.152
+ $X2=2.585 $Y2=0.152
r275 111 176 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.152
r276 111 113 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.825
r277 104 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0.152
+ $X2=1.22 $Y2=0.152
r278 103 176 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.152
+ $X2=2.5 $Y2=0.152
r279 99 175 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.152
r280 99 101 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.825
r281 94 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.152
+ $X2=1.22 $Y2=0.152
r282 90 92 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r283 88 90 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r284 88 95 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r285 88 186 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.855 $Y=0.152 $X2=9.795
+ $Y2=0.152
r286 88 194 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=0.17
+ $X2=9.855 $Y2=0.17
r287 88 192 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=0.17
+ $X2=0.335 $Y2=0.17
r288 88 141 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.52 $Y2=0.305
r289 88 133 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.435 $Y2=0.152
r290 88 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.605 $Y2=0.152
r291 88 117 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.02 $Y2=0.305
r292 88 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=2.935 $Y2=0.152
r293 88 122 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.105 $Y2=0.152
r294 88 166 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=9.625 $Y2=0.152
r295 88 167 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.835 $Y2=0.152
r296 88 154 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.665 $Y2=0.152
r297 88 155 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=7.815 $Y=0.152
+ $X2=7.555 $Y2=0.152
r298 88 145 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.385 $Y2=0.152
r299 88 146 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.605 $Y2=0.152
r300 88 133 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.435 $Y2=0.152
r301 88 134 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.855 $Y2=0.152
r302 88 121 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=4.685 $Y2=0.152
r303 88 122 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.105 $Y2=0.152
r304 88 103 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.415 $Y2=0.152
r305 88 104 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.305 $Y2=0.152
r306 88 94 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.135 $Y2=0.152
r307 88 95 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r308 9 173 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=9.57
+ $Y=0.575 $X2=9.71 $Y2=0.825
r309 8 164 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.61
+ $Y=0.575 $X2=8.75 $Y2=0.825
r310 7 152 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.825
r311 6 143 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.825
r312 5 131 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.575 $X2=4.77 $Y2=0.825
r313 4 119 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.575 $X2=3.02 $Y2=0.825
r314 3 113 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.5 $Y2=0.825
r315 2 101 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.575 $X2=1.22 $Y2=0.825
r316 1 92 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%VDD 1 2 3 4 5 6 7 67 71 75 83 87 93 97
+ 105 109 117 121 127 131 139 154 159 163
c145 139 0 1.98165e-19 $X=9.71 $Y=3.455
r146 159 163 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=6.49
+ $X2=9.855 $Y2=6.49
r147 154 159 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=6.507
+ $X2=9.855 $Y2=6.507
r148 154 157 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=6.49
+ $X2=0.335 $Y2=6.49
r149 151 163 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.795 $Y=6.507
+ $X2=9.855 $Y2=6.507
r150 151 152 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=6.507
+ $X2=9.71 $Y2=6.507
r151 139 142 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=9.71 $Y=3.455
+ $X2=9.71 $Y2=5.835
r152 137 152 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.71 $Y=6.355
+ $X2=9.71 $Y2=6.507
r153 137 142 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.71 $Y=6.355
+ $X2=9.71 $Y2=5.835
r154 134 136 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=8.495 $Y=6.507
+ $X2=9.175 $Y2=6.507
r155 132 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=6.507
+ $X2=7.9 $Y2=6.507
r156 132 134 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=7.985 $Y=6.507
+ $X2=8.495 $Y2=6.507
r157 131 152 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=6.507
+ $X2=9.71 $Y2=6.507
r158 131 136 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.625 $Y=6.507
+ $X2=9.175 $Y2=6.507
r159 127 130 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=5.835
r160 125 150 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=6.507
r161 125 130 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=5.835
r162 122 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=6.507
+ $X2=6.52 $Y2=6.507
r163 122 124 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=6.605 $Y=6.507
+ $X2=7.135 $Y2=6.507
r164 121 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.9 $Y2=6.507
r165 121 124 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.135 $Y2=6.507
r166 117 120 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.52 $Y=3.455
+ $X2=6.52 $Y2=5.835
r167 115 148 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.52 $Y=6.355
+ $X2=6.52 $Y2=6.507
r168 115 120 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.52 $Y=6.355
+ $X2=6.52 $Y2=5.835
r169 112 114 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=6.507
+ $X2=5.775 $Y2=6.507
r170 110 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=6.507
+ $X2=4.77 $Y2=6.507
r171 110 112 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=4.855 $Y=6.507
+ $X2=5.095 $Y2=6.507
r172 109 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=6.507
+ $X2=6.52 $Y2=6.507
r173 109 114 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=6.435 $Y=6.507
+ $X2=5.775 $Y2=6.507
r174 105 108 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.77 $Y=3.795
+ $X2=4.77 $Y2=5.835
r175 103 146 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.77 $Y=6.355
+ $X2=4.77 $Y2=6.507
r176 103 108 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.77 $Y=6.355
+ $X2=4.77 $Y2=5.835
r177 100 102 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=6.507
+ $X2=4.415 $Y2=6.507
r178 98 145 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=6.507
+ $X2=3.02 $Y2=6.507
r179 98 100 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.105 $Y=6.507
+ $X2=3.735 $Y2=6.507
r180 97 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=6.507
+ $X2=4.77 $Y2=6.507
r181 97 102 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.685 $Y=6.507
+ $X2=4.415 $Y2=6.507
r182 93 96 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=3.02 $Y=3.795
+ $X2=3.02 $Y2=5.835
r183 91 145 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.02 $Y=6.355
+ $X2=3.02 $Y2=6.507
r184 91 96 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.02 $Y=6.355
+ $X2=3.02 $Y2=5.835
r185 88 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=6.507
+ $X2=2.07 $Y2=6.507
r186 88 90 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.155 $Y=6.507
+ $X2=2.375 $Y2=6.507
r187 87 145 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=6.507
+ $X2=3.02 $Y2=6.507
r188 87 90 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=2.935 $Y=6.507
+ $X2=2.375 $Y2=6.507
r189 83 86 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.07 $Y=4.135
+ $X2=2.07 $Y2=5.835
r190 81 143 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.07 $Y=6.355
+ $X2=2.07 $Y2=6.507
r191 81 86 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.07 $Y=6.355
+ $X2=2.07 $Y2=5.835
r192 78 80 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=6.507
+ $X2=1.695 $Y2=6.507
r193 76 157 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r194 76 78 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.015 $Y2=6.507
r195 75 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=6.507
+ $X2=2.07 $Y2=6.507
r196 75 80 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.985 $Y=6.507
+ $X2=1.695 $Y2=6.507
r197 71 74 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r198 69 157 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r199 69 74 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r200 67 157 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=6.355 $X2=0.335 $Y2=6.44
r201 67 163 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=9.65 $Y=6.355 $X2=9.855 $Y2=6.44
r202 67 150 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=6.355 $X2=7.815 $Y2=6.44
r203 67 148 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=6.355 $X2=6.455 $Y2=6.44
r204 67 145 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=6.355 $X2=3.055 $Y2=6.44
r205 67 136 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=6.355 $X2=9.175 $Y2=6.44
r206 67 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=6.355 $X2=8.495 $Y2=6.44
r207 67 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=6.355 $X2=7.135 $Y2=6.44
r208 67 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=6.355 $X2=5.775 $Y2=6.44
r209 67 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=6.355 $X2=5.095 $Y2=6.44
r210 67 102 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=6.355 $X2=4.415 $Y2=6.44
r211 67 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=6.355 $X2=3.735 $Y2=6.44
r212 67 90 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=6.355 $X2=2.375 $Y2=6.44
r213 67 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=6.355 $X2=1.695 $Y2=6.44
r214 67 78 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=6.355 $X2=1.015 $Y2=6.44
r215 7 142 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=9.57
+ $Y=3.085 $X2=9.71 $Y2=5.835
r216 7 139 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=9.57
+ $Y=3.085 $X2=9.71 $Y2=3.455
r217 6 130 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=7.76
+ $Y=3.085 $X2=7.9 $Y2=5.835
r218 6 127 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=7.76
+ $Y=3.085 $X2=7.9 $Y2=4.135
r219 5 120 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=5.835
r220 5 117 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=3.455
r221 4 108 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=4.63 $Y=3.085 $X2=4.77 $Y2=5.835
r222 4 105 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=4.63 $Y=3.085 $X2=4.77 $Y2=3.795
r223 3 96 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=2.895 $Y=3.085 $X2=3.02 $Y2=5.835
r224 3 93 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=2.895 $Y=3.085 $X2=3.02 $Y2=3.795
r225 2 86 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=5.835
r226 2 83 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=4.135
r227 1 74 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r228 1 71 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%RN 3 5 7 9 16 17
c40 17 0 7.48684e-20 $X=0.325 $Y=3.33
c41 3 0 1.63751e-20 $X=0.475 $Y=1.075
r42 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=2.305 $X2=0.53 $Y2=2.305
r44 10 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=2.47 $X2=0.32
+ $Y2=3.33
r45 9 12 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=2.305
+ $X2=0.53 $Y2=2.305
r46 9 10 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.305
+ $X2=0.32 $Y2=2.47
r47 5 13 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.53 $Y2=2.305
r48 5 7 1084.5 $w=1.5e-07 $l=2.115e-06 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=4.585
r49 1 13 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.53 $Y2=2.305
r50 1 3 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_110_115# 1 2 8 11 13 15 16 18 21 24
+ 27 29 33 37 42 43 44 50 52 53 59 60 63 65 68
c207 53 0 1.63751e-20 $X=1.375 $Y=1.48
c208 50 0 7.48684e-20 $X=0.87 $Y=2.74
c209 43 0 1.90798e-19 $X=1.145 $Y=1.59
c210 29 0 1.09867e-19 $X=8.545 $Y=2.75
c211 24 0 1.70295e-19 $X=8.8 $Y=2.605
r212 68 71 12.05 $w=2.4e-07 $l=6e-08 $layer=POLY_cond $X=8.8 $Y=1.59 $X2=8.86
+ $Y2=1.59
r213 64 65 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.23 $Y=1.59 $X2=1.29
+ $Y2=1.59
r214 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.59 $X2=1.23 $Y2=1.59
r215 60 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.86
+ $Y=1.59 $X2=8.86 $Y2=1.59
r216 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.86 $Y=1.48
+ $X2=8.86 $Y2=1.48
r217 56 63 6.15596 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=1.27 $Y=1.48
+ $X2=1.27 $Y2=1.59
r218 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.48
+ $X2=1.23 $Y2=1.48
r219 53 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.375 $Y=1.48
+ $X2=1.23 $Y2=1.48
r220 52 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.715 $Y=1.48
+ $X2=8.86 $Y2=1.48
r221 52 53 7.06756 $w=1.7e-07 $l=7.34e-06 $layer=MET1_cond $X=8.715 $Y=1.48
+ $X2=1.375 $Y2=1.48
r222 48 50 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.74
+ $X2=0.87 $Y2=2.74
r223 45 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.87 $Y2=1.59
r224 44 47 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.59
+ $X2=0.87 $Y2=1.59
r225 43 63 2.19618 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=1.27 $Y2=1.59
r226 43 44 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=0.955 $Y2=1.59
r227 42 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.655
+ $X2=0.87 $Y2=2.74
r228 41 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=1.59
r229 41 42 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=2.655
r230 37 39 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r231 35 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=2.74
r232 35 37 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=3.455
r233 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=1.59
r234 31 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=0.825
r235 29 30 60.25 $w=2.04e-07 $l=2.55e-07 $layer=POLY_cond $X=8.545 $Y=2.75
+ $X2=8.8 $Y2=2.75
r236 25 27 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.29 $Y=2.82
+ $X2=1.425 $Y2=2.82
r237 24 30 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.8 $Y=2.605
+ $X2=8.8 $Y2=2.75
r238 23 68 13.7767 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=1.755
+ $X2=8.8 $Y2=1.59
r239 23 24 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=8.8 $Y=1.755
+ $X2=8.8 $Y2=2.605
r240 19 29 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.545 $Y=2.895
+ $X2=8.545 $Y2=2.75
r241 19 21 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=8.545 $Y=2.895
+ $X2=8.545 $Y2=4.585
r242 16 68 53.2208 $w=2.4e-07 $l=3.37565e-07 $layer=POLY_cond $X=8.535 $Y=1.425
+ $X2=8.8 $Y2=1.59
r243 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.535 $Y=1.425
+ $X2=8.535 $Y2=0.945
r244 13 65 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.435 $Y=1.425
+ $X2=1.29 $Y2=1.59
r245 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.435 $Y=1.425
+ $X2=1.435 $Y2=0.945
r246 9 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=2.895
+ $X2=1.425 $Y2=2.82
r247 9 11 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=1.425 $Y=2.895
+ $X2=1.425 $Y2=4.585
r248 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=2.745
+ $X2=1.29 $Y2=2.82
r249 7 65 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.755
+ $X2=1.29 $Y2=1.59
r250 7 8 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=1.29 $Y=1.755
+ $X2=1.29 $Y2=2.745
r251 2 39 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r252 2 37 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r253 1 33 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%SN 1 2 5 9 13 17 22 29 30 32 33 36 39
+ 41 45
c172 33 0 2.97185e-19 $X=1.855 $Y=2.96
r173 45 46 5.53115 $w=3.05e-07 $l=3.5e-08 $layer=POLY_cond $X=1.855 $Y=2.37
+ $X2=1.89 $Y2=2.37
r174 39 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.935 $Y=2.96
+ $X2=7.935 $Y2=2.96
r175 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=2.96
+ $X2=1.71 $Y2=2.96
r176 33 35 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=2.96
+ $X2=1.71 $Y2=2.96
r177 32 39 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.79 $Y=2.96
+ $X2=7.935 $Y2=2.96
r178 32 33 5.71471 $w=1.7e-07 $l=5.935e-06 $layer=MET1_cond $X=7.79 $Y=2.96
+ $X2=1.855 $Y2=2.96
r179 30 49 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=2.255
+ $X2=8.035 $Y2=2.42
r180 30 48 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=2.255
+ $X2=8.035 $Y2=2.09
r181 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.025
+ $Y=2.255 $X2=8.025 $Y2=2.255
r182 26 41 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.935 $Y=2.42
+ $X2=7.935 $Y2=2.96
r183 25 29 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=8.025 $Y2=2.295
r184 25 26 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=7.935 $Y2=2.42
r185 23 45 22.9148 $w=3.05e-07 $l=1.45e-07 $layer=POLY_cond $X=1.71 $Y=2.37
+ $X2=1.855 $Y2=2.37
r186 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=2.37 $X2=1.71 $Y2=2.37
r187 20 36 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.71 $Y=2.455
+ $X2=1.71 $Y2=2.96
r188 20 22 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.455
+ $X2=1.71 $Y2=2.37
r189 17 49 1110.14 $w=1.5e-07 $l=2.165e-06 $layer=POLY_cond $X=8.115 $Y=4.585
+ $X2=8.115 $Y2=2.42
r190 13 48 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=8.045 $Y=1.075
+ $X2=8.045 $Y2=2.09
r191 9 19 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=1.925 $Y=1.075
+ $X2=1.925 $Y2=1.775
r192 3 45 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=2.535
+ $X2=1.855 $Y2=2.37
r193 3 5 1051.17 $w=1.5e-07 $l=2.05e-06 $layer=POLY_cond $X=1.855 $Y=2.535
+ $X2=1.855 $Y2=4.585
r194 2 46 10.4756 $w=2.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=2.205
+ $X2=1.89 $Y2=2.37
r195 1 19 38.6248 $w=2.2e-07 $l=1.1e-07 $layer=POLY_cond $X=1.89 $Y=1.885
+ $X2=1.89 $Y2=1.775
r196 1 2 93.3405 $w=2.2e-07 $l=3.2e-07 $layer=POLY_cond $X=1.89 $Y=1.885
+ $X2=1.89 $Y2=2.205
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_432_520# 1 2 9 13 18 19 20 21 22 23
+ 25 28 32 37
c90 37 0 1.71621e-19 $X=3.887 $Y=1.415
c91 20 0 1.29912e-19 $X=3.71 $Y=1.765
c92 19 0 1.52962e-19 $X=2.295 $Y=2.765
c93 13 0 1.44224e-19 $X=2.285 $Y=4.585
c94 9 0 1.32807e-19 $X=2.285 $Y=1.075
r95 36 37 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.887 $Y=1.245
+ $X2=3.887 $Y2=1.415
r96 32 34 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=3.895 $Y=3.455
+ $X2=3.895 $Y2=5.835
r97 30 32 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=3.895 $Y=3.375
+ $X2=3.895 $Y2=3.455
r98 28 36 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=3.895 $Y=0.825
+ $X2=3.895 $Y2=1.245
r99 25 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.795 $Y=1.68
+ $X2=3.795 $Y2=1.415
r100 22 30 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=3.725 $Y=3.185
+ $X2=3.895 $Y2=3.375
r101 22 23 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=3.725 $Y=3.185
+ $X2=2.38 $Y2=3.185
r102 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=1.765
+ $X2=3.795 $Y2=1.68
r103 20 21 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.71 $Y=1.765
+ $X2=2.38 $Y2=1.765
r104 19 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.765
+ $X2=2.295 $Y2=2.93
r105 19 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.765
+ $X2=2.295 $Y2=2.6
r106 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=2.765 $X2=2.295 $Y2=2.765
r107 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=3.1
+ $X2=2.38 $Y2=3.185
r108 16 18 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.295 $Y=3.1
+ $X2=2.295 $Y2=2.765
r109 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=1.85
+ $X2=2.38 $Y2=1.765
r110 15 18 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.295 $Y=1.85
+ $X2=2.295 $Y2=2.765
r111 13 40 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.285 $Y=4.585
+ $X2=2.285 $Y2=2.93
r112 9 39 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=2.285 $Y=1.075
+ $X2=2.285 $Y2=2.6
r113 2 34 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=3.67
+ $Y=3.085 $X2=3.895 $Y2=5.835
r114 2 32 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=3.67
+ $Y=3.085 $X2=3.895 $Y2=3.455
r115 1 28 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=3.67
+ $Y=0.575 $X2=3.895 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%D 3 7 10 12 16
c39 16 0 1.12321e-19 $X=3.295 $Y=2.22
c40 10 0 1.41836e-19 $X=3.295 $Y=2.22
r41 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=2.22
+ $X2=3.295 $Y2=2.385
r42 16 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=2.22
+ $X2=3.295 $Y2=2.055
r43 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=2.22 $X2=3.295 $Y2=2.22
r44 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.295 $Y=2.22
+ $X2=3.295 $Y2=2.22
r45 7 18 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=3.235 $Y=4.585
+ $X2=3.235 $Y2=2.385
r46 3 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.235 $Y=1.075
+ $X2=3.235 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%CK 3 7 10 13 17 18 20 23 24 25 26 30 31
+ 35 36 38 39 40 41 42 43 46 50 52 54 59 63 66 70
c233 63 0 1.29912e-19 $X=4.135 $Y=1.685
c234 59 0 1.41836e-19 $X=3.655 $Y=2.765
c235 39 0 6.79641e-20 $X=5.49 $Y=2.59
c236 30 0 1.98654e-19 $X=4.135 $Y=1.85
c237 26 0 1.86602e-19 $X=4.05 $Y=2.59
r238 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=2.765 $X2=6.88 $Y2=2.765
r239 70 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=2.765
+ $X2=5.885 $Y2=2.93
r240 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=2.765 $X2=5.885 $Y2=2.765
r241 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=2.765
+ $X2=3.655 $Y2=2.93
r242 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=2.765 $X2=3.655 $Y2=2.765
r243 54 74 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.88 $Y=2.59
+ $X2=6.88 $Y2=2.765
r244 52 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.88 $Y=2.59
+ $X2=6.88 $Y2=2.59
r245 50 69 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.885 $Y=2.59
+ $X2=5.885 $Y2=2.765
r246 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=2.59
+ $X2=5.885 $Y2=2.59
r247 46 58 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.655 $Y=2.59
+ $X2=3.655 $Y2=2.765
r248 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.655 $Y=2.59
+ $X2=3.655 $Y2=2.59
r249 43 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.03 $Y=2.59
+ $X2=5.885 $Y2=2.59
r250 42 52 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.735 $Y=2.59
+ $X2=6.88 $Y2=2.59
r251 42 43 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.735 $Y=2.59
+ $X2=6.03 $Y2=2.59
r252 41 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.8 $Y=2.59
+ $X2=3.655 $Y2=2.59
r253 40 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.74 $Y=2.59
+ $X2=5.885 $Y2=2.59
r254 40 41 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.74 $Y=2.59
+ $X2=3.8 $Y2=2.59
r255 38 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.59
+ $X2=5.885 $Y2=2.59
r256 38 39 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.8 $Y=2.59
+ $X2=5.49 $Y2=2.59
r257 36 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.85
+ $X2=5.405 $Y2=1.685
r258 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.85 $X2=5.405 $Y2=1.85
r259 33 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.405 $Y=2.505
+ $X2=5.49 $Y2=2.59
r260 33 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.405 $Y=2.505
+ $X2=5.405 $Y2=1.85
r261 31 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.85
+ $X2=4.135 $Y2=1.685
r262 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.85 $X2=4.135 $Y2=1.85
r263 28 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.135 $Y=2.505
+ $X2=4.135 $Y2=1.85
r264 27 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=2.59
+ $X2=3.655 $Y2=2.59
r265 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.05 $Y=2.59
+ $X2=4.135 $Y2=2.505
r266 26 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.05 $Y=2.59
+ $X2=3.74 $Y2=2.59
r267 24 25 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.762 $Y=1.685
+ $X2=6.762 $Y2=1.835
r268 23 75 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.79 $Y=2.6
+ $X2=6.837 $Y2=2.765
r269 23 25 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.79 $Y=2.6
+ $X2=6.79 $Y2=1.835
r270 18 75 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.735 $Y=2.93
+ $X2=6.837 $Y2=2.765
r271 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=6.735 $Y=2.93
+ $X2=6.735 $Y2=4.585
r272 17 24 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.735 $Y=1.075
+ $X2=6.735 $Y2=1.685
r273 13 72 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.945 $Y=4.585
+ $X2=5.945 $Y2=2.93
r274 10 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.345 $Y=1.075
+ $X2=5.345 $Y2=1.685
r275 7 63 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.195 $Y=1.075
+ $X2=4.195 $Y2=1.685
r276 3 61 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.595 $Y=4.585
+ $X2=3.595 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_217_617# 1 2 9 13 17 21 23 24 25 26
+ 29 33 34 37 41 42 48 49 56
c165 56 0 1.63226e-19 $X=1.71 $Y=0.825
c166 42 0 1.32807e-19 $X=1.855 $Y=1.85
c167 41 0 2.71143e-19 $X=4.49 $Y=1.85
c168 37 0 1.5821e-19 $X=4.725 $Y=2.765
c169 26 0 6.79641e-20 $X=4.91 $Y=2.765
c170 24 0 1.86602e-19 $X=4.63 $Y=2.765
c171 21 0 6.36774e-20 $X=4.985 $Y=4.585
c172 13 0 6.36774e-20 $X=4.555 $Y=4.585
r173 49 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=1.85 $X2=4.725 $Y2=1.85
r174 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.85
+ $X2=4.635 $Y2=1.85
r175 45 56 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=1.71 $Y=1.85
+ $X2=1.71 $Y2=0.825
r176 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.85
+ $X2=1.71 $Y2=1.85
r177 42 44 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.85
+ $X2=1.71 $Y2=1.85
r178 41 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.49 $Y=1.85
+ $X2=4.635 $Y2=1.85
r179 41 42 2.53719 $w=1.7e-07 $l=2.635e-06 $layer=MET1_cond $X=4.49 $Y=1.85
+ $X2=1.855 $Y2=1.85
r180 40 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.935
+ $X2=1.71 $Y2=1.85
r181 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=2.765 $X2=4.725 $Y2=2.765
r182 35 49 2.3025 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.725 $Y=1.935
+ $X2=4.635 $Y2=1.81
r183 35 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.725 $Y=1.935
+ $X2=4.725 $Y2=2.765
r184 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=2.02
+ $X2=1.71 $Y2=1.935
r185 33 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.625 $Y=2.02
+ $X2=1.295 $Y2=2.02
r186 29 31 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.21 $Y=3.795
+ $X2=1.21 $Y2=5.835
r187 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.295 $Y2=2.02
r188 27 29 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.21 $Y2=3.795
r189 26 38 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=2.765
+ $X2=4.725 $Y2=2.765
r190 25 53 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=1.85
+ $X2=4.725 $Y2=1.85
r191 24 38 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=2.765
+ $X2=4.725 $Y2=2.765
r192 23 53 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=1.85
+ $X2=4.725 $Y2=1.85
r193 19 26 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.985 $Y=2.9
+ $X2=4.91 $Y2=2.765
r194 19 21 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.985 $Y=2.9
+ $X2=4.985 $Y2=4.585
r195 15 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.985 $Y=1.715
+ $X2=4.91 $Y2=1.85
r196 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.985 $Y=1.715
+ $X2=4.985 $Y2=1.075
r197 11 24 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.63 $Y2=2.765
r198 11 13 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.555 $Y2=4.585
r199 7 23 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.63 $Y2=1.85
r200 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.555 $Y2=1.075
r201 2 31 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=1.085 $Y=3.085 $X2=1.21 $Y2=5.835
r202 2 29 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=1.085 $Y=3.085 $X2=1.21 $Y2=3.795
r203 1 56 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.575 $X2=1.71 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_704_89# 1 2 7 9 11 12 13 16 18 22 24
+ 27 30 33 35 36 37 40 44 47 50 55 56 59 63 66
c191 33 0 1.98654e-19 $X=3.715 $Y=1.76
c192 16 0 1.12321e-19 $X=4.195 $Y=4.585
r193 61 63 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=3.185
+ $X2=7.22 $Y2=3.185
r194 57 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=2.19
+ $X2=7.22 $Y2=2.19
r195 55 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=3.1
+ $X2=7.22 $Y2=3.185
r196 54 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.275
+ $X2=7.22 $Y2=2.19
r197 54 55 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=7.22 $Y=2.275
+ $X2=7.22 $Y2=3.1
r198 50 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.95 $Y=3.455
+ $X2=6.95 $Y2=5.835
r199 48 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=3.27
+ $X2=6.95 $Y2=3.185
r200 48 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.95 $Y=3.27
+ $X2=6.95 $Y2=3.455
r201 47 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=2.105
+ $X2=6.95 $Y2=2.19
r202 46 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.935
+ $X2=6.95 $Y2=1.85
r203 46 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.95 $Y=1.935
+ $X2=6.95 $Y2=2.105
r204 42 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.765
+ $X2=6.95 $Y2=1.85
r205 42 44 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.95 $Y=1.765
+ $X2=6.95 $Y2=0.825
r206 40 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.85
+ $X2=5.885 $Y2=2.015
r207 40 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.85
+ $X2=5.885 $Y2=1.685
r208 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=1.85 $X2=5.885 $Y2=1.85
r209 37 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=1.85
+ $X2=6.95 $Y2=1.85
r210 37 39 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.865 $Y=1.85
+ $X2=5.885 $Y2=1.85
r211 31 33 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.595 $Y=1.76
+ $X2=3.715 $Y2=1.76
r212 30 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.945 $Y=1.075
+ $X2=5.945 $Y2=1.685
r213 27 67 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.825 $Y=2.225
+ $X2=5.825 $Y2=2.015
r214 25 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=2.3
+ $X2=5.345 $Y2=2.3
r215 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.75 $Y=2.3
+ $X2=5.825 $Y2=2.225
r216 24 25 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.75 $Y=2.3
+ $X2=5.42 $Y2=2.3
r217 20 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.345 $Y=2.375
+ $X2=5.345 $Y2=2.3
r218 20 22 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=5.345 $Y=2.375
+ $X2=5.345 $Y2=4.585
r219 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=2.3
+ $X2=4.195 $Y2=2.3
r220 18 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=2.3
+ $X2=5.345 $Y2=2.3
r221 18 19 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.27 $Y=2.3 $X2=4.27
+ $Y2=2.3
r222 14 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=2.375
+ $X2=4.195 $Y2=2.3
r223 14 16 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=4.195 $Y=2.375
+ $X2=4.195 $Y2=4.585
r224 12 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=2.3
+ $X2=4.195 $Y2=2.3
r225 12 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.12 $Y=2.3
+ $X2=3.79 $Y2=2.3
r226 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=2.225
+ $X2=3.79 $Y2=2.3
r227 10 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.715 $Y=1.835
+ $X2=3.715 $Y2=1.76
r228 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.715 $Y=1.835
+ $X2=3.715 $Y2=2.225
r229 7 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.685
+ $X2=3.595 $Y2=1.76
r230 7 9 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.595 $Y=1.685
+ $X2=3.595 $Y2=1.075
r231 2 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.81
+ $Y=3.085 $X2=6.95 $Y2=5.835
r232 2 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.81
+ $Y=3.085 $X2=6.95 $Y2=3.455
r233 1 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.81
+ $Y=0.575 $X2=6.95 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_1246_89# 1 2 9 13 21 24 25 26 27 28
+ 31 35 39 42 43 46 49 50 54 59 60
c173 59 0 2.20654e-19 $X=9.38 $Y=2.19
c174 31 0 1.63226e-19 $X=8.26 $Y=0.825
c175 27 0 8.77106e-20 $X=9.47 $Y=2.855
r176 59 61 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=2.19
+ $X2=9.382 $Y2=2.355
r177 59 60 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=2.19
+ $X2=9.382 $Y2=2.025
r178 54 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=2.19
+ $X2=6.365 $Y2=2.355
r179 54 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=2.19
+ $X2=6.365 $Y2=2.025
r180 50 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.38
+ $Y=2.19 $X2=9.38 $Y2=2.19
r181 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.38 $Y=2.19
+ $X2=9.38 $Y2=2.19
r182 46 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=2.19 $X2=6.365 $Y2=2.19
r183 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.365 $Y=2.19
+ $X2=6.365 $Y2=2.19
r184 43 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.51 $Y=2.19
+ $X2=6.365 $Y2=2.19
r185 42 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.235 $Y=2.19
+ $X2=9.38 $Y2=2.19
r186 42 43 2.62385 $w=1.7e-07 $l=2.725e-06 $layer=MET1_cond $X=9.235 $Y=2.19
+ $X2=6.51 $Y2=2.19
r187 39 50 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.845 $Y=2.19
+ $X2=9.38 $Y2=2.19
r188 35 37 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=8.76 $Y=3.795
+ $X2=8.76 $Y2=5.835
r189 33 39 5.37722 $w=2.41e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=2.275
+ $X2=8.845 $Y2=2.19
r190 33 35 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=8.76 $Y=2.275
+ $X2=8.76 $Y2=3.795
r191 29 33 25.3112 $w=2.41e-07 $l=6.89202e-07 $layer=LI1_cond $X=8.26 $Y=1.825
+ $X2=8.76 $Y2=2.275
r192 29 31 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=8.26 $Y=1.825
+ $X2=8.26 $Y2=0.825
r193 27 28 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=2.855
+ $X2=9.47 $Y2=3.005
r194 27 61 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.445 $Y=2.855
+ $X2=9.445 $Y2=2.355
r195 26 60 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.445 $Y=1.8
+ $X2=9.445 $Y2=2.025
r196 25 26 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=1.65 $X2=9.47
+ $Y2=1.8
r197 24 28 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=9.495 $Y=4.585
+ $X2=9.495 $Y2=3.005
r198 21 25 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.495 $Y=1.075
+ $X2=9.495 $Y2=1.65
r199 13 56 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=6.305 $Y=4.585
+ $X2=6.305 $Y2=2.355
r200 9 55 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.305 $Y=1.075
+ $X2=6.305 $Y2=2.025
r201 2 37 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=8.62
+ $Y=3.085 $X2=8.76 $Y2=5.835
r202 2 35 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=8.62
+ $Y=3.085 $X2=8.76 $Y2=3.795
r203 1 31 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=8.12
+ $Y=0.575 $X2=8.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_1084_115# 1 2 8 9 11 14 18 20 21 22
+ 23 26 30 36 37 40 43 44 51
c157 40 0 1.57671e-19 $X=5.065 $Y=1.85
c158 37 0 1.5821e-19 $X=5.21 $Y=1.85
c159 20 0 1.67294e-19 $X=5.475 $Y=1.43
c160 14 0 6.36774e-20 $X=7.685 $Y=4.585
r161 50 51 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=2.765
+ $X2=7.685 $Y2=2.765
r162 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=2.765 $X2=7.595 $Y2=2.765
r163 46 50 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=2.765
+ $X2=7.595 $Y2=2.765
r164 44 49 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.595 $Y=1.85
+ $X2=7.595 $Y2=2.765
r165 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=1.85
+ $X2=7.595 $Y2=1.85
r166 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.065 $Y=1.85
+ $X2=5.065 $Y2=1.85
r167 37 39 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.21 $Y=1.85
+ $X2=5.065 $Y2=1.85
r168 36 43 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=1.85
+ $X2=7.595 $Y2=1.85
r169 36 37 2.15686 $w=1.7e-07 $l=2.24e-06 $layer=MET1_cond $X=7.45 $Y=1.85
+ $X2=5.21 $Y2=1.85
r170 35 40 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.065 $Y=3.1
+ $X2=5.065 $Y2=1.85
r171 34 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.065 $Y=1.515
+ $X2=5.065 $Y2=1.85
r172 30 32 69.1466 $w=3.38e-07 $l=2.04e-06 $layer=LI1_cond $X=5.645 $Y=3.795
+ $X2=5.645 $Y2=5.835
r173 28 30 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=5.645 $Y=3.27
+ $X2=5.645 $Y2=3.795
r174 24 26 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=5.645 $Y=1.345
+ $X2=5.645 $Y2=0.825
r175 23 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.15 $Y=3.185
+ $X2=5.065 $Y2=3.1
r176 22 28 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=3.185
+ $X2=5.645 $Y2=3.27
r177 22 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=3.185
+ $X2=5.15 $Y2=3.185
r178 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.15 $Y=1.43
+ $X2=5.065 $Y2=1.515
r179 20 24 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=1.43
+ $X2=5.645 $Y2=1.345
r180 20 21 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=1.43
+ $X2=5.15 $Y2=1.43
r181 16 18 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=7.505 $Y=1.77
+ $X2=7.685 $Y2=1.77
r182 12 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.685 $Y=2.9
+ $X2=7.685 $Y2=2.765
r183 12 14 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=7.685 $Y=2.9
+ $X2=7.685 $Y2=4.585
r184 9 18 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.685 $Y=1.69
+ $X2=7.685 $Y2=1.77
r185 9 11 197.62 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=7.685 $Y=1.69
+ $X2=7.685 $Y2=1.075
r186 8 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.505 $Y=2.63
+ $X2=7.505 $Y2=2.765
r187 7 16 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.505 $Y=1.85
+ $X2=7.505 $Y2=1.77
r188 7 8 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.505 $Y=1.85
+ $X2=7.505 $Y2=2.63
r189 2 32 171.429 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=3 $X=5.42
+ $Y=3.085 $X2=5.645 $Y2=5.835
r190 2 30 171.429 $w=1.7e-07 $l=8.1477e-07 $layer=licon1_PDIFF $count=3 $X=5.42
+ $Y=3.085 $X2=5.645 $Y2=3.795
r191 1 26 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=5.42
+ $Y=0.575 $X2=5.645 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%QN 1 2 9 13 17 19 20 21 22 26 27 31 32
c81 32 0 8.77106e-20 $X=9.285 $Y=2.96
c82 31 0 1.09867e-19 $X=9.28 $Y=2.96
c83 27 0 1.98165e-19 $X=9.865 $Y=2.395
c84 21 0 9.99996e-20 $X=9.78 $Y=2.765
c85 19 0 1.20654e-19 $X=9.78 $Y=1.85
c86 17 0 1.70295e-19 $X=9.28 $Y=0.825
r87 39 41 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=9.28 $Y=3.455
+ $X2=9.28 $Y2=5.835
r88 31 39 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.28 $Y=2.96
+ $X2=9.28 $Y2=3.455
r89 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=2.96
+ $X2=9.28 $Y2=2.96
r90 28 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.28 $Y=2.85
+ $X2=9.28 $Y2=2.96
r91 27 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=2.395
+ $X2=9.865 $Y2=2.56
r92 27 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=2.395
+ $X2=9.865 $Y2=2.23
r93 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.865
+ $Y=2.395 $X2=9.865 $Y2=2.395
r94 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.865 $Y=2.68
+ $X2=9.865 $Y2=2.395
r95 23 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.865 $Y=1.935
+ $X2=9.865 $Y2=2.395
r96 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.365 $Y=2.765
+ $X2=9.28 $Y2=2.85
r97 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=2.765
+ $X2=9.865 $Y2=2.68
r98 21 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=2.765
+ $X2=9.365 $Y2=2.765
r99 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.85
+ $X2=9.865 $Y2=1.935
r100 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=1.85
+ $X2=9.365 $Y2=1.85
r101 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=1.765
+ $X2=9.365 $Y2=1.85
r102 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.28 $Y=1.765
+ $X2=9.28 $Y2=0.825
r103 13 36 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=9.925 $Y=4.585
+ $X2=9.925 $Y2=2.56
r104 9 35 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.925 $Y=1.075
+ $X2=9.925 $Y2=2.23
r105 2 41 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=9.155
+ $Y=3.085 $X2=9.28 $Y2=5.835
r106 2 39 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=9.155
+ $Y=3.085 $X2=9.28 $Y2=3.455
r107 1 17 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=9.155
+ $Y=0.575 $X2=9.28 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_300_617# 1 2 9 13 14 17
r20 17 19 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.5 $Y=3.795
+ $X2=2.5 $Y2=5.835
r21 15 17 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.5 $Y=3.715 $X2=2.5
+ $Y2=3.795
r22 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=3.63
+ $X2=2.5 $Y2=3.715
r23 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.415 $Y=3.63
+ $X2=1.725 $Y2=3.63
r24 9 11 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.64 $Y=3.795
+ $X2=1.64 $Y2=5.835
r25 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.715
+ $X2=1.725 $Y2=3.63
r26 7 9 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.64 $Y=3.715 $X2=1.64
+ $Y2=3.795
r27 2 19 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.36
+ $Y=3.085 $X2=2.5 $Y2=5.835
r28 2 17 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=2.36
+ $Y=3.085 $X2=2.5 $Y2=3.795
r29 1 11 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=5.835
r30 1 9 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%A_1469_617# 1 2 9 13 14 17
r19 17 19 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=8.33 $Y=3.795
+ $X2=8.33 $Y2=5.835
r20 15 17 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=8.33 $Y=3.715 $X2=8.33
+ $Y2=3.795
r21 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.245 $Y=3.63
+ $X2=8.33 $Y2=3.715
r22 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.245 $Y=3.63
+ $X2=7.555 $Y2=3.63
r23 9 11 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=7.47 $Y=3.795
+ $X2=7.47 $Y2=5.835
r24 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=3.715
+ $X2=7.555 $Y2=3.63
r25 7 9 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.47 $Y=3.715 $X2=7.47
+ $Y2=3.795
r26 2 19 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=8.19
+ $Y=3.085 $X2=8.33 $Y2=5.835
r27 2 17 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=8.19
+ $Y=3.085 $X2=8.33 $Y2=3.795
r28 1 11 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=7.345
+ $Y=3.085 $X2=7.47 $Y2=5.835
r29 1 9 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=7.345
+ $Y=3.085 $X2=7.47 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__DFFSR_1%Q 1 2 9 12 15 20 23 25
r20 25 30 163.428 $w=1.68e-07 $l=2.505e-06 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.14 $Y2=5.835
r21 23 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.14 $Y=3.33
+ $X2=10.14 $Y2=3.33
r22 18 25 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.14 $Y=3.175
+ $X2=10.14 $Y2=3.33
r23 17 20 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=3.09
+ $X2=10.255 $Y2=3.09
r24 17 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=3.09
+ $X2=10.14 $Y2=3.175
r25 13 15 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=1.515
+ $X2=10.255 $Y2=1.515
r26 12 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=3.005
+ $X2=10.255 $Y2=3.09
r27 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=1.6
+ $X2=10.255 $Y2=1.515
r28 11 12 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=10.255 $Y=1.6
+ $X2=10.255 $Y2=3.005
r29 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=1.43
+ $X2=10.14 $Y2=1.515
r30 7 9 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=10.14 $Y=1.43
+ $X2=10.14 $Y2=0.825
r31 2 30 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=10
+ $Y=3.085 $X2=10.14 $Y2=5.835
r32 2 25 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=10
+ $Y=3.085 $X2=10.14 $Y2=3.455
r33 1 9 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=10 $Y=0.575
+ $X2=10.14 $Y2=0.825
.ends

