* File: sky130_osu_sc_12T_ms__inv_2.pxi.spice
* Created: Fri Nov 12 15:24:10 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__INV_2%GND N_GND_M1000_d N_GND_M1002_d N_GND_M1000_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_MS__INV_2%GND
x_PM_SKY130_OSU_SC_12T_MS__INV_2%VDD N_VDD_M1001_s N_VDD_M1003_s N_VDD_M1001_b
+ N_VDD_c_28_p N_VDD_c_29_p N_VDD_c_35_p VDD N_VDD_c_30_p
+ PM_SKY130_OSU_SC_12T_MS__INV_2%VDD
x_PM_SKY130_OSU_SC_12T_MS__INV_2%A N_A_c_48_n N_A_M1000_g N_A_c_52_n N_A_c_66_n
+ N_A_M1001_g N_A_c_53_n N_A_c_54_n N_A_c_55_n N_A_M1002_g N_A_c_71_n
+ N_A_M1003_g N_A_c_59_n N_A_c_60_n N_A_c_61_n N_A_c_62_n N_A_c_63_n N_A_c_64_n
+ N_A_c_65_n A PM_SKY130_OSU_SC_12T_MS__INV_2%A
x_PM_SKY130_OSU_SC_12T_MS__INV_2%Y N_Y_M1000_s N_Y_M1001_d N_Y_c_115_n
+ N_Y_c_123_n Y N_Y_c_119_n N_Y_c_126_n PM_SKY130_OSU_SC_12T_MS__INV_2%Y
cc_1 N_GND_M1000_b N_A_c_48_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.22
cc_2 N_GND_c_2_p N_A_c_48_n 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=1.22
cc_3 N_GND_c_3_p N_A_c_48_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.22
cc_4 N_GND_c_4_p N_A_c_48_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.22
cc_5 N_GND_M1000_b N_A_c_52_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.33
cc_6 N_GND_M1000_b N_A_c_53_n 0.0349926f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.295
cc_7 N_GND_M1000_b N_A_c_54_n 0.0263741f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.405
cc_8 N_GND_M1000_b N_A_c_55_n 0.0208613f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.22
cc_9 N_GND_c_3_p N_A_c_55_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.22
cc_10 N_GND_c_10_p N_A_c_55_n 0.00502587f $X=1.12 $Y=0.755 $X2=0.905 $Y2=1.22
cc_11 N_GND_c_4_p N_A_c_55_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=1.22
cc_12 N_GND_M1000_b N_A_c_59_n 0.0104975f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.295
cc_13 N_GND_M1000_b N_A_c_60_n 0.0348407f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_14 N_GND_M1000_b N_A_c_61_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.66
cc_15 N_GND_M1000_b N_A_c_62_n 0.00422485f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.405
cc_16 N_GND_M1000_b N_A_c_63_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.85
cc_17 N_GND_M1000_b N_A_c_64_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.825
cc_18 N_GND_M1000_b N_A_c_65_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_19 N_GND_M1000_b N_Y_c_115_n 0.00154299f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.755
cc_20 N_GND_c_3_p N_Y_c_115_n 0.00740081f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.755
cc_21 N_GND_c_4_p N_Y_c_115_n 0.0047139f $X=1.02 $Y=0.19 $X2=0.69 $Y2=0.755
cc_22 N_GND_M1000_b Y 0.0458015f $X=-0.045 $Y=0 $X2=0.76 $Y2=1.72
cc_23 N_GND_M1000_b N_Y_c_119_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1
cc_24 N_GND_c_2_p N_Y_c_119_n 0.00125659f $X=0.26 $Y=0.755 $X2=0.69 $Y2=1
cc_25 N_GND_c_3_p N_Y_c_119_n 0.00245319f $X=1.035 $Y=0.152 $X2=0.69 $Y2=1
cc_26 N_GND_c_10_p N_Y_c_119_n 0.00125659f $X=1.12 $Y=0.755 $X2=0.69 $Y2=1
cc_27 N_VDD_M1001_b N_A_c_66_n 0.0181616f $X=-0.045 $Y=2.425 $X2=0.475 $Y2=2.48
cc_28 N_VDD_c_28_p N_A_c_66_n 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=2.48
cc_29 N_VDD_c_29_p N_A_c_66_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=2.48
cc_30 N_VDD_c_30_p N_A_c_66_n 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=2.48
cc_31 N_VDD_M1001_b N_A_c_54_n 0.00833572f $X=-0.045 $Y=2.425 $X2=0.83 $Y2=2.405
cc_32 N_VDD_M1001_b N_A_c_71_n 0.0207946f $X=-0.045 $Y=2.425 $X2=0.905 $Y2=2.48
cc_33 N_VDD_c_28_p N_A_c_71_n 3.67508e-19 $X=0.26 $Y=3.635 $X2=0.905 $Y2=2.48
cc_34 N_VDD_c_29_p N_A_c_71_n 0.00610567f $X=1.035 $Y=4.287 $X2=0.905 $Y2=2.48
cc_35 N_VDD_c_35_p N_A_c_71_n 0.00656078f $X=1.12 $Y=2.955 $X2=0.905 $Y2=2.48
cc_36 N_VDD_c_30_p N_A_c_71_n 0.00470215f $X=1.02 $Y=4.25 $X2=0.905 $Y2=2.48
cc_37 N_VDD_M1001_b N_A_c_62_n 0.00244597f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.405
cc_38 N_VDD_M1001_s N_A_c_63_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.85
cc_39 N_VDD_M1001_b N_A_c_63_n 0.00618364f $X=-0.045 $Y=2.425 $X2=0.32 $Y2=2.85
cc_40 N_VDD_c_28_p N_A_c_63_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_41 N_VDD_M1001_s A 0.0162774f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.845
cc_42 N_VDD_c_28_p A 0.00522047f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.845
cc_43 N_VDD_c_35_p A 9.09141e-19 $X=1.12 $Y=2.955 $X2=0.32 $Y2=2.845
cc_44 N_VDD_M1001_b N_Y_c_123_n 0.00361433f $X=-0.045 $Y=2.425 $X2=0.69 $Y2=2.48
cc_45 N_VDD_c_29_p N_Y_c_123_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69 $Y2=2.48
cc_46 N_VDD_c_30_p N_Y_c_123_n 0.00475776f $X=1.02 $Y=4.25 $X2=0.69 $Y2=2.48
cc_47 N_VDD_M1001_b N_Y_c_126_n 0.00248543f $X=-0.045 $Y=2.425 $X2=0.69 $Y2=2.48
cc_48 A N_Y_M1001_d 0.00250716f $X=0.32 $Y=2.845 $X2=0.55 $Y2=2.605
cc_49 N_A_c_48_n N_Y_c_115_n 0.00182852f $X=0.475 $Y=1.22 $X2=0.69 $Y2=0.755
cc_50 N_A_c_53_n N_Y_c_115_n 0.00251439f $X=0.83 $Y=1.295 $X2=0.69 $Y2=0.755
cc_51 N_A_c_55_n N_Y_c_115_n 0.00182852f $X=0.905 $Y=1.22 $X2=0.69 $Y2=0.755
cc_52 N_A_c_65_n N_Y_c_115_n 0.00109947f $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.755
cc_53 N_A_c_66_n N_Y_c_123_n 0.00183112f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.48
cc_54 N_A_c_54_n N_Y_c_123_n 0.00839237f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.48
cc_55 N_A_c_71_n N_Y_c_123_n 0.00335296f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.48
cc_56 N_A_c_60_n N_Y_c_123_n 2.38128e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_57 N_A_c_63_n N_Y_c_123_n 0.0226156f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_58 N_A_c_65_n N_Y_c_123_n 0.00165526f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_59 A N_Y_c_123_n 0.00938699f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.48
cc_60 N_A_c_48_n Y 0.00150089f $X=0.475 $Y=1.22 $X2=0.76 $Y2=1.72
cc_61 N_A_c_52_n Y 0.00792324f $X=0.475 $Y=2.33 $X2=0.76 $Y2=1.72
cc_62 N_A_c_53_n Y 0.0155521f $X=0.83 $Y=1.295 $X2=0.76 $Y2=1.72
cc_63 N_A_c_54_n Y 0.00371247f $X=0.83 $Y=2.405 $X2=0.76 $Y2=1.72
cc_64 N_A_c_55_n Y 0.00150089f $X=0.905 $Y=1.22 $X2=0.76 $Y2=1.72
cc_65 N_A_c_60_n Y 0.00610708f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_66 N_A_c_61_n Y 0.00675469f $X=0.535 $Y=1.66 $X2=0.76 $Y2=1.72
cc_67 N_A_c_63_n Y 0.0182346f $X=0.32 $Y=2.85 $X2=0.76 $Y2=1.72
cc_68 N_A_c_65_n Y 0.0178517f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_69 N_A_c_48_n N_Y_c_119_n 0.0084937f $X=0.475 $Y=1.22 $X2=0.69 $Y2=1
cc_70 N_A_c_55_n N_Y_c_119_n 0.0084676f $X=0.905 $Y=1.22 $X2=0.69 $Y2=1
cc_71 N_A_c_60_n N_Y_c_119_n 6.32153e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=1
cc_72 N_A_c_66_n N_Y_c_126_n 0.00166042f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.48
cc_73 N_A_c_54_n N_Y_c_126_n 0.00715376f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.48
cc_74 N_A_c_71_n N_Y_c_126_n 0.00524573f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.48
cc_75 N_A_c_60_n N_Y_c_126_n 2.98633e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_76 N_A_c_62_n N_Y_c_126_n 9.8958e-19 $X=0.475 $Y=2.405 $X2=0.69 $Y2=2.48
cc_77 N_A_c_63_n N_Y_c_126_n 0.00637867f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_78 N_A_c_65_n N_Y_c_126_n 0.00173027f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_79 A N_Y_c_126_n 0.00805971f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.48
