* File: sky130_osu_sc_18T_ls__buf_6.pxi.spice
* Created: Fri Nov 12 14:15:03 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_1 N_noxref_1_M1005_d N_noxref_1_M1001_s
+ N_noxref_1_M1010_s N_noxref_1_M1013_s N_noxref_1_M1005_b N_noxref_1_c_2_p
+ N_noxref_1_c_3_p N_noxref_1_c_9_p N_noxref_1_c_13_p N_noxref_1_c_21_p
+ N_noxref_1_c_26_p N_noxref_1_c_32_p N_noxref_1_c_38_p N_noxref_1_c_85_p
+ N_noxref_1_c_86_p PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_1
x_PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_2 N_noxref_2_M1004_d N_noxref_2_M1003_s
+ N_noxref_2_M1007_s N_noxref_2_M1012_s N_noxref_2_M1004_b N_noxref_2_c_88_p
+ N_noxref_2_c_89_p N_noxref_2_c_97_p N_noxref_2_c_101_p N_noxref_2_c_107_p
+ N_noxref_2_c_111_p N_noxref_2_c_116_p N_noxref_2_c_120_p N_noxref_2_c_144_p
+ N_noxref_2_c_145_p N_noxref_2_c_146_p PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_2
x_PM_SKY130_OSU_SC_18T_LS__BUF_6%A N_A_M1005_g N_A_M1004_g N_A_c_151_n
+ N_A_c_152_n A PM_SKY130_OSU_SC_18T_LS__BUF_6%A
x_PM_SKY130_OSU_SC_18T_LS__BUF_6%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1004_s N_A_27_115#_M1000_g N_A_27_115#_c_232_n
+ N_A_27_115#_M1002_g N_A_27_115#_c_190_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_235_n N_A_27_115#_M1003_g N_A_27_115#_c_194_n
+ N_A_27_115#_c_196_n N_A_27_115#_c_197_n N_A_27_115#_c_198_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_242_n N_A_27_115#_M1006_g
+ N_A_27_115#_c_202_n N_A_27_115#_c_203_n N_A_27_115#_M1010_g
+ N_A_27_115#_c_246_n N_A_27_115#_M1007_g N_A_27_115#_c_207_n
+ N_A_27_115#_c_209_n N_A_27_115#_M1011_g N_A_27_115#_c_213_n
+ N_A_27_115#_c_251_n N_A_27_115#_M1009_g N_A_27_115#_c_214_n
+ N_A_27_115#_c_215_n N_A_27_115#_M1013_g N_A_27_115#_c_255_n
+ N_A_27_115#_M1012_g N_A_27_115#_c_219_n N_A_27_115#_c_220_n
+ N_A_27_115#_c_221_n N_A_27_115#_c_222_n N_A_27_115#_c_223_n
+ N_A_27_115#_c_224_n N_A_27_115#_c_225_n N_A_27_115#_c_227_n
+ N_A_27_115#_c_228_n N_A_27_115#_c_230_n N_A_27_115#_c_231_n
+ PM_SKY130_OSU_SC_18T_LS__BUF_6%A_27_115#
x_PM_SKY130_OSU_SC_18T_LS__BUF_6%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1011_d
+ N_Y_M1002_d N_Y_M1006_d N_Y_M1009_d N_Y_c_364_n N_Y_c_392_n N_Y_c_367_n
+ N_Y_c_394_n N_Y_c_371_n N_Y_c_396_n N_Y_c_374_n N_Y_c_377_n Y N_Y_c_379_n
+ N_Y_c_399_n N_Y_c_381_n N_Y_c_382_n N_Y_c_384_n N_Y_c_401_n N_Y_c_387_n
+ N_Y_c_388_n N_Y_c_391_n PM_SKY130_OSU_SC_18T_LS__BUF_6%Y
cc_1 N_noxref_1_M1005_b N_A_M1005_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=1.075
cc_2 N_noxref_1_c_2_p N_A_M1005_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475
+ $Y2=1.075
cc_3 N_noxref_1_c_3_p N_A_M1005_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475
+ $Y2=1.075
cc_4 N_noxref_1_M1005_b N_A_M1004_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=4.585
cc_5 N_noxref_1_M1005_b N_A_c_151_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_6 N_noxref_1_M1005_b N_A_c_152_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635
+ $Y2=2.48
cc_7 N_noxref_1_M1005_b N_A_27_115#_M1000_g 0.0207501f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=1.075
cc_8 N_noxref_1_c_3_p N_A_27_115#_M1000_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=1.075
cc_9 N_noxref_1_c_9_p N_A_27_115#_M1000_g 0.00606474f $X=1.465 $Y=0.152
+ $X2=0.905 $Y2=1.075
cc_10 N_noxref_1_M1005_b N_A_27_115#_c_190_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.86
cc_11 N_noxref_1_M1005_b N_A_27_115#_M1001_g 0.020212f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_12 N_noxref_1_c_9_p N_A_27_115#_M1001_g 0.00606474f $X=1.465 $Y=0.152
+ $X2=1.335 $Y2=1.075
cc_13 N_noxref_1_c_13_p N_A_27_115#_M1001_g 0.00356864f $X=1.55 $Y=0.825
+ $X2=1.335 $Y2=1.075
cc_14 N_noxref_1_M1005_b N_A_27_115#_c_194_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.845
cc_15 N_noxref_1_c_13_p N_A_27_115#_c_194_n 0.00256938f $X=1.55 $Y=0.825
+ $X2=1.69 $Y2=1.845
cc_16 N_noxref_1_M1005_b N_A_27_115#_c_196_n 0.0429274f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.845
cc_17 N_noxref_1_M1005_b N_A_27_115#_c_197_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.935
cc_18 N_noxref_1_M1005_b N_A_27_115#_c_198_n 0.0196789f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.935
cc_19 N_noxref_1_M1005_b N_A_27_115#_M1008_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_20 N_noxref_1_c_13_p N_A_27_115#_M1008_g 0.00356864f $X=1.55 $Y=0.825
+ $X2=1.765 $Y2=1.075
cc_21 N_noxref_1_c_21_p N_A_27_115#_M1008_g 0.00606474f $X=2.325 $Y=0.152
+ $X2=1.765 $Y2=1.075
cc_22 N_noxref_1_M1005_b N_A_27_115#_c_202_n 0.0195339f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.845
cc_23 N_noxref_1_M1005_b N_A_27_115#_c_203_n 0.0107618f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.935
cc_24 N_noxref_1_M1005_b N_A_27_115#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.075
cc_25 N_noxref_1_c_21_p N_A_27_115#_M1010_g 0.00606474f $X=2.325 $Y=0.152
+ $X2=2.195 $Y2=1.075
cc_26 N_noxref_1_c_26_p N_A_27_115#_M1010_g 0.00356864f $X=2.41 $Y=0.825
+ $X2=2.195 $Y2=1.075
cc_27 N_noxref_1_M1005_b N_A_27_115#_c_207_n 0.0165886f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.845
cc_28 N_noxref_1_c_26_p N_A_27_115#_c_207_n 0.00256938f $X=2.41 $Y=0.825
+ $X2=2.55 $Y2=1.845
cc_29 N_noxref_1_M1005_b N_A_27_115#_c_209_n 0.0109555f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.935
cc_30 N_noxref_1_M1005_b N_A_27_115#_M1011_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.075
cc_31 N_noxref_1_c_26_p N_A_27_115#_M1011_g 0.00356864f $X=2.41 $Y=0.825
+ $X2=2.625 $Y2=1.075
cc_32 N_noxref_1_c_32_p N_A_27_115#_M1011_g 0.00606474f $X=3.185 $Y=0.152
+ $X2=2.625 $Y2=1.075
cc_33 N_noxref_1_M1005_b N_A_27_115#_c_213_n 0.0668243f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.86
cc_34 N_noxref_1_M1005_b N_A_27_115#_c_214_n 0.0385034f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.845
cc_35 N_noxref_1_M1005_b N_A_27_115#_c_215_n 0.0221499f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.935
cc_36 N_noxref_1_M1005_b N_A_27_115#_M1013_g 0.0264941f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.075
cc_37 N_noxref_1_c_32_p N_A_27_115#_M1013_g 0.00606474f $X=3.185 $Y=0.152
+ $X2=3.055 $Y2=1.075
cc_38 N_noxref_1_c_38_p N_A_27_115#_M1013_g 0.00713292f $X=3.27 $Y=0.825
+ $X2=3.055 $Y2=1.075
cc_39 N_noxref_1_M1005_b N_A_27_115#_c_219_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.845
cc_40 N_noxref_1_M1005_b N_A_27_115#_c_220_n 0.00890086f $X=-0.045 $Y=0
+ $X2=1.765 $Y2=2.935
cc_41 N_noxref_1_M1005_b N_A_27_115#_c_221_n 0.0106787f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.845
cc_42 N_noxref_1_M1005_b N_A_27_115#_c_222_n 0.00890086f $X=-0.045 $Y=0
+ $X2=2.195 $Y2=2.935
cc_43 N_noxref_1_M1005_b N_A_27_115#_c_223_n 0.0023879f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.845
cc_44 N_noxref_1_M1005_b N_A_27_115#_c_224_n 7.16371e-19 $X=-0.045 $Y=0
+ $X2=2.625 $Y2=2.935
cc_45 N_noxref_1_M1005_b N_A_27_115#_c_225_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_46 N_noxref_1_c_2_p N_A_27_115#_c_225_n 0.00736239f $X=0.605 $Y=0.152
+ $X2=0.26 $Y2=0.825
cc_47 N_noxref_1_M1005_b N_A_27_115#_c_227_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.455
cc_48 N_noxref_1_M1005_b N_A_27_115#_c_228_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.935
cc_49 N_noxref_1_c_3_p N_A_27_115#_c_228_n 0.00702738f $X=0.69 $Y=0.825 $X2=0.88
+ $Y2=1.935
cc_50 N_noxref_1_M1005_b N_A_27_115#_c_230_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.935
cc_51 N_noxref_1_M1005_b N_A_27_115#_c_231_n 0.00592383f $X=-0.045 $Y=0
+ $X2=0.965 $Y2=1.935
cc_52 N_noxref_1_M1005_b N_Y_c_364_n 0.00155118f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.825
cc_53 N_noxref_1_c_9_p N_Y_c_364_n 0.00734006f $X=1.465 $Y=0.152 $X2=1.12
+ $Y2=0.825
cc_54 N_noxref_1_c_13_p N_Y_c_364_n 8.14297e-19 $X=1.55 $Y=0.825 $X2=1.12
+ $Y2=0.825
cc_55 N_noxref_1_M1005_b N_Y_c_367_n 0.00155118f $X=-0.045 $Y=0 $X2=1.98
+ $Y2=0.825
cc_56 N_noxref_1_c_13_p N_Y_c_367_n 8.14297e-19 $X=1.55 $Y=0.825 $X2=1.98
+ $Y2=0.825
cc_57 N_noxref_1_c_21_p N_Y_c_367_n 0.00754406f $X=2.325 $Y=0.152 $X2=1.98
+ $Y2=0.825
cc_58 N_noxref_1_c_26_p N_Y_c_367_n 8.14297e-19 $X=2.41 $Y=0.825 $X2=1.98
+ $Y2=0.825
cc_59 N_noxref_1_M1005_b N_Y_c_371_n 0.00155118f $X=-0.045 $Y=0 $X2=2.84
+ $Y2=0.825
cc_60 N_noxref_1_c_26_p N_Y_c_371_n 8.14297e-19 $X=2.41 $Y=0.825 $X2=2.84
+ $Y2=0.825
cc_61 N_noxref_1_c_32_p N_Y_c_371_n 0.00746708f $X=3.185 $Y=0.152 $X2=2.84
+ $Y2=0.825
cc_62 N_noxref_1_M1005_b N_Y_c_374_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=1.595
cc_63 N_noxref_1_c_3_p N_Y_c_374_n 0.00134236f $X=0.69 $Y=0.825 $X2=1.12
+ $Y2=1.595
cc_64 N_noxref_1_c_13_p N_Y_c_374_n 7.53951e-19 $X=1.55 $Y=0.825 $X2=1.12
+ $Y2=1.595
cc_65 N_noxref_1_M1005_b N_Y_c_377_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=2.845
cc_66 N_noxref_1_M1005_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=2.27
cc_67 N_noxref_1_M1001_s N_Y_c_379_n 0.0127884f $X=1.41 $Y=0.575 $X2=1.835
+ $Y2=1.48
cc_68 N_noxref_1_c_13_p N_Y_c_379_n 0.0142303f $X=1.55 $Y=0.825 $X2=1.835
+ $Y2=1.48
cc_69 N_noxref_1_M1005_b N_Y_c_381_n 0.0437239f $X=-0.045 $Y=0 $X2=1.98
+ $Y2=2.845
cc_70 N_noxref_1_M1010_s N_Y_c_382_n 0.0127884f $X=2.27 $Y=0.575 $X2=2.695
+ $Y2=1.48
cc_71 N_noxref_1_c_26_p N_Y_c_382_n 0.0142303f $X=2.41 $Y=0.825 $X2=2.695
+ $Y2=1.48
cc_72 N_noxref_1_M1005_b N_Y_c_384_n 0.00409378f $X=-0.045 $Y=0 $X2=2.125
+ $Y2=1.48
cc_73 N_noxref_1_c_13_p N_Y_c_384_n 7.53951e-19 $X=1.55 $Y=0.825 $X2=2.125
+ $Y2=1.48
cc_74 N_noxref_1_c_26_p N_Y_c_384_n 7.53951e-19 $X=2.41 $Y=0.825 $X2=2.125
+ $Y2=1.48
cc_75 N_noxref_1_M1005_b N_Y_c_387_n 0.00560779f $X=-0.045 $Y=0 $X2=2.125
+ $Y2=2.96
cc_76 N_noxref_1_M1005_b N_Y_c_388_n 0.00409378f $X=-0.045 $Y=0 $X2=2.84
+ $Y2=1.595
cc_77 N_noxref_1_c_26_p N_Y_c_388_n 7.53951e-19 $X=2.41 $Y=0.825 $X2=2.84
+ $Y2=1.595
cc_78 N_noxref_1_c_38_p N_Y_c_388_n 0.00134236f $X=3.27 $Y=0.825 $X2=2.84
+ $Y2=1.595
cc_79 N_noxref_1_M1005_b N_Y_c_391_n 0.0625307f $X=-0.045 $Y=0 $X2=2.84
+ $Y2=2.845
cc_80 N_noxref_1_M1005_b GND 0.251858f $X=-0.045 $Y=0 $X2=0.34 $Y2=0.22
cc_81 N_noxref_1_c_2_p GND 0.0440059f $X=0.605 $Y=0.152 $X2=0.34 $Y2=0.22
cc_82 N_noxref_1_c_9_p GND 0.0435303f $X=1.465 $Y=0.152 $X2=0.34 $Y2=0.22
cc_83 N_noxref_1_c_21_p GND 0.042979f $X=2.325 $Y=0.152 $X2=0.34 $Y2=0.22
cc_84 N_noxref_1_c_32_p GND 0.0887744f $X=3.185 $Y=0.152 $X2=0.34 $Y2=0.22
cc_85 N_noxref_1_c_85_p GND 0.0189324f $X=0.69 $Y=0.152 $X2=0.34 $Y2=0.22
cc_86 N_noxref_1_c_86_p GND 0.0189324f $X=1.55 $Y=0.152 $X2=0.34 $Y2=0.22
cc_87 N_noxref_2_M1004_b N_A_M1004_g 0.0245629f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_88 N_noxref_2_c_88_p N_A_M1004_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_89 N_noxref_2_c_89_p N_A_M1004_g 0.00354579f $X=0.69 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_90 N_noxref_2_M1004_d N_A_c_152_n 0.00628533f $X=0.55 $Y=3.085 $X2=0.635
+ $Y2=2.48
cc_91 N_noxref_2_M1004_b N_A_c_152_n 0.00328912f $X=-0.045 $Y=2.905 $X2=0.635
+ $Y2=2.48
cc_92 N_noxref_2_c_89_p N_A_c_152_n 0.00264661f $X=0.69 $Y=4.135 $X2=0.635
+ $Y2=2.48
cc_93 N_noxref_2_M1004_d A 0.00797576f $X=0.55 $Y=3.085 $X2=0.635 $Y2=3.33
cc_94 N_noxref_2_c_89_p A 0.00510982f $X=0.69 $Y=4.135 $X2=0.635 $Y2=3.33
cc_95 N_noxref_2_M1004_b N_A_27_115#_c_232_n 0.014249f $X=-0.045 $Y=2.905
+ $X2=0.905 $Y2=3.01
cc_96 N_noxref_2_c_89_p N_A_27_115#_c_232_n 0.00354579f $X=0.69 $Y=4.135
+ $X2=0.905 $Y2=3.01
cc_97 N_noxref_2_c_97_p N_A_27_115#_c_232_n 0.00606474f $X=1.465 $Y=6.507
+ $X2=0.905 $Y2=3.01
cc_98 N_noxref_2_M1004_b N_A_27_115#_c_235_n 0.0141063f $X=-0.045 $Y=2.905
+ $X2=1.335 $Y2=3.01
cc_99 N_noxref_2_c_89_p N_A_27_115#_c_235_n 3.67508e-19 $X=0.69 $Y=4.135
+ $X2=1.335 $Y2=3.01
cc_100 N_noxref_2_c_97_p N_A_27_115#_c_235_n 0.00610567f $X=1.465 $Y=6.507
+ $X2=1.335 $Y2=3.01
cc_101 N_noxref_2_c_101_p N_A_27_115#_c_235_n 0.00373985f $X=1.55 $Y=3.455
+ $X2=1.335 $Y2=3.01
cc_102 N_noxref_2_M1004_b N_A_27_115#_c_197_n 0.00647677f $X=-0.045 $Y=2.905
+ $X2=1.69 $Y2=2.935
cc_103 N_noxref_2_c_101_p N_A_27_115#_c_197_n 0.00364479f $X=1.55 $Y=3.455
+ $X2=1.69 $Y2=2.935
cc_104 N_noxref_2_M1004_b N_A_27_115#_c_198_n 0.0113915f $X=-0.045 $Y=2.905
+ $X2=1.41 $Y2=2.935
cc_105 N_noxref_2_M1004_b N_A_27_115#_c_242_n 0.0137901f $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=3.01
cc_106 N_noxref_2_c_101_p N_A_27_115#_c_242_n 0.00354579f $X=1.55 $Y=3.455
+ $X2=1.765 $Y2=3.01
cc_107 N_noxref_2_c_107_p N_A_27_115#_c_242_n 0.00606474f $X=2.325 $Y=6.507
+ $X2=1.765 $Y2=3.01
cc_108 N_noxref_2_M1004_b N_A_27_115#_c_203_n 0.00596183f $X=-0.045 $Y=2.905
+ $X2=2.12 $Y2=2.935
cc_109 N_noxref_2_M1004_b N_A_27_115#_c_246_n 0.0137901f $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=3.01
cc_110 N_noxref_2_c_107_p N_A_27_115#_c_246_n 0.00606474f $X=2.325 $Y=6.507
+ $X2=2.195 $Y2=3.01
cc_111 N_noxref_2_c_111_p N_A_27_115#_c_246_n 0.00354579f $X=2.41 $Y=3.455
+ $X2=2.195 $Y2=3.01
cc_112 N_noxref_2_M1004_b N_A_27_115#_c_209_n 0.00647677f $X=-0.045 $Y=2.905
+ $X2=2.55 $Y2=2.935
cc_113 N_noxref_2_c_111_p N_A_27_115#_c_209_n 0.00364479f $X=2.41 $Y=3.455
+ $X2=2.55 $Y2=2.935
cc_114 N_noxref_2_M1004_b N_A_27_115#_c_251_n 0.0137901f $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=3.01
cc_115 N_noxref_2_c_111_p N_A_27_115#_c_251_n 0.00354579f $X=2.41 $Y=3.455
+ $X2=2.625 $Y2=3.01
cc_116 N_noxref_2_c_116_p N_A_27_115#_c_251_n 0.00606474f $X=3.185 $Y=6.507
+ $X2=2.625 $Y2=3.01
cc_117 N_noxref_2_M1004_b N_A_27_115#_c_215_n 0.0134369f $X=-0.045 $Y=2.905
+ $X2=2.98 $Y2=2.935
cc_118 N_noxref_2_M1004_b N_A_27_115#_c_255_n 0.0166569f $X=-0.045 $Y=2.905
+ $X2=3.055 $Y2=3.01
cc_119 N_noxref_2_c_116_p N_A_27_115#_c_255_n 0.00606474f $X=3.185 $Y=6.507
+ $X2=3.055 $Y2=3.01
cc_120 N_noxref_2_c_120_p N_A_27_115#_c_255_n 0.00713292f $X=3.27 $Y=3.455
+ $X2=3.055 $Y2=3.01
cc_121 N_noxref_2_M1004_b N_A_27_115#_c_220_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.935
cc_122 N_noxref_2_M1004_b N_A_27_115#_c_222_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.935
cc_123 N_noxref_2_M1004_b N_A_27_115#_c_224_n 0.00167153f $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=2.935
cc_124 N_noxref_2_M1004_b N_A_27_115#_c_227_n 0.00996008f $X=-0.045 $Y=2.905
+ $X2=0.26 $Y2=3.455
cc_125 N_noxref_2_c_88_p N_A_27_115#_c_227_n 0.00736239f $X=0.605 $Y=6.507
+ $X2=0.26 $Y2=3.455
cc_126 N_noxref_2_M1004_b N_Y_c_392_n 0.00290209f $X=-0.045 $Y=2.905 $X2=1.12
+ $Y2=2.96
cc_127 N_noxref_2_c_97_p N_Y_c_392_n 0.00734006f $X=1.465 $Y=6.507 $X2=1.12
+ $Y2=2.96
cc_128 N_noxref_2_M1004_b N_Y_c_394_n 0.00337919f $X=-0.045 $Y=2.905 $X2=1.98
+ $Y2=2.96
cc_129 N_noxref_2_c_107_p N_Y_c_394_n 0.00754406f $X=2.325 $Y=6.507 $X2=1.98
+ $Y2=2.96
cc_130 N_noxref_2_M1004_b N_Y_c_396_n 0.00337919f $X=-0.045 $Y=2.905 $X2=2.84
+ $Y2=2.96
cc_131 N_noxref_2_c_116_p N_Y_c_396_n 0.00746708f $X=3.185 $Y=6.507 $X2=2.84
+ $Y2=2.96
cc_132 N_noxref_2_M1004_b N_Y_c_377_n 0.00409378f $X=-0.045 $Y=2.905 $X2=1.12
+ $Y2=2.845
cc_133 N_noxref_2_M1004_b N_Y_c_399_n 0.00520877f $X=-0.045 $Y=2.905 $X2=1.835
+ $Y2=2.96
cc_134 N_noxref_2_c_101_p N_Y_c_399_n 0.0090257f $X=1.55 $Y=3.455 $X2=1.835
+ $Y2=2.96
cc_135 N_noxref_2_M1004_b N_Y_c_401_n 0.00520877f $X=-0.045 $Y=2.905 $X2=2.695
+ $Y2=2.96
cc_136 N_noxref_2_c_111_p N_Y_c_401_n 0.0090257f $X=2.41 $Y=3.455 $X2=2.695
+ $Y2=2.96
cc_137 N_noxref_2_M1004_b N_Y_c_387_n 0.00409378f $X=-0.045 $Y=2.905 $X2=2.125
+ $Y2=2.96
cc_138 N_noxref_2_M1004_b N_Y_c_391_n 0.00409378f $X=-0.045 $Y=2.905 $X2=2.84
+ $Y2=2.845
cc_139 N_noxref_2_M1004_b VDD 0.269451f $X=-0.045 $Y=2.905 $X2=0.34 $Y2=6.44
cc_140 N_noxref_2_c_88_p VDD 0.0439891f $X=0.605 $Y=6.507 $X2=0.34 $Y2=6.44
cc_141 N_noxref_2_c_97_p VDD 0.0435303f $X=1.465 $Y=6.507 $X2=0.34 $Y2=6.44
cc_142 N_noxref_2_c_107_p VDD 0.042979f $X=2.325 $Y=6.507 $X2=0.34 $Y2=6.44
cc_143 N_noxref_2_c_116_p VDD 0.0887744f $X=3.185 $Y=6.507 $X2=0.34 $Y2=6.44
cc_144 N_noxref_2_c_144_p VDD 0.0189324f $X=0.69 $Y=6.507 $X2=0.34 $Y2=6.44
cc_145 N_noxref_2_c_145_p VDD 0.0189324f $X=1.55 $Y=6.507 $X2=0.34 $Y2=6.44
cc_146 N_noxref_2_c_146_p VDD 0.0189324f $X=2.38 $Y=6.44 $X2=0.34 $Y2=6.44
cc_147 A N_A_27_115#_M1004_s 0.00414531f $X=0.635 $Y=3.33 $X2=0.135 $Y2=3.085
cc_148 N_A_M1005_g N_A_27_115#_M1000_g 0.0387262f $X=0.475 $Y=1.075 $X2=0.905
+ $Y2=1.075
cc_149 A N_A_27_115#_c_232_n 0.00419145f $X=0.635 $Y=3.33 $X2=0.905 $Y2=3.01
cc_150 N_A_M1005_g N_A_27_115#_c_190_n 0.00260138f $X=0.475 $Y=1.075 $X2=1.18
+ $Y2=2.86
cc_151 N_A_M1004_g N_A_27_115#_c_190_n 0.00209773f $X=0.475 $Y=4.585 $X2=1.18
+ $Y2=2.86
cc_152 N_A_c_151_n N_A_27_115#_c_190_n 0.0139096f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_153 N_A_c_152_n N_A_27_115#_c_190_n 0.00361737f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_154 N_A_M1004_g N_A_27_115#_c_198_n 0.0499373f $X=0.475 $Y=4.585 $X2=1.41
+ $Y2=2.935
cc_155 N_A_c_152_n N_A_27_115#_c_198_n 0.00477416f $X=0.635 $Y=2.48 $X2=1.41
+ $Y2=2.935
cc_156 N_A_M1005_g N_A_27_115#_c_225_n 0.0148408f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_157 N_A_M1005_g N_A_27_115#_c_227_n 0.0337582f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=3.455
cc_158 N_A_c_152_n N_A_27_115#_c_227_n 0.0548951f $X=0.635 $Y=2.48 $X2=0.26
+ $Y2=3.455
cc_159 A N_A_27_115#_c_227_n 0.0155137f $X=0.635 $Y=3.33 $X2=0.26 $Y2=3.455
cc_160 N_A_M1005_g N_A_27_115#_c_228_n 0.0207696f $X=0.475 $Y=1.075 $X2=0.88
+ $Y2=1.935
cc_161 N_A_c_151_n N_A_27_115#_c_228_n 0.00273049f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_162 N_A_c_152_n N_A_27_115#_c_228_n 0.00886797f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_163 N_A_M1005_g N_A_27_115#_c_231_n 6.59135e-19 $X=0.475 $Y=1.075 $X2=0.965
+ $Y2=1.935
cc_164 N_A_c_152_n N_Y_c_392_n 0.0135622f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_165 A N_Y_c_392_n 0.00731851f $X=0.635 $Y=3.33 $X2=1.12 $Y2=2.96
cc_166 N_A_M1005_g N_Y_c_374_n 8.23842e-19 $X=0.475 $Y=1.075 $X2=1.12 $Y2=1.595
cc_167 N_A_c_152_n N_Y_c_377_n 0.00677552f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.845
cc_168 N_A_M1005_g Y 0.00310306f $X=0.475 $Y=1.075 $X2=1.055 $Y2=2.27
cc_169 N_A_c_151_n Y 0.00441844f $X=0.635 $Y=2.48 $X2=1.055 $Y2=2.27
cc_170 N_A_c_152_n Y 0.0200396f $X=0.635 $Y=2.48 $X2=1.055 $Y2=2.27
cc_171 N_A_M1005_g GND 0.00468827f $X=0.475 $Y=1.075 $X2=0.34 $Y2=0.22
cc_172 N_A_M1004_g VDD 0.00468827f $X=0.475 $Y=4.585 $X2=0.34 $Y2=6.44
cc_173 N_A_27_115#_M1000_g N_Y_c_364_n 0.00231637f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_174 N_A_27_115#_M1001_g N_Y_c_364_n 0.00231637f $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=0.825
cc_175 N_A_27_115#_c_196_n N_Y_c_364_n 0.0030245f $X=1.41 $Y=1.845 $X2=1.12
+ $Y2=0.825
cc_176 N_A_27_115#_c_231_n N_Y_c_364_n 7.32051e-19 $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_177 N_A_27_115#_c_232_n N_Y_c_392_n 0.00155107f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_178 N_A_27_115#_c_235_n N_Y_c_392_n 0.00250481f $X=1.335 $Y=3.01 $X2=1.12
+ $Y2=2.96
cc_179 N_A_27_115#_c_198_n N_Y_c_392_n 0.0126676f $X=1.41 $Y=2.935 $X2=1.12
+ $Y2=2.96
cc_180 N_A_27_115#_M1008_g N_Y_c_367_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.98
+ $Y2=0.825
cc_181 N_A_27_115#_c_202_n N_Y_c_367_n 0.00280419f $X=2.12 $Y=1.845 $X2=1.98
+ $Y2=0.825
cc_182 N_A_27_115#_M1010_g N_Y_c_367_n 0.00231637f $X=2.195 $Y=1.075 $X2=1.98
+ $Y2=0.825
cc_183 N_A_27_115#_c_242_n N_Y_c_394_n 0.00250481f $X=1.765 $Y=3.01 $X2=1.98
+ $Y2=2.96
cc_184 N_A_27_115#_c_203_n N_Y_c_394_n 0.0138847f $X=2.12 $Y=2.935 $X2=1.98
+ $Y2=2.96
cc_185 N_A_27_115#_c_246_n N_Y_c_394_n 0.00250481f $X=2.195 $Y=3.01 $X2=1.98
+ $Y2=2.96
cc_186 N_A_27_115#_M1011_g N_Y_c_371_n 0.00231637f $X=2.625 $Y=1.075 $X2=2.84
+ $Y2=0.825
cc_187 N_A_27_115#_c_214_n N_Y_c_371_n 0.00280419f $X=2.98 $Y=1.845 $X2=2.84
+ $Y2=0.825
cc_188 N_A_27_115#_M1013_g N_Y_c_371_n 0.00231637f $X=3.055 $Y=1.075 $X2=2.84
+ $Y2=0.825
cc_189 N_A_27_115#_c_251_n N_Y_c_396_n 0.00250481f $X=2.625 $Y=3.01 $X2=2.84
+ $Y2=2.96
cc_190 N_A_27_115#_c_215_n N_Y_c_396_n 0.013404f $X=2.98 $Y=2.935 $X2=2.84
+ $Y2=2.96
cc_191 N_A_27_115#_c_255_n N_Y_c_396_n 0.00250481f $X=3.055 $Y=3.01 $X2=2.84
+ $Y2=2.96
cc_192 N_A_27_115#_M1000_g N_Y_c_374_n 0.00541983f $X=0.905 $Y=1.075 $X2=1.12
+ $Y2=1.595
cc_193 N_A_27_115#_M1001_g N_Y_c_374_n 0.00262362f $X=1.335 $Y=1.075 $X2=1.12
+ $Y2=1.595
cc_194 N_A_27_115#_c_231_n N_Y_c_374_n 0.00278861f $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=1.595
cc_195 N_A_27_115#_c_232_n N_Y_c_377_n 0.00120715f $X=0.905 $Y=3.01 $X2=1.12
+ $Y2=2.845
cc_196 N_A_27_115#_c_190_n N_Y_c_377_n 0.00215118f $X=1.18 $Y=2.86 $X2=1.12
+ $Y2=2.845
cc_197 N_A_27_115#_c_235_n N_Y_c_377_n 0.00113627f $X=1.335 $Y=3.01 $X2=1.12
+ $Y2=2.845
cc_198 N_A_27_115#_c_198_n N_Y_c_377_n 0.00372325f $X=1.41 $Y=2.935 $X2=1.12
+ $Y2=2.845
cc_199 N_A_27_115#_M1000_g Y 0.00251111f $X=0.905 $Y=1.075 $X2=1.055 $Y2=2.27
cc_200 N_A_27_115#_c_190_n Y 0.0314621f $X=1.18 $Y=2.86 $X2=1.055 $Y2=2.27
cc_201 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.055 $Y2=2.27
cc_202 N_A_27_115#_c_196_n Y 0.0166018f $X=1.41 $Y=1.845 $X2=1.055 $Y2=2.27
cc_203 N_A_27_115#_c_228_n Y 8.73078e-19 $X=0.88 $Y=1.935 $X2=1.055 $Y2=2.27
cc_204 N_A_27_115#_c_231_n Y 0.0121742f $X=0.965 $Y=1.935 $X2=1.055 $Y2=2.27
cc_205 N_A_27_115#_M1001_g N_Y_c_379_n 0.0133661f $X=1.335 $Y=1.075 $X2=1.835
+ $Y2=1.48
cc_206 N_A_27_115#_c_194_n N_Y_c_379_n 0.00213861f $X=1.69 $Y=1.845 $X2=1.835
+ $Y2=1.48
cc_207 N_A_27_115#_M1008_g N_Y_c_379_n 0.0130095f $X=1.765 $Y=1.075 $X2=1.835
+ $Y2=1.48
cc_208 N_A_27_115#_c_235_n N_Y_c_399_n 0.00639369f $X=1.335 $Y=3.01 $X2=1.835
+ $Y2=2.96
cc_209 N_A_27_115#_c_197_n N_Y_c_399_n 0.0125005f $X=1.69 $Y=2.935 $X2=1.835
+ $Y2=2.96
cc_210 N_A_27_115#_c_198_n N_Y_c_399_n 0.00627763f $X=1.41 $Y=2.935 $X2=1.835
+ $Y2=2.96
cc_211 N_A_27_115#_c_242_n N_Y_c_399_n 0.00639369f $X=1.765 $Y=3.01 $X2=1.835
+ $Y2=2.96
cc_212 N_A_27_115#_c_220_n N_Y_c_399_n 0.00580646f $X=1.765 $Y=2.935 $X2=1.835
+ $Y2=2.96
cc_213 N_A_27_115#_c_196_n N_Y_c_381_n 0.013329f $X=1.41 $Y=1.845 $X2=1.98
+ $Y2=2.845
cc_214 N_A_27_115#_M1008_g N_Y_c_381_n 0.00251111f $X=1.765 $Y=1.075 $X2=1.98
+ $Y2=2.845
cc_215 N_A_27_115#_c_202_n N_Y_c_381_n 0.0178059f $X=2.12 $Y=1.845 $X2=1.98
+ $Y2=2.845
cc_216 N_A_27_115#_M1010_g N_Y_c_381_n 0.00251111f $X=2.195 $Y=1.075 $X2=1.98
+ $Y2=2.845
cc_217 N_A_27_115#_c_213_n N_Y_c_381_n 0.0137936f $X=2.625 $Y=2.86 $X2=1.98
+ $Y2=2.845
cc_218 N_A_27_115#_M1010_g N_Y_c_382_n 0.0130095f $X=2.195 $Y=1.075 $X2=2.695
+ $Y2=1.48
cc_219 N_A_27_115#_c_207_n N_Y_c_382_n 0.00213861f $X=2.55 $Y=1.845 $X2=2.695
+ $Y2=1.48
cc_220 N_A_27_115#_M1011_g N_Y_c_382_n 0.0136594f $X=2.625 $Y=1.075 $X2=2.695
+ $Y2=1.48
cc_221 N_A_27_115#_M1008_g N_Y_c_384_n 0.00259902f $X=1.765 $Y=1.075 $X2=2.125
+ $Y2=1.48
cc_222 N_A_27_115#_M1010_g N_Y_c_384_n 0.00259902f $X=2.195 $Y=1.075 $X2=2.125
+ $Y2=1.48
cc_223 N_A_27_115#_c_246_n N_Y_c_401_n 0.00639369f $X=2.195 $Y=3.01 $X2=2.695
+ $Y2=2.96
cc_224 N_A_27_115#_c_209_n N_Y_c_401_n 0.0130313f $X=2.55 $Y=2.935 $X2=2.695
+ $Y2=2.96
cc_225 N_A_27_115#_c_251_n N_Y_c_401_n 0.00639369f $X=2.625 $Y=3.01 $X2=2.695
+ $Y2=2.96
cc_226 N_A_27_115#_c_222_n N_Y_c_401_n 0.00580646f $X=2.195 $Y=2.935 $X2=2.695
+ $Y2=2.96
cc_227 N_A_27_115#_c_224_n N_Y_c_401_n 0.00666531f $X=2.625 $Y=2.935 $X2=2.695
+ $Y2=2.96
cc_228 N_A_27_115#_c_242_n N_Y_c_387_n 0.00113627f $X=1.765 $Y=3.01 $X2=2.125
+ $Y2=2.96
cc_229 N_A_27_115#_c_203_n N_Y_c_387_n 0.00364679f $X=2.12 $Y=2.935 $X2=2.125
+ $Y2=2.96
cc_230 N_A_27_115#_c_246_n N_Y_c_387_n 0.00113627f $X=2.195 $Y=3.01 $X2=2.125
+ $Y2=2.96
cc_231 N_A_27_115#_c_220_n N_Y_c_387_n 6.99501e-19 $X=1.765 $Y=2.935 $X2=2.125
+ $Y2=2.96
cc_232 N_A_27_115#_c_222_n N_Y_c_387_n 6.99501e-19 $X=2.195 $Y=2.935 $X2=2.125
+ $Y2=2.96
cc_233 N_A_27_115#_M1011_g N_Y_c_388_n 0.00262362f $X=2.625 $Y=1.075 $X2=2.84
+ $Y2=1.595
cc_234 N_A_27_115#_M1013_g N_Y_c_388_n 0.00939545f $X=3.055 $Y=1.075 $X2=2.84
+ $Y2=1.595
cc_235 N_A_27_115#_M1011_g N_Y_c_391_n 0.00251111f $X=2.625 $Y=1.075 $X2=2.84
+ $Y2=2.845
cc_236 N_A_27_115#_c_213_n N_Y_c_391_n 0.0185925f $X=2.625 $Y=2.86 $X2=2.84
+ $Y2=2.845
cc_237 N_A_27_115#_c_251_n N_Y_c_391_n 0.00113627f $X=2.625 $Y=3.01 $X2=2.84
+ $Y2=2.845
cc_238 N_A_27_115#_c_214_n N_Y_c_391_n 0.0170354f $X=2.98 $Y=1.845 $X2=2.84
+ $Y2=2.845
cc_239 N_A_27_115#_c_215_n N_Y_c_391_n 0.00966211f $X=2.98 $Y=2.935 $X2=2.84
+ $Y2=2.845
cc_240 N_A_27_115#_M1013_g N_Y_c_391_n 0.00251111f $X=3.055 $Y=1.075 $X2=2.84
+ $Y2=2.845
cc_241 N_A_27_115#_c_255_n N_Y_c_391_n 0.0031083f $X=3.055 $Y=3.01 $X2=2.84
+ $Y2=2.845
cc_242 N_A_27_115#_c_224_n N_Y_c_391_n 6.59375e-19 $X=2.625 $Y=2.935 $X2=2.84
+ $Y2=2.845
cc_243 N_A_27_115#_M1000_g GND 0.00468827f $X=0.905 $Y=1.075 $X2=0.34 $Y2=0.22
cc_244 N_A_27_115#_M1001_g GND 0.00468827f $X=1.335 $Y=1.075 $X2=0.34 $Y2=0.22
cc_245 N_A_27_115#_M1008_g GND 0.00468827f $X=1.765 $Y=1.075 $X2=0.34 $Y2=0.22
cc_246 N_A_27_115#_M1010_g GND 0.00468827f $X=2.195 $Y=1.075 $X2=0.34 $Y2=0.22
cc_247 N_A_27_115#_M1011_g GND 0.00468827f $X=2.625 $Y=1.075 $X2=0.34 $Y2=0.22
cc_248 N_A_27_115#_M1013_g GND 0.00468827f $X=3.055 $Y=1.075 $X2=0.34 $Y2=0.22
cc_249 N_A_27_115#_c_225_n GND 0.00476261f $X=0.26 $Y=0.825 $X2=0.34 $Y2=0.22
cc_250 N_A_27_115#_c_232_n VDD 0.00468827f $X=0.905 $Y=3.01 $X2=0.34 $Y2=6.44
cc_251 N_A_27_115#_c_235_n VDD 0.00470215f $X=1.335 $Y=3.01 $X2=0.34 $Y2=6.44
cc_252 N_A_27_115#_c_242_n VDD 0.00468827f $X=1.765 $Y=3.01 $X2=0.34 $Y2=6.44
cc_253 N_A_27_115#_c_246_n VDD 0.00468827f $X=2.195 $Y=3.01 $X2=0.34 $Y2=6.44
cc_254 N_A_27_115#_c_251_n VDD 0.00468827f $X=2.625 $Y=3.01 $X2=0.34 $Y2=6.44
cc_255 N_A_27_115#_c_255_n VDD 0.00468827f $X=3.055 $Y=3.01 $X2=0.34 $Y2=6.44
cc_256 N_A_27_115#_c_227_n VDD 0.00476261f $X=0.26 $Y=3.455 $X2=0.34 $Y2=6.44
cc_257 N_Y_c_364_n GND 0.00475776f $X=1.12 $Y=0.825 $X2=0.34 $Y2=0.22
cc_258 N_Y_c_367_n GND 0.00475776f $X=1.98 $Y=0.825 $X2=0.34 $Y2=0.22
cc_259 N_Y_c_371_n GND 0.00475776f $X=2.84 $Y=0.825 $X2=0.34 $Y2=0.22
cc_260 N_Y_c_392_n VDD 0.00475776f $X=1.12 $Y=2.96 $X2=0.34 $Y2=6.44
cc_261 N_Y_c_394_n VDD 0.00475776f $X=1.98 $Y=2.96 $X2=0.34 $Y2=6.44
cc_262 N_Y_c_396_n VDD 0.00475776f $X=2.84 $Y=2.96 $X2=0.34 $Y2=6.44
