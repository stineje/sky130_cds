* File: sky130_osu_sc_18T_hs__dffsr_1.spice
* Created: Fri Nov 12 13:49:33 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_hs__dffsr_1.pex.spice"
.subckt sky130_osu_sc_18T_hs__dffsr_1  GND VDD RN SN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* RN	RN
* VDD	VDD
* GND	GND
MM1021 N_A_110_115#_M1021_d N_RN_M1021_g N_GND_M1021_s N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1033 N_A_217_617#_M1033_d N_A_110_115#_M1033_g N_GND_M1033_s N_GND_M1021_b
+ NLOWVT L=0.15 W=0.74 AD=0.136305 AS=0.1961 PD=1.13977 PS=2.01 NRD=9.72 NRS=0
+ M=1 R=4.93333 SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1018 A_400_115# N_SN_M1018_g N_A_217_617#_M1033_d N_GND_M1021_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.184195 PD=1.21 PS=1.54023 NRD=5.988 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1006 N_GND_M1006_d N_A_432_520#_M1006_g A_400_115# N_GND_M1021_b NLOWVT L=0.15
+ W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 A_662_115# N_D_M1009_g N_GND_M1009_s N_GND_M1021_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1035 N_A_432_520#_M1035_d N_A_704_89#_M1035_g A_662_115# N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1
+ R=6.66667 SA=75000.5 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1031 A_854_115# N_CK_M1031_g N_A_432_520#_M1035_d N_GND_M1021_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.1 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1025 N_GND_M1025_d N_A_217_617#_M1025_g A_854_115# N_GND_M1021_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.5
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1029 A_1012_115# N_A_217_617#_M1029_g N_GND_M1025_d N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1026 N_A_1084_115#_M1026_d N_CK_M1026_g A_1012_115# N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1
+ R=6.66667 SA=75002.3 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1022 A_1204_115# N_A_704_89#_M1022_g N_A_1084_115#_M1026_d N_GND_M1021_b
+ NLOWVT L=0.15 W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1
+ R=6.66667 SA=75002.9 SB=75001 A=0.15 P=2.3 MULT=1
MM1010 N_GND_M1010_d N_A_1246_89#_M1010_g A_1204_115# N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667
+ SA=75003.3 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_A_704_89#_M1015_d N_CK_M1015_g N_GND_M1010_d N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1016 A_1552_115# N_A_1084_115#_M1016_g N_GND_M1016_s N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1007 N_A_1246_89#_M1007_d N_SN_M1007_g A_1552_115# N_GND_M1021_b NLOWVT L=0.15
+ W=1 AD=0.184195 AS=0.105 PD=1.54023 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667
+ SA=75000.5 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1027 N_GND_M1027_d N_A_110_115#_M1027_g N_A_1246_89#_M1007_d N_GND_M1021_b
+ NLOWVT L=0.15 W=0.74 AD=0.1961 AS=0.136305 PD=2.01 PS=1.13977 NRD=0 NRS=9.72
+ M=1 R=4.93333 SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_GND_M1011_d N_A_1246_89#_M1011_g N_QN_M1011_s N_GND_M1021_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_Q_M1013_d N_QN_M1013_g N_GND_M1011_d N_GND_M1021_b NLOWVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1019 N_A_110_115#_M1019_d N_RN_M1019_g N_VDD_M1019_s N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1017 N_A_300_617#_M1017_d N_A_110_115#_M1017_g N_A_217_617#_M1017_s
+ N_VDD_M1019_b PSHORT L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0
+ M=1 R=20 SA=75000.2 SB=75001 A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_SN_M1000_g N_A_300_617#_M1017_d N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1001 N_A_300_617#_M1001_d N_A_432_520#_M1001_g N_VDD_M1000_d N_VDD_M1019_b
+ PSHORT L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20
+ SA=75001 SB=75000.2 A=0.45 P=6.3 MULT=1
MM1003 A_662_617# N_D_M1003_g N_VDD_M1003_s N_VDD_M1019_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.2
+ SB=75003.7 A=0.45 P=6.3 MULT=1
MM1032 N_A_432_520#_M1032_d N_CK_M1032_g A_662_617# N_VDD_M1019_b PSHORT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75000.5 SB=75003.3 A=0.45 P=6.3 MULT=1
MM1030 A_854_617# N_A_704_89#_M1030_g N_A_432_520#_M1032_d N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75001.1 SB=75002.7 A=0.45 P=6.3 MULT=1
MM1023 N_VDD_M1023_d N_A_217_617#_M1023_g A_854_617# N_VDD_M1019_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.5
+ SB=75002.4 A=0.45 P=6.3 MULT=1
MM1028 A_1012_617# N_A_217_617#_M1028_g N_VDD_M1023_d N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20
+ SA=75001.9 SB=75001.9 A=0.45 P=6.3 MULT=1
MM1024 N_A_1084_115#_M1024_d N_A_704_89#_M1024_g A_1012_617# N_VDD_M1019_b
+ PSHORT L=0.15 W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1
+ R=20 SA=75002.3 SB=75001.6 A=0.45 P=6.3 MULT=1
MM1020 A_1204_617# N_CK_M1020_g N_A_1084_115#_M1024_d N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75002.9 SB=75001 A=0.45 P=6.3 MULT=1
MM1004 N_VDD_M1004_d N_A_1246_89#_M1004_g A_1204_617# N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20
+ SA=75003.3 SB=75000.6 A=0.45 P=6.3 MULT=1
MM1012 N_A_704_89#_M1012_d N_CK_M1012_g N_VDD_M1004_d N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.7
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1014 N_VDD_M1014_d N_A_1084_115#_M1014_g N_A_1469_617#_M1014_s N_VDD_M1019_b
+ PSHORT L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20
+ SA=75000.2 SB=75001 A=0.45 P=6.3 MULT=1
MM1034 N_A_1469_617#_M1034_d N_SN_M1034_g N_VDD_M1014_d N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1002 N_A_1246_89#_M1002_d N_A_110_115#_M1002_g N_A_1469_617#_M1034_d
+ N_VDD_M1019_b PSHORT L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0
+ M=1 R=20 SA=75001 SB=75000.2 A=0.45 P=6.3 MULT=1
MM1005 N_VDD_M1005_d N_A_1246_89#_M1005_g N_QN_M1005_s N_VDD_M1019_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1008 N_Q_M1008_d N_QN_M1008_g N_VDD_M1005_d N_VDD_M1019_b PSHORT L=0.15 W=3
+ AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX36_noxref N_GND_M1021_b N_VDD_M1019_b NWDIODE A=39.9 P=28.6
pX37_noxref noxref_27 RN RN PROBETYPE=1
pX38_noxref noxref_28 D D PROBETYPE=1
pX39_noxref noxref_29 CK CK PROBETYPE=1
pX40_noxref noxref_30 SN SN PROBETYPE=1
pX41_noxref noxref_31 QN QN PROBETYPE=1
pX42_noxref noxref_32 Q Q PROBETYPE=1
c_1965 A_1012_617# 0 1.57671e-19 $X=5.06 $Y=3.085
*
.include "sky130_osu_sc_18T_hs__dffsr_1.pxi.spice"
*
.ends
*
*
