magic
tech sky130A
magscale 1 2
timestamp 1641997726
<< nwell >>
rect 50 1089 330 1090
rect 50 529 1020 1089
<< nmoslvt >>
rect 171 115 201 263
rect 257 115 287 263
rect 329 115 359 263
rect 449 115 479 263
rect 521 115 551 263
rect 607 115 637 263
rect 815 115 845 263
rect 901 115 931 263
<< pmos >>
rect 171 565 201 965
rect 257 565 287 965
rect 329 565 359 965
rect 449 565 479 965
rect 521 565 551 965
rect 607 565 637 965
rect 815 565 845 965
rect 901 565 931 965
<< ndiff >>
rect 118 215 171 263
rect 118 131 126 215
rect 160 131 171 215
rect 118 115 171 131
rect 201 215 257 263
rect 201 131 212 215
rect 246 131 257 215
rect 201 115 257 131
rect 287 115 329 263
rect 359 215 449 263
rect 359 131 370 215
rect 438 131 449 215
rect 359 115 449 131
rect 479 115 521 263
rect 551 215 607 263
rect 551 131 562 215
rect 596 131 607 215
rect 551 115 607 131
rect 637 215 690 263
rect 637 131 648 215
rect 682 131 690 215
rect 637 115 690 131
rect 762 215 815 263
rect 762 131 770 215
rect 804 131 815 215
rect 762 115 815 131
rect 845 215 901 263
rect 845 131 856 215
rect 890 131 901 215
rect 845 115 901 131
rect 931 215 984 263
rect 931 131 942 215
rect 976 131 984 215
rect 931 115 984 131
<< pdiff >>
rect 118 949 171 965
rect 118 673 126 949
rect 160 673 171 949
rect 118 565 171 673
rect 201 949 257 965
rect 201 673 212 949
rect 246 673 257 949
rect 201 565 257 673
rect 287 565 329 965
rect 359 949 449 965
rect 359 605 370 949
rect 438 605 449 949
rect 359 565 449 605
rect 479 565 521 965
rect 551 949 607 965
rect 551 605 562 949
rect 596 605 607 949
rect 551 565 607 605
rect 637 949 690 965
rect 637 605 648 949
rect 682 605 690 949
rect 637 565 690 605
rect 762 949 815 965
rect 762 605 770 949
rect 804 605 815 949
rect 762 565 815 605
rect 845 949 901 965
rect 845 605 856 949
rect 890 605 901 949
rect 845 565 901 605
rect 931 949 984 965
rect 931 605 942 949
rect 976 605 984 949
rect 931 565 984 605
<< ndiffc >>
rect 126 131 160 215
rect 212 131 246 215
rect 370 131 438 215
rect 562 131 596 215
rect 648 131 682 215
rect 770 131 804 215
rect 856 131 890 215
rect 942 131 976 215
<< pdiffc >>
rect 126 673 160 949
rect 212 673 246 949
rect 370 605 438 949
rect 562 605 596 949
rect 648 605 682 949
rect 770 605 804 949
rect 856 605 890 949
rect 942 605 976 949
<< psubdiff >>
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
<< nsubdiff >>
rect 163 1019 187 1053
rect 221 1019 245 1053
rect 299 1019 323 1053
rect 357 1019 381 1053
rect 435 1019 459 1053
rect 493 1019 517 1053
rect 571 1019 595 1053
rect 629 1019 653 1053
rect 707 1019 731 1053
rect 765 1019 789 1053
rect 843 1019 867 1053
rect 901 1019 925 1053
<< psubdiffcont >>
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
<< nsubdiffcont >>
rect 187 1019 221 1053
rect 323 1019 357 1053
rect 459 1019 493 1053
rect 595 1019 629 1053
rect 731 1019 765 1053
rect 867 1019 901 1053
<< poly >>
rect 171 965 201 991
rect 257 965 287 991
rect 329 965 359 991
rect 449 965 479 991
rect 521 965 551 991
rect 607 965 637 991
rect 815 965 845 991
rect 901 965 931 991
rect 171 543 201 565
rect 161 509 201 543
rect 161 351 191 509
rect 257 466 287 565
rect 329 534 359 565
rect 449 534 479 565
rect 329 518 383 534
rect 329 484 339 518
rect 373 484 383 518
rect 329 468 383 484
rect 425 518 479 534
rect 425 484 435 518
rect 469 484 479 518
rect 425 468 479 484
rect 233 450 287 466
rect 233 416 243 450
rect 277 416 287 450
rect 425 423 455 468
rect 233 400 287 416
rect 161 335 215 351
rect 161 301 171 335
rect 205 301 215 335
rect 161 285 215 301
rect 171 263 201 285
rect 257 263 287 400
rect 329 393 455 423
rect 521 425 551 565
rect 607 534 637 565
rect 815 549 845 565
rect 607 504 648 534
rect 521 409 575 425
rect 329 263 359 393
rect 521 375 531 409
rect 565 375 575 409
rect 521 359 575 375
rect 425 335 479 351
rect 425 301 435 335
rect 469 301 479 335
rect 425 285 479 301
rect 449 263 479 285
rect 521 263 551 359
rect 618 351 648 504
rect 805 519 845 549
rect 805 425 835 519
rect 901 425 931 565
rect 780 409 835 425
rect 780 375 790 409
rect 824 375 835 409
rect 780 359 835 375
rect 877 409 931 425
rect 877 375 887 409
rect 921 375 931 409
rect 877 359 931 375
rect 618 335 680 351
rect 618 311 632 335
rect 607 301 632 311
rect 666 301 680 335
rect 607 281 680 301
rect 805 308 835 359
rect 607 263 637 281
rect 805 278 845 308
rect 815 263 845 278
rect 901 263 931 359
rect 171 89 201 115
rect 257 89 287 115
rect 329 89 359 115
rect 449 89 479 115
rect 521 89 551 115
rect 607 89 637 115
rect 815 89 845 115
rect 901 89 931 115
<< polycont >>
rect 339 484 373 518
rect 435 484 469 518
rect 243 416 277 450
rect 171 301 205 335
rect 531 375 565 409
rect 435 301 469 335
rect 790 375 824 409
rect 887 375 921 409
rect 632 301 666 335
<< locali >>
rect 50 1059 1018 1080
rect 50 1019 187 1059
rect 221 1019 323 1059
rect 357 1019 459 1059
rect 493 1019 595 1059
rect 629 1019 731 1059
rect 765 1019 867 1059
rect 901 1019 1018 1059
rect 126 949 160 965
rect 103 673 126 739
rect 103 656 160 673
rect 212 949 246 1019
rect 212 657 246 673
rect 370 949 438 965
rect 103 409 137 656
rect 370 602 438 605
rect 103 244 137 375
rect 171 568 438 602
rect 562 949 596 1019
rect 562 589 596 605
rect 648 949 682 965
rect 171 335 205 568
rect 435 518 469 534
rect 323 484 339 518
rect 373 484 389 518
rect 243 400 277 416
rect 355 335 389 484
rect 435 483 469 484
rect 648 483 682 605
rect 770 949 804 965
rect 770 557 804 605
rect 856 949 890 1019
rect 856 589 890 605
rect 942 949 976 965
rect 976 597 989 614
rect 942 580 989 597
rect 770 518 804 523
rect 770 484 921 518
rect 648 419 682 449
rect 515 375 531 409
rect 565 375 581 409
rect 648 385 736 419
rect 887 409 921 484
rect 632 335 666 351
rect 205 301 314 335
rect 355 301 435 335
rect 469 301 485 335
rect 171 285 205 301
rect 280 251 314 301
rect 632 285 666 301
rect 103 215 160 244
rect 103 210 126 215
rect 126 115 160 131
rect 212 215 246 231
rect 280 217 438 251
rect 702 249 736 385
rect 774 375 790 409
rect 824 375 840 409
rect 887 335 921 375
rect 212 61 246 131
rect 370 215 438 217
rect 370 115 438 131
rect 562 215 596 231
rect 562 61 596 131
rect 648 215 736 249
rect 770 301 921 335
rect 770 215 804 301
rect 955 267 989 580
rect 942 233 989 267
rect 648 115 682 131
rect 770 115 804 131
rect 856 215 890 231
rect 856 61 890 131
rect 942 215 976 233
rect 942 115 976 131
rect 50 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1018 61
rect 50 0 1018 21
<< viali >>
rect 187 1053 221 1059
rect 187 1025 221 1053
rect 323 1053 357 1059
rect 323 1025 357 1053
rect 459 1053 493 1059
rect 459 1025 493 1053
rect 595 1053 629 1059
rect 595 1025 629 1053
rect 731 1053 765 1059
rect 731 1025 765 1053
rect 867 1053 901 1059
rect 867 1025 901 1053
rect 103 375 137 409
rect 243 450 277 484
rect 435 449 469 483
rect 942 605 976 631
rect 942 597 976 605
rect 770 523 804 557
rect 648 449 682 483
rect 531 375 565 409
rect 435 301 469 335
rect 632 301 666 335
rect 790 375 824 409
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
<< metal1 >>
rect 50 1059 1018 1080
rect 50 1025 187 1059
rect 221 1025 323 1059
rect 357 1025 459 1059
rect 493 1025 595 1059
rect 629 1025 731 1059
rect 765 1025 867 1059
rect 901 1025 1018 1059
rect 50 1019 1018 1025
rect 930 631 988 637
rect 907 597 942 631
rect 976 597 988 631
rect 930 591 988 597
rect 758 557 816 563
rect 751 556 770 557
rect 736 524 770 556
rect 751 523 770 524
rect 804 523 816 557
rect 758 517 816 523
rect 231 484 290 490
rect 231 450 243 484
rect 277 450 310 484
rect 423 483 481 489
rect 636 483 694 489
rect 231 444 290 450
rect 423 449 435 483
rect 469 449 648 483
rect 682 449 694 483
rect 423 443 481 449
rect 636 443 694 449
rect 90 409 149 415
rect 90 375 103 409
rect 137 402 149 409
rect 519 409 578 415
rect 519 402 531 409
rect 137 375 531 402
rect 565 406 578 409
rect 778 409 836 415
rect 778 406 790 409
rect 565 378 790 406
rect 565 375 578 378
rect 90 374 578 375
rect 90 369 149 374
rect 519 369 578 374
rect 778 375 790 378
rect 824 375 836 409
rect 778 369 836 375
rect 423 335 482 342
rect 615 336 674 341
rect 615 335 683 336
rect 400 301 435 335
rect 469 301 632 335
rect 666 301 683 335
rect 423 295 482 301
rect 615 294 674 301
rect 50 55 1018 61
rect 50 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1018 55
rect 50 0 1018 21
<< labels >>
rlabel viali 260 466 260 466 1 D
port 1 n
rlabel viali 959 614 959 614 1 Q
port 2 n
rlabel viali 788 540 788 540 1 QN
port 3 n
rlabel viali 452 318 452 318 1 CK
port 4 n
rlabel nwell 204 1041 208 1042 1 vdd
rlabel nwell 342 1043 346 1044 1 vdd
rlabel viali 476 1043 476 1043 1 vdd
rlabel viali 611 1045 611 1045 1 vdd
rlabel viali 747 1046 747 1046 1 vdd
rlabel viali 885 1044 885 1044 1 vdd
rlabel viali 204 42 204 42 1 gnd
rlabel viali 337 38 337 38 1 gnd
rlabel viali 475 36 475 36 1 gnd
rlabel viali 611 36 611 36 1 gnd
rlabel viali 745 34 745 34 1 gnd
rlabel viali 886 34 886 34 1 gnd
<< end >>
