magic
tech sky130A
magscale 1 2
timestamp 1612373629
<< nwell >>
rect -9 529 462 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 252 115 282 243
rect 338 115 368 243
<< pmos >>
rect 80 565 110 965
rect 152 565 182 965
rect 252 565 282 965
rect 324 565 354 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 165 166 243
rect 110 131 121 165
rect 155 131 166 165
rect 110 115 166 131
rect 196 215 252 243
rect 196 131 207 215
rect 241 131 252 215
rect 196 115 252 131
rect 282 215 338 243
rect 282 181 293 215
rect 327 181 338 215
rect 282 115 338 181
rect 368 165 421 243
rect 368 131 379 165
rect 413 131 421 165
rect 368 115 421 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 565 152 965
rect 182 949 252 965
rect 182 673 200 949
rect 234 673 252 949
rect 182 565 252 673
rect 282 565 324 965
rect 354 949 407 965
rect 354 741 365 949
rect 399 741 407 949
rect 354 565 407 741
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 165
rect 207 131 241 215
rect 293 181 327 215
rect 379 131 413 165
<< pdiffc >>
rect 35 741 69 949
rect 200 673 234 949
rect 365 741 399 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
<< poly >>
rect 80 965 110 991
rect 152 965 182 991
rect 252 965 282 991
rect 324 965 354 991
rect 80 533 110 565
rect 56 517 110 533
rect 56 483 66 517
rect 100 483 110 517
rect 56 467 110 483
rect 56 318 86 467
rect 152 419 182 565
rect 130 409 196 419
rect 130 375 146 409
rect 180 375 196 409
rect 130 365 196 375
rect 56 288 110 318
rect 80 243 110 288
rect 166 243 196 365
rect 252 361 282 565
rect 324 540 354 565
rect 324 510 368 540
rect 338 426 368 510
rect 338 410 430 426
rect 338 376 384 410
rect 418 376 430 410
rect 238 345 292 361
rect 238 311 248 345
rect 282 311 292 345
rect 238 295 292 311
rect 338 360 430 376
rect 252 243 282 295
rect 338 243 368 360
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
rect 338 89 368 115
<< polycont >>
rect 66 483 100 517
rect 146 375 180 409
rect 384 376 418 410
rect 248 311 282 345
<< locali >>
rect 0 1089 462 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 462 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 200 949 234 965
rect 365 949 399 1049
rect 365 725 399 741
rect 200 648 234 673
rect 200 614 350 648
rect 66 517 100 597
rect 66 467 100 483
rect 146 523 162 557
rect 146 409 180 523
rect 146 359 180 375
rect 223 361 257 449
rect 223 345 282 361
rect 223 311 248 345
rect 223 295 282 311
rect 316 335 350 614
rect 384 410 418 426
rect 384 360 418 376
rect 35 215 241 249
rect 35 115 69 131
rect 121 165 155 181
rect 121 61 155 131
rect 293 227 316 261
rect 293 215 327 227
rect 293 165 327 181
rect 379 165 413 181
rect 207 129 241 131
rect 379 129 413 131
rect 207 95 413 129
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 462 61
rect 0 0 462 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 66 597 100 631
rect 162 523 196 557
rect 223 449 257 483
rect 384 376 418 410
rect 316 301 350 335
rect 316 227 350 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
<< metal1 >>
rect 0 1089 462 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 462 1089
rect 0 1049 462 1055
rect 54 631 112 637
rect 54 597 66 631
rect 100 597 134 631
rect 54 591 112 597
rect 150 557 208 563
rect 150 523 162 557
rect 196 523 230 557
rect 150 517 208 523
rect 211 483 269 489
rect 189 449 223 483
rect 257 449 269 483
rect 211 443 269 449
rect 372 410 430 416
rect 350 376 384 410
rect 418 376 430 410
rect 372 370 430 376
rect 304 335 362 341
rect 304 301 316 335
rect 350 301 362 335
rect 304 295 362 301
rect 316 267 350 295
rect 304 261 362 267
rect 304 227 316 261
rect 350 227 362 261
rect 304 221 362 227
rect 0 55 462 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 462 55
rect 0 0 462 21
<< labels >>
rlabel viali 240 466 240 466 1 B0
port 4 n
rlabel viali 179 540 179 540 1 A1
port 2 n
rlabel viali 83 614 83 614 1 A0
port 1 n
rlabel viali 333 318 333 318 1 Y
port 3 n
rlabel viali 401 393 401 393 1 B1
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
