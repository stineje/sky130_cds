* File: sky130_osu_sc_12T_ls__buf_6.pxi.spice
* Created: Fri Nov 12 15:35:22 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__BUF_6%noxref_1 N_noxref_1_M1006_d N_noxref_1_M1001_s
+ N_noxref_1_M1010_s N_noxref_1_M1013_s N_noxref_1_M1006_b N_noxref_1_c_2_p
+ N_noxref_1_c_3_p N_noxref_1_c_9_p N_noxref_1_c_13_p N_noxref_1_c_21_p
+ N_noxref_1_c_26_p N_noxref_1_c_32_p N_noxref_1_c_38_p N_noxref_1_c_92_p
+ N_noxref_1_c_93_p PM_SKY130_OSU_SC_12T_LS__BUF_6%noxref_1
x_PM_SKY130_OSU_SC_12T_LS__BUF_6%noxref_2 N_noxref_2_M1004_d N_noxref_2_M1003_s
+ N_noxref_2_M1007_s N_noxref_2_M1012_s N_noxref_2_M1004_b N_noxref_2_c_95_p
+ N_noxref_2_c_96_p N_noxref_2_c_104_p N_noxref_2_c_108_p N_noxref_2_c_114_p
+ N_noxref_2_c_118_p N_noxref_2_c_123_p N_noxref_2_c_127_p N_noxref_2_c_151_p
+ N_noxref_2_c_152_p N_noxref_2_c_153_p PM_SKY130_OSU_SC_12T_LS__BUF_6%noxref_2
x_PM_SKY130_OSU_SC_12T_LS__BUF_6%A N_A_M1006_g N_A_M1004_g N_A_c_158_n
+ N_A_c_159_n A PM_SKY130_OSU_SC_12T_LS__BUF_6%A
x_PM_SKY130_OSU_SC_12T_LS__BUF_6%A_27_115# N_A_27_115#_M1006_s
+ N_A_27_115#_M1004_s N_A_27_115#_M1000_g N_A_27_115#_c_239_n
+ N_A_27_115#_M1002_g N_A_27_115#_c_197_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_242_n N_A_27_115#_M1003_g N_A_27_115#_c_201_n
+ N_A_27_115#_c_203_n N_A_27_115#_c_204_n N_A_27_115#_c_205_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_249_n N_A_27_115#_M1005_g
+ N_A_27_115#_c_209_n N_A_27_115#_c_210_n N_A_27_115#_M1010_g
+ N_A_27_115#_c_253_n N_A_27_115#_M1007_g N_A_27_115#_c_214_n
+ N_A_27_115#_c_216_n N_A_27_115#_M1011_g N_A_27_115#_c_220_n
+ N_A_27_115#_c_258_n N_A_27_115#_M1009_g N_A_27_115#_c_221_n
+ N_A_27_115#_c_222_n N_A_27_115#_M1013_g N_A_27_115#_c_262_n
+ N_A_27_115#_M1012_g N_A_27_115#_c_226_n N_A_27_115#_c_227_n
+ N_A_27_115#_c_228_n N_A_27_115#_c_229_n N_A_27_115#_c_230_n
+ N_A_27_115#_c_231_n N_A_27_115#_c_232_n N_A_27_115#_c_234_n
+ N_A_27_115#_c_235_n N_A_27_115#_c_237_n N_A_27_115#_c_238_n
+ PM_SKY130_OSU_SC_12T_LS__BUF_6%A_27_115#
x_PM_SKY130_OSU_SC_12T_LS__BUF_6%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1011_d
+ N_Y_M1002_d N_Y_M1005_d N_Y_M1009_d N_Y_c_371_n N_Y_c_406_n N_Y_c_374_n
+ N_Y_c_408_n N_Y_c_378_n N_Y_c_410_n N_Y_c_381_n N_Y_c_385_n Y N_Y_c_387_n
+ N_Y_c_413_n N_Y_c_391_n N_Y_c_392_n N_Y_c_396_n N_Y_c_415_n N_Y_c_400_n
+ N_Y_c_401_n N_Y_c_405_n PM_SKY130_OSU_SC_12T_LS__BUF_6%Y
cc_1 N_noxref_1_M1006_b N_A_M1006_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=0.835
cc_2 N_noxref_1_c_2_p N_A_M1006_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475
+ $Y2=0.835
cc_3 N_noxref_1_c_3_p N_A_M1006_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.475
+ $Y2=0.835
cc_4 N_noxref_1_M1006_b N_A_M1004_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=3.235
cc_5 N_noxref_1_M1006_b N_A_c_158_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_6 N_noxref_1_M1006_b N_A_c_159_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_7 N_noxref_1_M1006_b N_A_27_115#_M1000_g 0.0207501f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.835
cc_8 N_noxref_1_c_3_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.905
+ $Y2=0.835
cc_9 N_noxref_1_c_9_p N_A_27_115#_M1000_g 0.00606474f $X=1.465 $Y=0.152
+ $X2=0.905 $Y2=0.835
cc_10 N_noxref_1_M1006_b N_A_27_115#_c_197_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.38
cc_11 N_noxref_1_M1006_b N_A_27_115#_M1001_g 0.020212f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.835
cc_12 N_noxref_1_c_9_p N_A_27_115#_M1001_g 0.00606474f $X=1.465 $Y=0.152
+ $X2=1.335 $Y2=0.835
cc_13 N_noxref_1_c_13_p N_A_27_115#_M1001_g 0.00311745f $X=1.55 $Y=0.755
+ $X2=1.335 $Y2=0.835
cc_14 N_noxref_1_M1006_b N_A_27_115#_c_201_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.365
cc_15 N_noxref_1_c_13_p N_A_27_115#_c_201_n 0.00256938f $X=1.55 $Y=0.755
+ $X2=1.69 $Y2=1.365
cc_16 N_noxref_1_M1006_b N_A_27_115#_c_203_n 0.0429274f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.365
cc_17 N_noxref_1_M1006_b N_A_27_115#_c_204_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.455
cc_18 N_noxref_1_M1006_b N_A_27_115#_c_205_n 0.0196789f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.455
cc_19 N_noxref_1_M1006_b N_A_27_115#_M1008_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.835
cc_20 N_noxref_1_c_13_p N_A_27_115#_M1008_g 0.00311745f $X=1.55 $Y=0.755
+ $X2=1.765 $Y2=0.835
cc_21 N_noxref_1_c_21_p N_A_27_115#_M1008_g 0.00606474f $X=2.325 $Y=0.152
+ $X2=1.765 $Y2=0.835
cc_22 N_noxref_1_M1006_b N_A_27_115#_c_209_n 0.0195339f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.365
cc_23 N_noxref_1_M1006_b N_A_27_115#_c_210_n 0.0107618f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.455
cc_24 N_noxref_1_M1006_b N_A_27_115#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.835
cc_25 N_noxref_1_c_21_p N_A_27_115#_M1010_g 0.00606474f $X=2.325 $Y=0.152
+ $X2=2.195 $Y2=0.835
cc_26 N_noxref_1_c_26_p N_A_27_115#_M1010_g 0.00311745f $X=2.41 $Y=0.755
+ $X2=2.195 $Y2=0.835
cc_27 N_noxref_1_M1006_b N_A_27_115#_c_214_n 0.0165886f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.365
cc_28 N_noxref_1_c_26_p N_A_27_115#_c_214_n 0.00256938f $X=2.41 $Y=0.755
+ $X2=2.55 $Y2=1.365
cc_29 N_noxref_1_M1006_b N_A_27_115#_c_216_n 0.0109555f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.455
cc_30 N_noxref_1_M1006_b N_A_27_115#_M1011_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.835
cc_31 N_noxref_1_c_26_p N_A_27_115#_M1011_g 0.00311745f $X=2.41 $Y=0.755
+ $X2=2.625 $Y2=0.835
cc_32 N_noxref_1_c_32_p N_A_27_115#_M1011_g 0.00606474f $X=3.185 $Y=0.152
+ $X2=2.625 $Y2=0.835
cc_33 N_noxref_1_M1006_b N_A_27_115#_c_220_n 0.0668243f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.38
cc_34 N_noxref_1_M1006_b N_A_27_115#_c_221_n 0.0385034f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.365
cc_35 N_noxref_1_M1006_b N_A_27_115#_c_222_n 0.0221499f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.455
cc_36 N_noxref_1_M1006_b N_A_27_115#_M1013_g 0.0264941f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.835
cc_37 N_noxref_1_c_32_p N_A_27_115#_M1013_g 0.00606474f $X=3.185 $Y=0.152
+ $X2=3.055 $Y2=0.835
cc_38 N_noxref_1_c_38_p N_A_27_115#_M1013_g 0.00502587f $X=3.27 $Y=0.755
+ $X2=3.055 $Y2=0.835
cc_39 N_noxref_1_M1006_b N_A_27_115#_c_226_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.365
cc_40 N_noxref_1_M1006_b N_A_27_115#_c_227_n 0.00890086f $X=-0.045 $Y=0
+ $X2=1.765 $Y2=2.455
cc_41 N_noxref_1_M1006_b N_A_27_115#_c_228_n 0.0106787f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.365
cc_42 N_noxref_1_M1006_b N_A_27_115#_c_229_n 0.00890086f $X=-0.045 $Y=0
+ $X2=2.195 $Y2=2.455
cc_43 N_noxref_1_M1006_b N_A_27_115#_c_230_n 0.0023879f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.365
cc_44 N_noxref_1_M1006_b N_A_27_115#_c_231_n 7.16371e-19 $X=-0.045 $Y=0
+ $X2=2.625 $Y2=2.455
cc_45 N_noxref_1_M1006_b N_A_27_115#_c_232_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_46 N_noxref_1_c_2_p N_A_27_115#_c_232_n 0.00736239f $X=0.605 $Y=0.152
+ $X2=0.26 $Y2=0.755
cc_47 N_noxref_1_M1006_b N_A_27_115#_c_234_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.955
cc_48 N_noxref_1_M1006_b N_A_27_115#_c_235_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.455
cc_49 N_noxref_1_c_3_p N_A_27_115#_c_235_n 0.00702738f $X=0.69 $Y=0.755 $X2=0.88
+ $Y2=1.455
cc_50 N_noxref_1_M1006_b N_A_27_115#_c_237_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.455
cc_51 N_noxref_1_M1006_b N_A_27_115#_c_238_n 0.00592383f $X=-0.045 $Y=0
+ $X2=0.965 $Y2=1.455
cc_52 N_noxref_1_M1006_b N_Y_c_371_n 0.00154299f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.755
cc_53 N_noxref_1_c_9_p N_Y_c_371_n 0.00718527f $X=1.465 $Y=0.152 $X2=1.12
+ $Y2=0.755
cc_54 N_noxref_1_c_13_p N_Y_c_371_n 8.14297e-19 $X=1.55 $Y=0.755 $X2=1.12
+ $Y2=0.755
cc_55 N_noxref_1_M1006_b N_Y_c_374_n 0.00154299f $X=-0.045 $Y=0 $X2=1.98
+ $Y2=0.755
cc_56 N_noxref_1_c_13_p N_Y_c_374_n 8.14297e-19 $X=1.55 $Y=0.755 $X2=1.98
+ $Y2=0.755
cc_57 N_noxref_1_c_21_p N_Y_c_374_n 0.00738926f $X=2.325 $Y=0.152 $X2=1.98
+ $Y2=0.755
cc_58 N_noxref_1_c_26_p N_Y_c_374_n 8.14297e-19 $X=2.41 $Y=0.755 $X2=1.98
+ $Y2=0.755
cc_59 N_noxref_1_M1006_b N_Y_c_378_n 0.00154299f $X=-0.045 $Y=0 $X2=2.84
+ $Y2=0.755
cc_60 N_noxref_1_c_26_p N_Y_c_378_n 8.14297e-19 $X=2.41 $Y=0.755 $X2=2.84
+ $Y2=0.755
cc_61 N_noxref_1_c_32_p N_Y_c_378_n 0.00731228f $X=3.185 $Y=0.152 $X2=2.84
+ $Y2=0.755
cc_62 N_noxref_1_M1006_b N_Y_c_381_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=1.115
cc_63 N_noxref_1_c_3_p N_Y_c_381_n 0.00134236f $X=0.69 $Y=0.755 $X2=1.12
+ $Y2=1.115
cc_64 N_noxref_1_c_9_p N_Y_c_381_n 0.00245319f $X=1.465 $Y=0.152 $X2=1.12
+ $Y2=1.115
cc_65 N_noxref_1_c_13_p N_Y_c_381_n 7.53951e-19 $X=1.55 $Y=0.755 $X2=1.12
+ $Y2=1.115
cc_66 N_noxref_1_M1006_b N_Y_c_385_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=2.365
cc_67 N_noxref_1_M1006_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=1.79
cc_68 N_noxref_1_M1001_s N_Y_c_387_n 0.0100329f $X=1.41 $Y=0.575 $X2=1.835 $Y2=1
cc_69 N_noxref_1_c_9_p N_Y_c_387_n 0.0028844f $X=1.465 $Y=0.152 $X2=1.835 $Y2=1
cc_70 N_noxref_1_c_13_p N_Y_c_387_n 0.0142303f $X=1.55 $Y=0.755 $X2=1.835 $Y2=1
cc_71 N_noxref_1_c_21_p N_Y_c_387_n 0.0028844f $X=2.325 $Y=0.152 $X2=1.835 $Y2=1
cc_72 N_noxref_1_M1006_b N_Y_c_391_n 0.0437239f $X=-0.045 $Y=0 $X2=1.98
+ $Y2=2.365
cc_73 N_noxref_1_M1010_s N_Y_c_392_n 0.0100329f $X=2.27 $Y=0.575 $X2=2.695 $Y2=1
cc_74 N_noxref_1_c_21_p N_Y_c_392_n 0.0028844f $X=2.325 $Y=0.152 $X2=2.695 $Y2=1
cc_75 N_noxref_1_c_26_p N_Y_c_392_n 0.0142303f $X=2.41 $Y=0.755 $X2=2.695 $Y2=1
cc_76 N_noxref_1_c_32_p N_Y_c_392_n 0.0028844f $X=3.185 $Y=0.152 $X2=2.695 $Y2=1
cc_77 N_noxref_1_M1006_b N_Y_c_396_n 0.00409378f $X=-0.045 $Y=0 $X2=2.125 $Y2=1
cc_78 N_noxref_1_c_13_p N_Y_c_396_n 7.53951e-19 $X=1.55 $Y=0.755 $X2=2.125 $Y2=1
cc_79 N_noxref_1_c_21_p N_Y_c_396_n 0.00245319f $X=2.325 $Y=0.152 $X2=2.125
+ $Y2=1
cc_80 N_noxref_1_c_26_p N_Y_c_396_n 7.53951e-19 $X=2.41 $Y=0.755 $X2=2.125 $Y2=1
cc_81 N_noxref_1_M1006_b N_Y_c_400_n 0.00560779f $X=-0.045 $Y=0 $X2=2.125
+ $Y2=2.48
cc_82 N_noxref_1_M1006_b N_Y_c_401_n 0.00409378f $X=-0.045 $Y=0 $X2=2.84
+ $Y2=1.115
cc_83 N_noxref_1_c_26_p N_Y_c_401_n 7.53951e-19 $X=2.41 $Y=0.755 $X2=2.84
+ $Y2=1.115
cc_84 N_noxref_1_c_32_p N_Y_c_401_n 0.00245319f $X=3.185 $Y=0.152 $X2=2.84
+ $Y2=1.115
cc_85 N_noxref_1_c_38_p N_Y_c_401_n 0.00134236f $X=3.27 $Y=0.755 $X2=2.84
+ $Y2=1.115
cc_86 N_noxref_1_M1006_b N_Y_c_405_n 0.0625307f $X=-0.045 $Y=0 $X2=2.84
+ $Y2=2.365
cc_87 N_noxref_1_M1006_b GND 0.251858f $X=-0.045 $Y=0 $X2=0.34 $Y2=0.22
cc_88 N_noxref_1_c_2_p GND 0.0440059f $X=0.605 $Y=0.152 $X2=0.34 $Y2=0.22
cc_89 N_noxref_1_c_9_p GND 0.0435303f $X=1.465 $Y=0.152 $X2=0.34 $Y2=0.22
cc_90 N_noxref_1_c_21_p GND 0.042979f $X=2.325 $Y=0.152 $X2=0.34 $Y2=0.22
cc_91 N_noxref_1_c_32_p GND 0.0887744f $X=3.185 $Y=0.152 $X2=0.34 $Y2=0.22
cc_92 N_noxref_1_c_92_p GND 0.0189324f $X=0.69 $Y=0.152 $X2=0.34 $Y2=0.22
cc_93 N_noxref_1_c_93_p GND 0.0189324f $X=1.55 $Y=0.152 $X2=0.34 $Y2=0.22
cc_94 N_noxref_2_M1004_b N_A_M1004_g 0.0245629f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_95 N_noxref_2_c_95_p N_A_M1004_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_96 N_noxref_2_c_96_p N_A_M1004_g 0.00337744f $X=0.69 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_97 N_noxref_2_M1004_d N_A_c_159_n 0.00628533f $X=0.55 $Y=2.605 $X2=0.635
+ $Y2=2
cc_98 N_noxref_2_M1004_b N_A_c_159_n 0.00328912f $X=-0.045 $Y=2.425 $X2=0.635
+ $Y2=2
cc_99 N_noxref_2_c_96_p N_A_c_159_n 0.00264661f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2
cc_100 N_noxref_2_M1004_d A 0.00797576f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2.85
cc_101 N_noxref_2_c_96_p A 0.00510982f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2.85
cc_102 N_noxref_2_M1004_b N_A_27_115#_c_239_n 0.014249f $X=-0.045 $Y=2.425
+ $X2=0.905 $Y2=2.53
cc_103 N_noxref_2_c_96_p N_A_27_115#_c_239_n 0.00337744f $X=0.69 $Y=3.635
+ $X2=0.905 $Y2=2.53
cc_104 N_noxref_2_c_104_p N_A_27_115#_c_239_n 0.00606474f $X=1.465 $Y=4.287
+ $X2=0.905 $Y2=2.53
cc_105 N_noxref_2_M1004_b N_A_27_115#_c_242_n 0.0141063f $X=-0.045 $Y=2.425
+ $X2=1.335 $Y2=2.53
cc_106 N_noxref_2_c_96_p N_A_27_115#_c_242_n 3.67508e-19 $X=0.69 $Y=3.635
+ $X2=1.335 $Y2=2.53
cc_107 N_noxref_2_c_104_p N_A_27_115#_c_242_n 0.00610567f $X=1.465 $Y=4.287
+ $X2=1.335 $Y2=2.53
cc_108 N_noxref_2_c_108_p N_A_27_115#_c_242_n 0.0035715f $X=1.55 $Y=2.955
+ $X2=1.335 $Y2=2.53
cc_109 N_noxref_2_M1004_b N_A_27_115#_c_204_n 0.00647677f $X=-0.045 $Y=2.425
+ $X2=1.69 $Y2=2.455
cc_110 N_noxref_2_c_108_p N_A_27_115#_c_204_n 0.00364479f $X=1.55 $Y=2.955
+ $X2=1.69 $Y2=2.455
cc_111 N_noxref_2_M1004_b N_A_27_115#_c_205_n 0.0113915f $X=-0.045 $Y=2.425
+ $X2=1.41 $Y2=2.455
cc_112 N_noxref_2_M1004_b N_A_27_115#_c_249_n 0.0137901f $X=-0.045 $Y=2.425
+ $X2=1.765 $Y2=2.53
cc_113 N_noxref_2_c_108_p N_A_27_115#_c_249_n 0.00337744f $X=1.55 $Y=2.955
+ $X2=1.765 $Y2=2.53
cc_114 N_noxref_2_c_114_p N_A_27_115#_c_249_n 0.00606474f $X=2.325 $Y=4.287
+ $X2=1.765 $Y2=2.53
cc_115 N_noxref_2_M1004_b N_A_27_115#_c_210_n 0.00596183f $X=-0.045 $Y=2.425
+ $X2=2.12 $Y2=2.455
cc_116 N_noxref_2_M1004_b N_A_27_115#_c_253_n 0.0137901f $X=-0.045 $Y=2.425
+ $X2=2.195 $Y2=2.53
cc_117 N_noxref_2_c_114_p N_A_27_115#_c_253_n 0.00606474f $X=2.325 $Y=4.287
+ $X2=2.195 $Y2=2.53
cc_118 N_noxref_2_c_118_p N_A_27_115#_c_253_n 0.00337744f $X=2.41 $Y=2.955
+ $X2=2.195 $Y2=2.53
cc_119 N_noxref_2_M1004_b N_A_27_115#_c_216_n 0.00647677f $X=-0.045 $Y=2.425
+ $X2=2.55 $Y2=2.455
cc_120 N_noxref_2_c_118_p N_A_27_115#_c_216_n 0.00364479f $X=2.41 $Y=2.955
+ $X2=2.55 $Y2=2.455
cc_121 N_noxref_2_M1004_b N_A_27_115#_c_258_n 0.0137901f $X=-0.045 $Y=2.425
+ $X2=2.625 $Y2=2.53
cc_122 N_noxref_2_c_118_p N_A_27_115#_c_258_n 0.00337744f $X=2.41 $Y=2.955
+ $X2=2.625 $Y2=2.53
cc_123 N_noxref_2_c_123_p N_A_27_115#_c_258_n 0.00606474f $X=3.185 $Y=4.287
+ $X2=2.625 $Y2=2.53
cc_124 N_noxref_2_M1004_b N_A_27_115#_c_222_n 0.0134369f $X=-0.045 $Y=2.425
+ $X2=2.98 $Y2=2.455
cc_125 N_noxref_2_M1004_b N_A_27_115#_c_262_n 0.0166569f $X=-0.045 $Y=2.425
+ $X2=3.055 $Y2=2.53
cc_126 N_noxref_2_c_123_p N_A_27_115#_c_262_n 0.00606474f $X=3.185 $Y=4.287
+ $X2=3.055 $Y2=2.53
cc_127 N_noxref_2_c_127_p N_A_27_115#_c_262_n 0.00636672f $X=3.27 $Y=2.955
+ $X2=3.055 $Y2=2.53
cc_128 N_noxref_2_M1004_b N_A_27_115#_c_227_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=1.765 $Y2=2.455
cc_129 N_noxref_2_M1004_b N_A_27_115#_c_229_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=2.195 $Y2=2.455
cc_130 N_noxref_2_M1004_b N_A_27_115#_c_231_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=2.625 $Y2=2.455
cc_131 N_noxref_2_M1004_b N_A_27_115#_c_234_n 0.00996008f $X=-0.045 $Y=2.425
+ $X2=0.26 $Y2=2.955
cc_132 N_noxref_2_c_95_p N_A_27_115#_c_234_n 0.00736239f $X=0.605 $Y=4.287
+ $X2=0.26 $Y2=2.955
cc_133 N_noxref_2_M1004_b N_Y_c_406_n 0.00290209f $X=-0.045 $Y=2.425 $X2=1.12
+ $Y2=2.48
cc_134 N_noxref_2_c_104_p N_Y_c_406_n 0.00734006f $X=1.465 $Y=4.287 $X2=1.12
+ $Y2=2.48
cc_135 N_noxref_2_M1004_b N_Y_c_408_n 0.00337919f $X=-0.045 $Y=2.425 $X2=1.98
+ $Y2=2.48
cc_136 N_noxref_2_c_114_p N_Y_c_408_n 0.00754406f $X=2.325 $Y=4.287 $X2=1.98
+ $Y2=2.48
cc_137 N_noxref_2_M1004_b N_Y_c_410_n 0.00337919f $X=-0.045 $Y=2.425 $X2=2.84
+ $Y2=2.48
cc_138 N_noxref_2_c_123_p N_Y_c_410_n 0.00746708f $X=3.185 $Y=4.287 $X2=2.84
+ $Y2=2.48
cc_139 N_noxref_2_M1004_b N_Y_c_385_n 0.00409378f $X=-0.045 $Y=2.425 $X2=1.12
+ $Y2=2.365
cc_140 N_noxref_2_M1004_b N_Y_c_413_n 0.00520877f $X=-0.045 $Y=2.425 $X2=1.835
+ $Y2=2.48
cc_141 N_noxref_2_c_108_p N_Y_c_413_n 0.0090257f $X=1.55 $Y=2.955 $X2=1.835
+ $Y2=2.48
cc_142 N_noxref_2_M1004_b N_Y_c_415_n 0.00520877f $X=-0.045 $Y=2.425 $X2=2.695
+ $Y2=2.48
cc_143 N_noxref_2_c_118_p N_Y_c_415_n 0.0090257f $X=2.41 $Y=2.955 $X2=2.695
+ $Y2=2.48
cc_144 N_noxref_2_M1004_b N_Y_c_400_n 0.00409378f $X=-0.045 $Y=2.425 $X2=2.125
+ $Y2=2.48
cc_145 N_noxref_2_M1004_b N_Y_c_405_n 0.00409378f $X=-0.045 $Y=2.425 $X2=2.84
+ $Y2=2.365
cc_146 N_noxref_2_M1004_b VDD 0.269451f $X=-0.045 $Y=2.425 $X2=0.34 $Y2=4.22
cc_147 N_noxref_2_c_95_p VDD 0.0439891f $X=0.605 $Y=4.287 $X2=0.34 $Y2=4.22
cc_148 N_noxref_2_c_104_p VDD 0.0435303f $X=1.465 $Y=4.287 $X2=0.34 $Y2=4.22
cc_149 N_noxref_2_c_114_p VDD 0.042979f $X=2.325 $Y=4.287 $X2=0.34 $Y2=4.22
cc_150 N_noxref_2_c_123_p VDD 0.0887744f $X=3.185 $Y=4.287 $X2=0.34 $Y2=4.22
cc_151 N_noxref_2_c_151_p VDD 0.0189324f $X=0.69 $Y=4.287 $X2=0.34 $Y2=4.22
cc_152 N_noxref_2_c_152_p VDD 0.0189324f $X=1.55 $Y=4.287 $X2=0.34 $Y2=4.22
cc_153 N_noxref_2_c_153_p VDD 0.0189324f $X=2.38 $Y=4.22 $X2=0.34 $Y2=4.22
cc_154 A N_A_27_115#_M1004_s 0.00410657f $X=0.635 $Y=2.85 $X2=0.135 $Y2=2.605
cc_155 N_A_M1006_g N_A_27_115#_M1000_g 0.0342527f $X=0.475 $Y=0.835 $X2=0.905
+ $Y2=0.835
cc_156 A N_A_27_115#_c_239_n 0.00419145f $X=0.635 $Y=2.85 $X2=0.905 $Y2=2.53
cc_157 N_A_M1006_g N_A_27_115#_c_197_n 0.00260138f $X=0.475 $Y=0.835 $X2=1.18
+ $Y2=2.38
cc_158 N_A_M1004_g N_A_27_115#_c_197_n 0.00209773f $X=0.475 $Y=3.235 $X2=1.18
+ $Y2=2.38
cc_159 N_A_c_158_n N_A_27_115#_c_197_n 0.0139096f $X=0.635 $Y=2 $X2=1.18
+ $Y2=2.38
cc_160 N_A_c_159_n N_A_27_115#_c_197_n 0.00361737f $X=0.635 $Y=2 $X2=1.18
+ $Y2=2.38
cc_161 N_A_M1004_g N_A_27_115#_c_205_n 0.0485392f $X=0.475 $Y=3.235 $X2=1.41
+ $Y2=2.455
cc_162 N_A_c_159_n N_A_27_115#_c_205_n 0.00477416f $X=0.635 $Y=2 $X2=1.41
+ $Y2=2.455
cc_163 N_A_M1006_g N_A_27_115#_c_232_n 0.0124465f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.755
cc_164 N_A_M1006_g N_A_27_115#_c_234_n 0.0330322f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=2.955
cc_165 N_A_c_159_n N_A_27_115#_c_234_n 0.0548951f $X=0.635 $Y=2 $X2=0.26
+ $Y2=2.955
cc_166 A N_A_27_115#_c_234_n 0.0155137f $X=0.635 $Y=2.85 $X2=0.26 $Y2=2.955
cc_167 N_A_M1006_g N_A_27_115#_c_235_n 0.0207696f $X=0.475 $Y=0.835 $X2=0.88
+ $Y2=1.455
cc_168 N_A_c_158_n N_A_27_115#_c_235_n 0.00273049f $X=0.635 $Y=2 $X2=0.88
+ $Y2=1.455
cc_169 N_A_c_159_n N_A_27_115#_c_235_n 0.00886797f $X=0.635 $Y=2 $X2=0.88
+ $Y2=1.455
cc_170 N_A_M1006_g N_A_27_115#_c_238_n 6.59135e-19 $X=0.475 $Y=0.835 $X2=0.965
+ $Y2=1.455
cc_171 N_A_c_159_n N_Y_c_406_n 0.0135622f $X=0.635 $Y=2 $X2=1.12 $Y2=2.48
cc_172 A N_Y_c_406_n 0.00731851f $X=0.635 $Y=2.85 $X2=1.12 $Y2=2.48
cc_173 N_A_M1006_g N_Y_c_381_n 8.01483e-19 $X=0.475 $Y=0.835 $X2=1.12 $Y2=1.115
cc_174 N_A_c_159_n N_Y_c_385_n 0.00677552f $X=0.635 $Y=2 $X2=1.12 $Y2=2.365
cc_175 N_A_M1006_g Y 0.00310306f $X=0.475 $Y=0.835 $X2=1.055 $Y2=1.79
cc_176 N_A_c_158_n Y 0.00441844f $X=0.635 $Y=2 $X2=1.055 $Y2=1.79
cc_177 N_A_c_159_n Y 0.0200396f $X=0.635 $Y=2 $X2=1.055 $Y2=1.79
cc_178 N_A_M1006_g GND 0.00468827f $X=0.475 $Y=0.835 $X2=0.34 $Y2=0.22
cc_179 N_A_M1004_g VDD 0.00468827f $X=0.475 $Y=3.235 $X2=0.34 $Y2=4.22
cc_180 N_A_27_115#_M1000_g N_Y_c_371_n 0.00182852f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_181 N_A_27_115#_M1001_g N_Y_c_371_n 0.00182852f $X=1.335 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_182 N_A_27_115#_c_203_n N_Y_c_371_n 0.00296072f $X=1.41 $Y=1.365 $X2=1.12
+ $Y2=0.755
cc_183 N_A_27_115#_c_238_n N_Y_c_371_n 7.29965e-19 $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=0.755
cc_184 N_A_27_115#_c_239_n N_Y_c_406_n 0.00138273f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_185 N_A_27_115#_c_242_n N_Y_c_406_n 0.00233646f $X=1.335 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_186 N_A_27_115#_c_205_n N_Y_c_406_n 0.0126676f $X=1.41 $Y=2.455 $X2=1.12
+ $Y2=2.48
cc_187 N_A_27_115#_M1008_g N_Y_c_374_n 0.00182852f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=0.755
cc_188 N_A_27_115#_c_209_n N_Y_c_374_n 0.00274041f $X=2.12 $Y=1.365 $X2=1.98
+ $Y2=0.755
cc_189 N_A_27_115#_M1010_g N_Y_c_374_n 0.00182852f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=0.755
cc_190 N_A_27_115#_c_249_n N_Y_c_408_n 0.00233646f $X=1.765 $Y=2.53 $X2=1.98
+ $Y2=2.48
cc_191 N_A_27_115#_c_210_n N_Y_c_408_n 0.0138847f $X=2.12 $Y=2.455 $X2=1.98
+ $Y2=2.48
cc_192 N_A_27_115#_c_253_n N_Y_c_408_n 0.00233646f $X=2.195 $Y=2.53 $X2=1.98
+ $Y2=2.48
cc_193 N_A_27_115#_M1011_g N_Y_c_378_n 0.00182852f $X=2.625 $Y=0.835 $X2=2.84
+ $Y2=0.755
cc_194 N_A_27_115#_c_221_n N_Y_c_378_n 0.00274041f $X=2.98 $Y=1.365 $X2=2.84
+ $Y2=0.755
cc_195 N_A_27_115#_M1013_g N_Y_c_378_n 0.00182852f $X=3.055 $Y=0.835 $X2=2.84
+ $Y2=0.755
cc_196 N_A_27_115#_c_258_n N_Y_c_410_n 0.00233646f $X=2.625 $Y=2.53 $X2=2.84
+ $Y2=2.48
cc_197 N_A_27_115#_c_222_n N_Y_c_410_n 0.013404f $X=2.98 $Y=2.455 $X2=2.84
+ $Y2=2.48
cc_198 N_A_27_115#_c_262_n N_Y_c_410_n 0.00233646f $X=3.055 $Y=2.53 $X2=2.84
+ $Y2=2.48
cc_199 N_A_27_115#_M1000_g N_Y_c_381_n 0.00480694f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=1.115
cc_200 N_A_27_115#_M1001_g N_Y_c_381_n 0.00201073f $X=1.335 $Y=0.835 $X2=1.12
+ $Y2=1.115
cc_201 N_A_27_115#_c_238_n N_Y_c_381_n 0.00278861f $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=1.115
cc_202 N_A_27_115#_c_239_n N_Y_c_385_n 0.00120715f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.365
cc_203 N_A_27_115#_c_197_n N_Y_c_385_n 0.00215118f $X=1.18 $Y=2.38 $X2=1.12
+ $Y2=2.365
cc_204 N_A_27_115#_c_242_n N_Y_c_385_n 0.00113627f $X=1.335 $Y=2.53 $X2=1.12
+ $Y2=2.365
cc_205 N_A_27_115#_c_205_n N_Y_c_385_n 0.00372325f $X=1.41 $Y=2.455 $X2=1.12
+ $Y2=2.365
cc_206 N_A_27_115#_M1000_g Y 0.00251111f $X=0.905 $Y=0.835 $X2=1.055 $Y2=1.79
cc_207 N_A_27_115#_c_197_n Y 0.0314621f $X=1.18 $Y=2.38 $X2=1.055 $Y2=1.79
cc_208 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=0.835 $X2=1.055 $Y2=1.79
cc_209 N_A_27_115#_c_203_n Y 0.0166018f $X=1.41 $Y=1.365 $X2=1.055 $Y2=1.79
cc_210 N_A_27_115#_c_235_n Y 8.73078e-19 $X=0.88 $Y=1.455 $X2=1.055 $Y2=1.79
cc_211 N_A_27_115#_c_238_n Y 0.0121742f $X=0.965 $Y=1.455 $X2=1.055 $Y2=1.79
cc_212 N_A_27_115#_M1001_g N_Y_c_387_n 0.00908832f $X=1.335 $Y=0.835 $X2=1.835
+ $Y2=1
cc_213 N_A_27_115#_c_201_n N_Y_c_387_n 0.00213861f $X=1.69 $Y=1.365 $X2=1.835
+ $Y2=1
cc_214 N_A_27_115#_M1008_g N_Y_c_387_n 0.00873177f $X=1.765 $Y=0.835 $X2=1.835
+ $Y2=1
cc_215 N_A_27_115#_c_242_n N_Y_c_413_n 0.00639369f $X=1.335 $Y=2.53 $X2=1.835
+ $Y2=2.48
cc_216 N_A_27_115#_c_204_n N_Y_c_413_n 0.0125005f $X=1.69 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_217 N_A_27_115#_c_205_n N_Y_c_413_n 0.00627763f $X=1.41 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_218 N_A_27_115#_c_249_n N_Y_c_413_n 0.00639369f $X=1.765 $Y=2.53 $X2=1.835
+ $Y2=2.48
cc_219 N_A_27_115#_c_227_n N_Y_c_413_n 0.00580646f $X=1.765 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_220 N_A_27_115#_c_203_n N_Y_c_391_n 0.013329f $X=1.41 $Y=1.365 $X2=1.98
+ $Y2=2.365
cc_221 N_A_27_115#_M1008_g N_Y_c_391_n 0.00251111f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=2.365
cc_222 N_A_27_115#_c_209_n N_Y_c_391_n 0.0178059f $X=2.12 $Y=1.365 $X2=1.98
+ $Y2=2.365
cc_223 N_A_27_115#_M1010_g N_Y_c_391_n 0.00251111f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=2.365
cc_224 N_A_27_115#_c_220_n N_Y_c_391_n 0.0137936f $X=2.625 $Y=2.38 $X2=1.98
+ $Y2=2.365
cc_225 N_A_27_115#_M1010_g N_Y_c_392_n 0.00873177f $X=2.195 $Y=0.835 $X2=2.695
+ $Y2=1
cc_226 N_A_27_115#_c_214_n N_Y_c_392_n 0.00213861f $X=2.55 $Y=1.365 $X2=2.695
+ $Y2=1
cc_227 N_A_27_115#_M1011_g N_Y_c_392_n 0.00938169f $X=2.625 $Y=0.835 $X2=2.695
+ $Y2=1
cc_228 N_A_27_115#_M1008_g N_Y_c_396_n 0.00198614f $X=1.765 $Y=0.835 $X2=2.125
+ $Y2=1
cc_229 N_A_27_115#_M1010_g N_Y_c_396_n 0.00198614f $X=2.195 $Y=0.835 $X2=2.125
+ $Y2=1
cc_230 N_A_27_115#_c_253_n N_Y_c_415_n 0.00639369f $X=2.195 $Y=2.53 $X2=2.695
+ $Y2=2.48
cc_231 N_A_27_115#_c_216_n N_Y_c_415_n 0.0130313f $X=2.55 $Y=2.455 $X2=2.695
+ $Y2=2.48
cc_232 N_A_27_115#_c_258_n N_Y_c_415_n 0.00639369f $X=2.625 $Y=2.53 $X2=2.695
+ $Y2=2.48
cc_233 N_A_27_115#_c_229_n N_Y_c_415_n 0.00580646f $X=2.195 $Y=2.455 $X2=2.695
+ $Y2=2.48
cc_234 N_A_27_115#_c_231_n N_Y_c_415_n 0.00666531f $X=2.625 $Y=2.455 $X2=2.695
+ $Y2=2.48
cc_235 N_A_27_115#_c_249_n N_Y_c_400_n 0.00113627f $X=1.765 $Y=2.53 $X2=2.125
+ $Y2=2.48
cc_236 N_A_27_115#_c_210_n N_Y_c_400_n 0.00364679f $X=2.12 $Y=2.455 $X2=2.125
+ $Y2=2.48
cc_237 N_A_27_115#_c_253_n N_Y_c_400_n 0.00113627f $X=2.195 $Y=2.53 $X2=2.125
+ $Y2=2.48
cc_238 N_A_27_115#_c_227_n N_Y_c_400_n 6.99501e-19 $X=1.765 $Y=2.455 $X2=2.125
+ $Y2=2.48
cc_239 N_A_27_115#_c_229_n N_Y_c_400_n 6.99501e-19 $X=2.195 $Y=2.455 $X2=2.125
+ $Y2=2.48
cc_240 N_A_27_115#_M1011_g N_Y_c_401_n 0.00201073f $X=2.625 $Y=0.835 $X2=2.84
+ $Y2=1.115
cc_241 N_A_27_115#_M1013_g N_Y_c_401_n 0.00878256f $X=3.055 $Y=0.835 $X2=2.84
+ $Y2=1.115
cc_242 N_A_27_115#_M1011_g N_Y_c_405_n 0.00251111f $X=2.625 $Y=0.835 $X2=2.84
+ $Y2=2.365
cc_243 N_A_27_115#_c_220_n N_Y_c_405_n 0.0185925f $X=2.625 $Y=2.38 $X2=2.84
+ $Y2=2.365
cc_244 N_A_27_115#_c_258_n N_Y_c_405_n 0.00113627f $X=2.625 $Y=2.53 $X2=2.84
+ $Y2=2.365
cc_245 N_A_27_115#_c_221_n N_Y_c_405_n 0.0170354f $X=2.98 $Y=1.365 $X2=2.84
+ $Y2=2.365
cc_246 N_A_27_115#_c_222_n N_Y_c_405_n 0.00966211f $X=2.98 $Y=2.455 $X2=2.84
+ $Y2=2.365
cc_247 N_A_27_115#_M1013_g N_Y_c_405_n 0.00251111f $X=3.055 $Y=0.835 $X2=2.84
+ $Y2=2.365
cc_248 N_A_27_115#_c_262_n N_Y_c_405_n 0.0031083f $X=3.055 $Y=2.53 $X2=2.84
+ $Y2=2.365
cc_249 N_A_27_115#_c_231_n N_Y_c_405_n 6.59375e-19 $X=2.625 $Y=2.455 $X2=2.84
+ $Y2=2.365
cc_250 N_A_27_115#_M1000_g GND 0.00468827f $X=0.905 $Y=0.835 $X2=0.34 $Y2=0.22
cc_251 N_A_27_115#_M1001_g GND 0.00468827f $X=1.335 $Y=0.835 $X2=0.34 $Y2=0.22
cc_252 N_A_27_115#_M1008_g GND 0.00468827f $X=1.765 $Y=0.835 $X2=0.34 $Y2=0.22
cc_253 N_A_27_115#_M1010_g GND 0.00468827f $X=2.195 $Y=0.835 $X2=0.34 $Y2=0.22
cc_254 N_A_27_115#_M1011_g GND 0.00468827f $X=2.625 $Y=0.835 $X2=0.34 $Y2=0.22
cc_255 N_A_27_115#_M1013_g GND 0.00468827f $X=3.055 $Y=0.835 $X2=0.34 $Y2=0.22
cc_256 N_A_27_115#_c_232_n GND 0.00476261f $X=0.26 $Y=0.755 $X2=0.34 $Y2=0.22
cc_257 N_A_27_115#_c_239_n VDD 0.00468827f $X=0.905 $Y=2.53 $X2=0.34 $Y2=4.22
cc_258 N_A_27_115#_c_242_n VDD 0.00470215f $X=1.335 $Y=2.53 $X2=0.34 $Y2=4.22
cc_259 N_A_27_115#_c_249_n VDD 0.00468827f $X=1.765 $Y=2.53 $X2=0.34 $Y2=4.22
cc_260 N_A_27_115#_c_253_n VDD 0.00468827f $X=2.195 $Y=2.53 $X2=0.34 $Y2=4.22
cc_261 N_A_27_115#_c_258_n VDD 0.00468827f $X=2.625 $Y=2.53 $X2=0.34 $Y2=4.22
cc_262 N_A_27_115#_c_262_n VDD 0.00468827f $X=3.055 $Y=2.53 $X2=0.34 $Y2=4.22
cc_263 N_A_27_115#_c_234_n VDD 0.00476261f $X=0.26 $Y=2.955 $X2=0.34 $Y2=4.22
cc_264 N_Y_c_371_n GND 0.0047139f $X=1.12 $Y=0.755 $X2=0.34 $Y2=0.22
cc_265 N_Y_c_374_n GND 0.0047139f $X=1.98 $Y=0.755 $X2=0.34 $Y2=0.22
cc_266 N_Y_c_378_n GND 0.0047139f $X=2.84 $Y=0.755 $X2=0.34 $Y2=0.22
cc_267 N_Y_c_406_n VDD 0.00475776f $X=1.12 $Y=2.48 $X2=0.34 $Y2=4.22
cc_268 N_Y_c_408_n VDD 0.00475776f $X=1.98 $Y=2.48 $X2=0.34 $Y2=4.22
cc_269 N_Y_c_410_n VDD 0.00475776f $X=2.84 $Y=2.48 $X2=0.34 $Y2=4.22
