* File: sky130_osu_sc_15T_ms__aoi22_l.pex.spice
* Created: Fri Nov 12 14:41:13 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%GND 1 2 27 31 33 44 56 58
c45 27 0 6.36774e-20 $X=-0.045 $Y=0
r46 56 58 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r47 42 52 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.152
r48 42 44 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.74
r49 33 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=0.152
+ $X2=1.91 $Y2=0.152
r50 29 31 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r51 27 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r52 27 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r53 27 29 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r54 27 34 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r55 27 33 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.825 $Y2=0.152
r56 27 34 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r57 2 44 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.77
+ $Y=0.575 $X2=1.91 $Y2=0.74
r58 1 31 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%VDD 1 17 19 26 34 39 43
r31 39 43 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.7 $Y2=5.397
r32 34 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=5.36 $X2=1.7
+ $Y2=5.36
r33 32 34 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=5.397
+ $X2=1.7 $Y2=5.397
r34 30 37 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r35 30 32 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r36 26 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=3.98
+ $X2=0.69 $Y2=4.66
r37 24 37 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r38 24 29 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.66
r39 21 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r40 19 37 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r41 19 21 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r42 17 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r43 17 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r44 17 21 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r45 1 29 400 $w=1.7e-07 $l=1.90371e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.66
r46 1 26 400 $w=1.7e-07 $l=1.223e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.98
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%A0 2 3 5 8 12 18 21 27
c35 8 0 6.36774e-20 $X=0.475 $Y=3.825
r36 24 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=3.07
+ $X2=0.385 $Y2=3.07
r37 21 24 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.385 $Y=2.505
+ $X2=0.385 $Y2=3.07
r38 17 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.505 $X2=0.385 $Y2=2.505
r39 17 18 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.505
+ $X2=0.475 $Y2=2.505
r40 14 17 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.505
+ $X2=0.385 $Y2=2.505
r41 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.51
+ $X2=0.475 $Y2=1.51
r42 6 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.64
+ $X2=0.475 $Y2=2.505
r43 6 8 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.475 $Y=2.64
+ $X2=0.475 $Y2=3.825
r44 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.43 $X2=0.475
+ $Y2=1.51
r45 3 5 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.475 $Y=1.43
+ $X2=0.475 $Y2=0.945
r46 2 14 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.37
+ $X2=0.295 $Y2=2.505
r47 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.59 $X2=0.295
+ $Y2=1.51
r48 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.59
+ $X2=0.295 $Y2=2.37
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%A1 3 5 7 12 18
r44 15 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.7
+ $X2=0.725 $Y2=2.7
r45 12 15 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.725 $Y=1.995
+ $X2=0.725 $Y2=2.7
r46 10 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.995 $X2=0.725 $Y2=1.995
r47 5 10 63.0864 $w=2.95e-07 $l=3.7229e-07 $layer=POLY_cond $X=0.905 $Y=2.31
+ $X2=0.78 $Y2=1.995
r48 5 7 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=0.905 $Y=2.31
+ $X2=0.905 $Y2=3.825
r49 1 10 38.578 $w=2.95e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.835 $Y=1.83
+ $X2=0.78 $Y2=1.995
r50 1 3 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=0.835 $Y=1.83
+ $X2=0.835 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%B0 3 7 10 15 17 21
c43 3 0 1.94783e-19 $X=1.335 $Y=0.945
r44 17 19 3.63576 $w=3.02e-07 $l=9e-08 $layer=LI1_cond $X=1.165 $Y=1.64
+ $X2=1.255 $Y2=1.64
r45 15 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.33
+ $X2=1.165 $Y2=2.33
r46 13 17 4.10007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=1.805
+ $X2=1.165 $Y2=1.64
r47 13 15 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.165 $Y=1.805
+ $X2=1.165 $Y2=2.33
r48 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.64 $X2=1.255 $Y2=1.64
r49 10 12 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.64
+ $X2=1.265 $Y2=1.805
r50 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.64
+ $X2=1.265 $Y2=1.475
r51 7 12 1035.79 $w=1.5e-07 $l=2.02e-06 $layer=POLY_cond $X=1.335 $Y=3.825
+ $X2=1.335 $Y2=1.805
r52 3 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=0.945
+ $X2=1.335 $Y2=1.475
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%B1 3 7 10 14 19
r27 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.935 $Y=1.965
+ $X2=1.935 $Y2=1.965
r28 12 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.965 $X2=1.935 $Y2=1.965
r29 10 12 26.0127 $w=3.15e-07 $l=1.7e-07 $layer=POLY_cond $X=1.765 $Y=1.945
+ $X2=1.935 $Y2=1.945
r30 9 10 10.7111 $w=3.15e-07 $l=7e-08 $layer=POLY_cond $X=1.695 $Y=1.945
+ $X2=1.765 $Y2=1.945
r31 5 10 20.1192 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.765 $Y=2.13
+ $X2=1.765 $Y2=1.945
r32 5 7 869.138 $w=1.5e-07 $l=1.695e-06 $layer=POLY_cond $X=1.765 $Y=2.13
+ $X2=1.765 $Y2=3.825
r33 1 9 20.1192 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.695 $Y=1.76
+ $X2=1.695 $Y2=1.945
r34 1 3 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.695 $Y=1.76
+ $X2=1.695 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%A_27_565# 1 2 3 13 15 17 23 24
r25 27 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.98 $Y=3.64
+ $X2=1.98 $Y2=4.66
r26 25 30 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.98 $Y=4.75 $X2=1.98
+ $Y2=4.66
r27 23 25 6.81835 $w=1.75e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.895 $Y=4.837
+ $X2=1.98 $Y2=4.75
r28 23 24 43.7299 $w=1.73e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=4.837
+ $X2=1.205 $Y2=4.837
r29 20 24 6.81835 $w=1.75e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.12 $Y=4.75
+ $X2=1.205 $Y2=4.837
r30 20 22 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.12 $Y=4.75 $X2=1.12
+ $Y2=4.66
r31 19 34 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=3.645
+ $X2=1.12 $Y2=3.56
r32 19 22 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=1.12 $Y=3.645
+ $X2=1.12 $Y2=4.66
r33 18 32 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=3.56
+ $X2=0.26 $Y2=3.56
r34 17 34 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=3.56
+ $X2=1.12 $Y2=3.56
r35 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.56
+ $X2=0.345 $Y2=3.56
r36 13 32 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=3.645
+ $X2=0.26 $Y2=3.56
r37 13 15 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=0.26 $Y=3.645
+ $X2=0.26 $Y2=4.66
r38 3 30 300 $w=1.7e-07 $l=1.90371e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.66
r39 3 27 300 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.64
r40 2 22 300 $w=1.7e-07 $l=1.90371e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.66
r41 2 34 300 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.64
r42 1 15 300 $w=1.7e-07 $l=1.89647e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.66
r43 1 32 300 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.64
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AOI22_L%Y 1 3 10 17 23 27 28 32 38
c39 32 0 5.84789e-20 $X=1.605 $Y=1.44
c40 28 0 1.94783e-19 $X=1.23 $Y=1.22
r41 38 39 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.595 $Y=1.59
+ $X2=1.595 $Y2=1.475
r42 32 39 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.605 $Y=1.44
+ $X2=1.605 $Y2=1.475
r43 29 32 0.129989 $w=1.7e-07 $l=1.35e-07 $layer=MET1_cond $X=1.605 $Y=1.305
+ $X2=1.605 $Y2=1.44
r44 28 35 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.23 $Y=1.22
+ $X2=1.085 $Y2=1.22
r45 27 29 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.52 $Y=1.22
+ $X2=1.605 $Y2=1.305
r46 27 28 0.279236 $w=1.7e-07 $l=2.9e-07 $layer=MET1_cond $X=1.52 $Y=1.22
+ $X2=1.23 $Y2=1.22
r47 25 26 9.11234 $w=2.13e-07 $l=1.7e-07 $layer=LI1_cond $X=1.572 $Y=2.9
+ $X2=1.572 $Y2=3.07
r48 23 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.595 $Y=1.59
+ $X2=1.595 $Y2=1.59
r49 23 25 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.595 $Y=1.59
+ $X2=1.595 $Y2=2.9
r50 17 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=3.64
+ $X2=1.55 $Y2=4.32
r51 17 26 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.55 $Y=3.64
+ $X2=1.55 $Y2=3.07
r52 13 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=1.22
+ $X2=1.085 $Y2=1.22
r53 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.085 $Y=0.74
+ $X2=1.085 $Y2=1.22
r54 3 19 400 $w=1.7e-07 $l=1.56343e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.32
r55 3 17 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.64
r56 1 10 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.085 $Y2=0.74
.ends

