* File: sky130_osu_sc_18T_ls__oai22_l.spice
* Created: Thu Oct 29 17:37:46 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ls__oai22_l.pex.spice"
.subckt sky130_osu_sc_18T_ls__oai22_l  GND VDD A0 A1 B0 B1 Y
* 
* Y	Y
* B1	B1
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A0_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1000 N_A_27_115#_M1000_d N_A1_M1000_g N_GND_M1004_d N_GND_M1004_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_B0_M1001_g N_A_27_115#_M1000_d N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_115#_M1007_d N_B1_M1007_g N_Y_M1001_d N_GND_M1004_b NSHORT L=0.15
+ W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 A_110_617# N_A0_M1003_g N_VDD_M1003_s N_VDD_M1003_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001.4 A=0.45 P=6.3 MULT=1
MM1002 N_Y_M1002_d N_A1_M1002_g A_110_617# N_VDD_M1003_b PHIGHVT L=0.15 W=3
+ AD=0.525 AS=0.315 PD=3.35 PS=3.21 NRD=2.2852 NRS=3.2702 M=1 R=20 SA=75000.5
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1005 A_282_617# N_B0_M1005_g N_Y_M1002_d N_VDD_M1003_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.525 PD=3.21 PS=3.35 NRD=3.2702 NRS=2.2852 M=1 R=20 SA=75001
+ SB=75000.5 A=0.45 P=6.3 MULT=1
MM1006 N_VDD_M1006_d N_B1_M1006_g A_282_617# N_VDD_M1003_b PHIGHVT L=0.15 W=3
+ AD=0.795 AS=0.315 PD=6.53 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.4
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX8_noxref N_GND_M1004_b N_VDD_M1003_b NWDIODE A=8.949 P=12.31
pX9_noxref noxref_11 A0 A0 PROBETYPE=1
pX10_noxref noxref_12 A1 A1 PROBETYPE=1
pX11_noxref noxref_13 B0 B0 PROBETYPE=1
pX12_noxref noxref_14 Y Y PROBETYPE=1
pX13_noxref noxref_15 B1 B1 PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__oai22_l.pxi.spice"
*
.ends
*
*
