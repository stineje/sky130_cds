* File: sky130_osu_sc_15T_hs__buf_8.pxi.spice
* Created: Fri Nov 12 14:28:34 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__BUF_8%GND N_GND_M1007_d N_GND_M1004_s N_GND_M1011_s
+ N_GND_M1013_s N_GND_M1015_s N_GND_M1007_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p
+ N_GND_c_15_p N_GND_c_24_p N_GND_c_30_p N_GND_c_37_p N_GND_c_44_p N_GND_c_51_p
+ N_GND_c_57_p GND N_GND_c_4_p PM_SKY130_OSU_SC_15T_HS__BUF_8%GND
x_PM_SKY130_OSU_SC_15T_HS__BUF_8%VDD N_VDD_M1009_d N_VDD_M1001_s N_VDD_M1005_s
+ N_VDD_M1010_s N_VDD_M1017_s N_VDD_M1009_b N_VDD_c_124_p N_VDD_c_125_p
+ N_VDD_c_134_p N_VDD_c_139_p N_VDD_c_146_p N_VDD_c_151_p N_VDD_c_157_p
+ N_VDD_c_162_p N_VDD_c_168_p N_VDD_c_173_p VDD N_VDD_c_126_p
+ PM_SKY130_OSU_SC_15T_HS__BUF_8%VDD
x_PM_SKY130_OSU_SC_15T_HS__BUF_8%A N_A_M1007_g N_A_M1009_g N_A_c_210_n
+ N_A_c_211_n A PM_SKY130_OSU_SC_15T_HS__BUF_8%A
x_PM_SKY130_OSU_SC_15T_HS__BUF_8%A_27_115# N_A_27_115#_M1007_s
+ N_A_27_115#_M1009_s N_A_27_115#_M1002_g N_A_27_115#_c_314_n
+ N_A_27_115#_M1000_g N_A_27_115#_c_249_n N_A_27_115#_M1004_g
+ N_A_27_115#_c_318_n N_A_27_115#_M1001_g N_A_27_115#_c_254_n
+ N_A_27_115#_c_256_n N_A_27_115#_c_257_n N_A_27_115#_c_258_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_326_n N_A_27_115#_M1003_g
+ N_A_27_115#_c_263_n N_A_27_115#_c_264_n N_A_27_115#_M1011_g
+ N_A_27_115#_c_331_n N_A_27_115#_M1005_g N_A_27_115#_c_269_n
+ N_A_27_115#_c_271_n N_A_27_115#_M1012_g N_A_27_115#_c_276_n
+ N_A_27_115#_c_337_n N_A_27_115#_M1006_g N_A_27_115#_c_277_n
+ N_A_27_115#_c_278_n N_A_27_115#_M1013_g N_A_27_115#_c_342_n
+ N_A_27_115#_M1010_g N_A_27_115#_c_283_n N_A_27_115#_c_285_n
+ N_A_27_115#_M1014_g N_A_27_115#_c_348_n N_A_27_115#_M1016_g
+ N_A_27_115#_c_290_n N_A_27_115#_c_291_n N_A_27_115#_M1015_g
+ N_A_27_115#_c_353_n N_A_27_115#_M1017_g N_A_27_115#_c_296_n
+ N_A_27_115#_c_297_n N_A_27_115#_c_298_n N_A_27_115#_c_299_n
+ N_A_27_115#_c_300_n N_A_27_115#_c_301_n N_A_27_115#_c_302_n
+ N_A_27_115#_c_303_n N_A_27_115#_c_304_n N_A_27_115#_c_305_n
+ N_A_27_115#_c_306_n N_A_27_115#_c_309_n N_A_27_115#_c_310_n
+ N_A_27_115#_c_312_n N_A_27_115#_c_313_n
+ PM_SKY130_OSU_SC_15T_HS__BUF_8%A_27_115#
x_PM_SKY130_OSU_SC_15T_HS__BUF_8%Y N_Y_M1002_d N_Y_M1008_d N_Y_M1012_d
+ N_Y_M1014_d N_Y_M1000_d N_Y_M1003_d N_Y_M1006_d N_Y_M1016_d N_Y_c_477_n
+ N_Y_c_523_n N_Y_c_481_n N_Y_c_526_n N_Y_c_486_n N_Y_c_529_n N_Y_c_491_n
+ N_Y_c_532_n N_Y_c_495_n N_Y_c_498_n Y N_Y_c_500_n N_Y_c_536_n N_Y_c_503_n
+ N_Y_c_504_n N_Y_c_507_n N_Y_c_538_n N_Y_c_510_n N_Y_c_511_n N_Y_c_512_n
+ N_Y_c_515_n N_Y_c_541_n N_Y_c_518_n N_Y_c_519_n N_Y_c_522_n
+ PM_SKY130_OSU_SC_15T_HS__BUF_8%Y
cc_1 N_GND_M1007_b N_A_M1007_g 0.0645234f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_A_M1007_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_A_M1007_g 0.00388248f $X=0.69 $Y=0.865 $X2=0.475 $Y2=0.895
cc_4 N_GND_c_4_p N_A_M1007_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.475 $Y2=0.895
cc_5 N_GND_M1007_b N_A_M1009_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_6 N_GND_M1007_b N_A_c_210_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.22
cc_7 N_GND_M1007_b N_A_c_211_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.22
cc_8 N_GND_M1007_b N_A_27_115#_M1002_g 0.0255964f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.895
cc_9 N_GND_c_3_p N_A_27_115#_M1002_g 0.00388248f $X=0.69 $Y=0.865 $X2=0.905
+ $Y2=0.895
cc_10 N_GND_c_10_p N_A_27_115#_M1002_g 0.00606474f $X=1.465 $Y=0.152 $X2=0.905
+ $Y2=0.895
cc_11 N_GND_c_4_p N_A_27_115#_M1002_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.905
+ $Y2=0.895
cc_12 N_GND_M1007_b N_A_27_115#_c_249_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.6
cc_13 N_GND_M1007_b N_A_27_115#_M1004_g 0.0245289f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.895
cc_14 N_GND_c_10_p N_A_27_115#_M1004_g 0.00606474f $X=1.465 $Y=0.152 $X2=1.335
+ $Y2=0.895
cc_15 N_GND_c_15_p N_A_27_115#_M1004_g 0.00390533f $X=1.55 $Y=0.865 $X2=1.335
+ $Y2=0.895
cc_16 N_GND_c_4_p N_A_27_115#_M1004_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.335
+ $Y2=0.895
cc_17 N_GND_M1007_b N_A_27_115#_c_254_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.585
cc_18 N_GND_c_15_p N_A_27_115#_c_254_n 0.00256938f $X=1.55 $Y=0.865 $X2=1.69
+ $Y2=1.585
cc_19 N_GND_M1007_b N_A_27_115#_c_256_n 0.0429274f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.585
cc_20 N_GND_M1007_b N_A_27_115#_c_257_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.675
cc_21 N_GND_M1007_b N_A_27_115#_c_258_n 0.0196789f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.675
cc_22 N_GND_M1007_b N_A_27_115#_M1008_g 0.0245289f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.895
cc_23 N_GND_c_15_p N_A_27_115#_M1008_g 0.00390533f $X=1.55 $Y=0.865 $X2=1.765
+ $Y2=0.895
cc_24 N_GND_c_24_p N_A_27_115#_M1008_g 0.00606474f $X=2.325 $Y=0.152 $X2=1.765
+ $Y2=0.895
cc_25 N_GND_c_4_p N_A_27_115#_M1008_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.765
+ $Y2=0.895
cc_26 N_GND_M1007_b N_A_27_115#_c_263_n 0.0195339f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_27 N_GND_M1007_b N_A_27_115#_c_264_n 0.0107618f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.675
cc_28 N_GND_M1007_b N_A_27_115#_M1011_g 0.0245289f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.895
cc_29 N_GND_c_24_p N_A_27_115#_M1011_g 0.00606474f $X=2.325 $Y=0.152 $X2=2.195
+ $Y2=0.895
cc_30 N_GND_c_30_p N_A_27_115#_M1011_g 0.00390533f $X=2.41 $Y=0.865 $X2=2.195
+ $Y2=0.895
cc_31 N_GND_c_4_p N_A_27_115#_M1011_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.195
+ $Y2=0.895
cc_32 N_GND_M1007_b N_A_27_115#_c_269_n 0.0165886f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.585
cc_33 N_GND_c_30_p N_A_27_115#_c_269_n 0.00256938f $X=2.41 $Y=0.865 $X2=2.55
+ $Y2=1.585
cc_34 N_GND_M1007_b N_A_27_115#_c_271_n 0.0109555f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.675
cc_35 N_GND_M1007_b N_A_27_115#_M1012_g 0.0245289f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.895
cc_36 N_GND_c_30_p N_A_27_115#_M1012_g 0.00390533f $X=2.41 $Y=0.865 $X2=2.625
+ $Y2=0.895
cc_37 N_GND_c_37_p N_A_27_115#_M1012_g 0.00606474f $X=3.185 $Y=0.152 $X2=2.625
+ $Y2=0.895
cc_38 N_GND_c_4_p N_A_27_115#_M1012_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.625
+ $Y2=0.895
cc_39 N_GND_M1007_b N_A_27_115#_c_276_n 0.0668243f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.6
cc_40 N_GND_M1007_b N_A_27_115#_c_277_n 0.0195339f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.585
cc_41 N_GND_M1007_b N_A_27_115#_c_278_n 0.0107618f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.675
cc_42 N_GND_M1007_b N_A_27_115#_M1013_g 0.0245289f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.895
cc_43 N_GND_c_37_p N_A_27_115#_M1013_g 0.00606474f $X=3.185 $Y=0.152 $X2=3.055
+ $Y2=0.895
cc_44 N_GND_c_44_p N_A_27_115#_M1013_g 0.00390533f $X=3.27 $Y=0.865 $X2=3.055
+ $Y2=0.895
cc_45 N_GND_c_4_p N_A_27_115#_M1013_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.055
+ $Y2=0.895
cc_46 N_GND_M1007_b N_A_27_115#_c_283_n 0.0215078f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.585
cc_47 N_GND_c_44_p N_A_27_115#_c_283_n 0.00256938f $X=3.27 $Y=0.865 $X2=3.41
+ $Y2=1.585
cc_48 N_GND_M1007_b N_A_27_115#_c_285_n 0.0158747f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.675
cc_49 N_GND_M1007_b N_A_27_115#_M1014_g 0.0245289f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=0.895
cc_50 N_GND_c_44_p N_A_27_115#_M1014_g 0.00390533f $X=3.27 $Y=0.865 $X2=3.485
+ $Y2=0.895
cc_51 N_GND_c_51_p N_A_27_115#_M1014_g 0.00606474f $X=4.045 $Y=0.152 $X2=3.485
+ $Y2=0.895
cc_52 N_GND_c_4_p N_A_27_115#_M1014_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.485
+ $Y2=0.895
cc_53 N_GND_M1007_b N_A_27_115#_c_290_n 0.0385034f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.585
cc_54 N_GND_M1007_b N_A_27_115#_c_291_n 0.0221499f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.675
cc_55 N_GND_M1007_b N_A_27_115#_M1015_g 0.0341369f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=0.895
cc_56 N_GND_c_51_p N_A_27_115#_M1015_g 0.00606474f $X=4.045 $Y=0.152 $X2=3.915
+ $Y2=0.895
cc_57 N_GND_c_57_p N_A_27_115#_M1015_g 0.00866533f $X=4.13 $Y=0.865 $X2=3.915
+ $Y2=0.895
cc_58 N_GND_c_4_p N_A_27_115#_M1015_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.915
+ $Y2=0.895
cc_59 N_GND_M1007_b N_A_27_115#_c_296_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.585
cc_60 N_GND_M1007_b N_A_27_115#_c_297_n 0.00890086f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.675
cc_61 N_GND_M1007_b N_A_27_115#_c_298_n 0.0106787f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.585
cc_62 N_GND_M1007_b N_A_27_115#_c_299_n 0.00890086f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.675
cc_63 N_GND_M1007_b N_A_27_115#_c_300_n 0.0023879f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.585
cc_64 N_GND_M1007_b N_A_27_115#_c_301_n 7.16371e-19 $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.675
cc_65 N_GND_M1007_b N_A_27_115#_c_302_n 0.0106787f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.585
cc_66 N_GND_M1007_b N_A_27_115#_c_303_n 0.00890086f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.675
cc_67 N_GND_M1007_b N_A_27_115#_c_304_n 0.0106787f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.585
cc_68 N_GND_M1007_b N_A_27_115#_c_305_n 0.00890086f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.675
cc_69 N_GND_M1007_b N_A_27_115#_c_306_n 0.0191914f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_70 N_GND_c_2_p N_A_27_115#_c_306_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_71 N_GND_c_4_p N_A_27_115#_c_306_n 0.00476261f $X=3.74 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_72 N_GND_M1007_b N_A_27_115#_c_309_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.205
cc_73 N_GND_M1007_b N_A_27_115#_c_310_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.675
cc_74 N_GND_c_3_p N_A_27_115#_c_310_n 0.00702738f $X=0.69 $Y=0.865 $X2=0.88
+ $Y2=1.675
cc_75 N_GND_M1007_b N_A_27_115#_c_312_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.675
cc_76 N_GND_M1007_b N_A_27_115#_c_313_n 0.00592383f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.675
cc_77 N_GND_M1007_b N_Y_c_477_n 0.00644861f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.865
cc_78 N_GND_c_10_p N_Y_c_477_n 0.00734006f $X=1.465 $Y=0.152 $X2=1.12 $Y2=0.865
cc_79 N_GND_c_15_p N_Y_c_477_n 8.14297e-19 $X=1.55 $Y=0.865 $X2=1.12 $Y2=0.865
cc_80 N_GND_c_4_p N_Y_c_477_n 0.00475776f $X=3.74 $Y=0.19 $X2=1.12 $Y2=0.865
cc_81 N_GND_M1007_b N_Y_c_481_n 0.00656459f $X=-0.045 $Y=0 $X2=1.98 $Y2=0.865
cc_82 N_GND_c_15_p N_Y_c_481_n 8.14297e-19 $X=1.55 $Y=0.865 $X2=1.98 $Y2=0.865
cc_83 N_GND_c_24_p N_Y_c_481_n 0.00754406f $X=2.325 $Y=0.152 $X2=1.98 $Y2=0.865
cc_84 N_GND_c_30_p N_Y_c_481_n 8.14297e-19 $X=2.41 $Y=0.865 $X2=1.98 $Y2=0.865
cc_85 N_GND_c_4_p N_Y_c_481_n 0.00475776f $X=3.74 $Y=0.19 $X2=1.98 $Y2=0.865
cc_86 N_GND_M1007_b N_Y_c_486_n 0.00656459f $X=-0.045 $Y=0 $X2=2.84 $Y2=0.865
cc_87 N_GND_c_30_p N_Y_c_486_n 8.14297e-19 $X=2.41 $Y=0.865 $X2=2.84 $Y2=0.865
cc_88 N_GND_c_37_p N_Y_c_486_n 0.00746708f $X=3.185 $Y=0.152 $X2=2.84 $Y2=0.865
cc_89 N_GND_c_44_p N_Y_c_486_n 8.14297e-19 $X=3.27 $Y=0.865 $X2=2.84 $Y2=0.865
cc_90 N_GND_c_4_p N_Y_c_486_n 0.00475776f $X=3.74 $Y=0.19 $X2=2.84 $Y2=0.865
cc_91 N_GND_M1007_b N_Y_c_491_n 0.00656459f $X=-0.045 $Y=0 $X2=3.7 $Y2=0.865
cc_92 N_GND_c_44_p N_Y_c_491_n 8.14297e-19 $X=3.27 $Y=0.865 $X2=3.7 $Y2=0.865
cc_93 N_GND_c_51_p N_Y_c_491_n 0.00734006f $X=4.045 $Y=0.152 $X2=3.7 $Y2=0.865
cc_94 N_GND_c_4_p N_Y_c_491_n 0.00475776f $X=3.74 $Y=0.19 $X2=3.7 $Y2=0.865
cc_95 N_GND_M1007_b N_Y_c_495_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.335
cc_96 N_GND_c_3_p N_Y_c_495_n 0.00134236f $X=0.69 $Y=0.865 $X2=1.12 $Y2=1.335
cc_97 N_GND_c_15_p N_Y_c_495_n 7.53951e-19 $X=1.55 $Y=0.865 $X2=1.12 $Y2=1.335
cc_98 N_GND_M1007_b N_Y_c_498_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.585
cc_99 N_GND_M1007_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=2.01
cc_100 N_GND_M1004_s N_Y_c_500_n 0.00418405f $X=1.41 $Y=0.575 $X2=1.835 $Y2=1.22
cc_101 N_GND_M1007_b N_Y_c_500_n 0.00793787f $X=-0.045 $Y=0 $X2=1.835 $Y2=1.22
cc_102 N_GND_c_15_p N_Y_c_500_n 0.0142303f $X=1.55 $Y=0.865 $X2=1.835 $Y2=1.22
cc_103 N_GND_M1007_b N_Y_c_503_n 0.0437239f $X=-0.045 $Y=0 $X2=1.98 $Y2=2.585
cc_104 N_GND_M1011_s N_Y_c_504_n 0.00418405f $X=2.27 $Y=0.575 $X2=2.695 $Y2=1.22
cc_105 N_GND_M1007_b N_Y_c_504_n 0.00793787f $X=-0.045 $Y=0 $X2=2.695 $Y2=1.22
cc_106 N_GND_c_30_p N_Y_c_504_n 0.0142303f $X=2.41 $Y=0.865 $X2=2.695 $Y2=1.22
cc_107 N_GND_M1007_b N_Y_c_507_n 0.00409378f $X=-0.045 $Y=0 $X2=2.125 $Y2=1.22
cc_108 N_GND_c_15_p N_Y_c_507_n 7.53951e-19 $X=1.55 $Y=0.865 $X2=2.125 $Y2=1.22
cc_109 N_GND_c_30_p N_Y_c_507_n 7.53951e-19 $X=2.41 $Y=0.865 $X2=2.125 $Y2=1.22
cc_110 N_GND_M1007_b N_Y_c_510_n 0.00560779f $X=-0.045 $Y=0 $X2=2.125 $Y2=2.7
cc_111 N_GND_M1007_b N_Y_c_511_n 0.0575129f $X=-0.045 $Y=0 $X2=2.84 $Y2=2.585
cc_112 N_GND_M1013_s N_Y_c_512_n 0.00418405f $X=3.13 $Y=0.575 $X2=3.555 $Y2=1.22
cc_113 N_GND_M1007_b N_Y_c_512_n 0.00793787f $X=-0.045 $Y=0 $X2=3.555 $Y2=1.22
cc_114 N_GND_c_44_p N_Y_c_512_n 0.0142303f $X=3.27 $Y=0.865 $X2=3.555 $Y2=1.22
cc_115 N_GND_M1007_b N_Y_c_515_n 0.00409378f $X=-0.045 $Y=0 $X2=2.985 $Y2=1.22
cc_116 N_GND_c_30_p N_Y_c_515_n 7.53951e-19 $X=2.41 $Y=0.865 $X2=2.985 $Y2=1.22
cc_117 N_GND_c_44_p N_Y_c_515_n 7.53951e-19 $X=3.27 $Y=0.865 $X2=2.985 $Y2=1.22
cc_118 N_GND_M1007_b N_Y_c_518_n 0.00485078f $X=-0.045 $Y=0 $X2=2.985 $Y2=2.7
cc_119 N_GND_M1007_b N_Y_c_519_n 0.00409378f $X=-0.045 $Y=0 $X2=3.7 $Y2=1.335
cc_120 N_GND_c_44_p N_Y_c_519_n 7.53951e-19 $X=3.27 $Y=0.865 $X2=3.7 $Y2=1.335
cc_121 N_GND_c_57_p N_Y_c_519_n 0.00134236f $X=4.13 $Y=0.865 $X2=3.7 $Y2=1.335
cc_122 N_GND_M1007_b N_Y_c_522_n 0.0800785f $X=-0.045 $Y=0 $X2=3.7 $Y2=2.585
cc_123 N_VDD_M1009_b N_A_M1009_g 0.024954f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_124 N_VDD_c_124_p N_A_M1009_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_125 N_VDD_c_125_p N_A_M1009_g 0.00362996f $X=0.69 $Y=3.885 $X2=0.475
+ $Y2=3.825
cc_126 N_VDD_c_126_p N_A_M1009_g 0.00429146f $X=3.74 $Y=5.36 $X2=0.475 $Y2=3.825
cc_127 N_VDD_M1009_d N_A_c_211_n 0.00628533f $X=0.55 $Y=2.825 $X2=0.635 $Y2=2.22
cc_128 N_VDD_M1009_b N_A_c_211_n 0.00328912f $X=-0.045 $Y=2.645 $X2=0.635
+ $Y2=2.22
cc_129 N_VDD_c_125_p N_A_c_211_n 0.00264661f $X=0.69 $Y=3.885 $X2=0.635 $Y2=2.22
cc_130 N_VDD_M1009_d A 0.00797576f $X=0.55 $Y=2.825 $X2=0.635 $Y2=3.07
cc_131 N_VDD_c_125_p A 0.00510982f $X=0.69 $Y=3.885 $X2=0.635 $Y2=3.07
cc_132 N_VDD_M1009_b N_A_27_115#_c_314_n 0.01464f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=2.75
cc_133 N_VDD_c_125_p N_A_27_115#_c_314_n 0.00362996f $X=0.69 $Y=3.885 $X2=0.905
+ $Y2=2.75
cc_134 N_VDD_c_134_p N_A_27_115#_c_314_n 0.00496961f $X=1.465 $Y=5.397 $X2=0.905
+ $Y2=2.75
cc_135 N_VDD_c_126_p N_A_27_115#_c_314_n 0.00429146f $X=3.74 $Y=5.36 $X2=0.905
+ $Y2=2.75
cc_136 N_VDD_M1009_b N_A_27_115#_c_318_n 0.0144912f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.75
cc_137 N_VDD_c_125_p N_A_27_115#_c_318_n 3.67508e-19 $X=0.69 $Y=3.885 $X2=1.335
+ $Y2=2.75
cc_138 N_VDD_c_134_p N_A_27_115#_c_318_n 0.00500229f $X=1.465 $Y=5.397 $X2=1.335
+ $Y2=2.75
cc_139 N_VDD_c_139_p N_A_27_115#_c_318_n 0.00382402f $X=1.55 $Y=3.205 $X2=1.335
+ $Y2=2.75
cc_140 N_VDD_c_126_p N_A_27_115#_c_318_n 0.00430409f $X=3.74 $Y=5.36 $X2=1.335
+ $Y2=2.75
cc_141 N_VDD_M1009_b N_A_27_115#_c_257_n 0.00647677f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.675
cc_142 N_VDD_c_139_p N_A_27_115#_c_257_n 0.00364479f $X=1.55 $Y=3.205 $X2=1.69
+ $Y2=2.675
cc_143 N_VDD_M1009_b N_A_27_115#_c_258_n 0.0113915f $X=-0.045 $Y=2.645 $X2=1.41
+ $Y2=2.675
cc_144 N_VDD_M1009_b N_A_27_115#_c_326_n 0.0141812f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.75
cc_145 N_VDD_c_139_p N_A_27_115#_c_326_n 0.00362996f $X=1.55 $Y=3.205 $X2=1.765
+ $Y2=2.75
cc_146 N_VDD_c_146_p N_A_27_115#_c_326_n 0.00496961f $X=2.325 $Y=5.397 $X2=1.765
+ $Y2=2.75
cc_147 N_VDD_c_126_p N_A_27_115#_c_326_n 0.00429146f $X=3.74 $Y=5.36 $X2=1.765
+ $Y2=2.75
cc_148 N_VDD_M1009_b N_A_27_115#_c_264_n 0.00596183f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.675
cc_149 N_VDD_M1009_b N_A_27_115#_c_331_n 0.0141812f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.75
cc_150 N_VDD_c_146_p N_A_27_115#_c_331_n 0.00496961f $X=2.325 $Y=5.397 $X2=2.195
+ $Y2=2.75
cc_151 N_VDD_c_151_p N_A_27_115#_c_331_n 0.00362996f $X=2.41 $Y=3.205 $X2=2.195
+ $Y2=2.75
cc_152 N_VDD_c_126_p N_A_27_115#_c_331_n 0.00429146f $X=3.74 $Y=5.36 $X2=2.195
+ $Y2=2.75
cc_153 N_VDD_M1009_b N_A_27_115#_c_271_n 0.00647677f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.675
cc_154 N_VDD_c_151_p N_A_27_115#_c_271_n 0.00364479f $X=2.41 $Y=3.205 $X2=2.55
+ $Y2=2.675
cc_155 N_VDD_M1009_b N_A_27_115#_c_337_n 0.0141812f $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.75
cc_156 N_VDD_c_151_p N_A_27_115#_c_337_n 0.00362996f $X=2.41 $Y=3.205 $X2=2.625
+ $Y2=2.75
cc_157 N_VDD_c_157_p N_A_27_115#_c_337_n 0.00496961f $X=3.185 $Y=5.397 $X2=2.625
+ $Y2=2.75
cc_158 N_VDD_c_126_p N_A_27_115#_c_337_n 0.00429146f $X=3.74 $Y=5.36 $X2=2.625
+ $Y2=2.75
cc_159 N_VDD_M1009_b N_A_27_115#_c_278_n 0.00596183f $X=-0.045 $Y=2.645 $X2=2.98
+ $Y2=2.675
cc_160 N_VDD_M1009_b N_A_27_115#_c_342_n 0.0141812f $X=-0.045 $Y=2.645 $X2=3.055
+ $Y2=2.75
cc_161 N_VDD_c_157_p N_A_27_115#_c_342_n 0.00496961f $X=3.185 $Y=5.397 $X2=3.055
+ $Y2=2.75
cc_162 N_VDD_c_162_p N_A_27_115#_c_342_n 0.00362996f $X=3.27 $Y=3.205 $X2=3.055
+ $Y2=2.75
cc_163 N_VDD_c_126_p N_A_27_115#_c_342_n 0.00429146f $X=3.74 $Y=5.36 $X2=3.055
+ $Y2=2.75
cc_164 N_VDD_M1009_b N_A_27_115#_c_285_n 0.00647677f $X=-0.045 $Y=2.645 $X2=3.41
+ $Y2=2.675
cc_165 N_VDD_c_162_p N_A_27_115#_c_285_n 0.00364479f $X=3.27 $Y=3.205 $X2=3.41
+ $Y2=2.675
cc_166 N_VDD_M1009_b N_A_27_115#_c_348_n 0.0141812f $X=-0.045 $Y=2.645 $X2=3.485
+ $Y2=2.75
cc_167 N_VDD_c_162_p N_A_27_115#_c_348_n 0.00362996f $X=3.27 $Y=3.205 $X2=3.485
+ $Y2=2.75
cc_168 N_VDD_c_168_p N_A_27_115#_c_348_n 0.00496961f $X=4.045 $Y=5.397 $X2=3.485
+ $Y2=2.75
cc_169 N_VDD_c_126_p N_A_27_115#_c_348_n 0.00429146f $X=3.74 $Y=5.36 $X2=3.485
+ $Y2=2.75
cc_170 N_VDD_M1009_b N_A_27_115#_c_291_n 0.0134369f $X=-0.045 $Y=2.645 $X2=3.84
+ $Y2=2.675
cc_171 N_VDD_M1009_b N_A_27_115#_c_353_n 0.017048f $X=-0.045 $Y=2.645 $X2=3.915
+ $Y2=2.75
cc_172 N_VDD_c_168_p N_A_27_115#_c_353_n 0.00496961f $X=4.045 $Y=5.397 $X2=3.915
+ $Y2=2.75
cc_173 N_VDD_c_173_p N_A_27_115#_c_353_n 0.00751602f $X=4.13 $Y=3.205 $X2=3.915
+ $Y2=2.75
cc_174 N_VDD_c_126_p N_A_27_115#_c_353_n 0.00429146f $X=3.74 $Y=5.36 $X2=3.915
+ $Y2=2.75
cc_175 N_VDD_M1009_b N_A_27_115#_c_297_n 0.00167153f $X=-0.045 $Y=2.645
+ $X2=1.765 $Y2=2.675
cc_176 N_VDD_M1009_b N_A_27_115#_c_299_n 0.00167153f $X=-0.045 $Y=2.645
+ $X2=2.195 $Y2=2.675
cc_177 N_VDD_M1009_b N_A_27_115#_c_301_n 0.00167153f $X=-0.045 $Y=2.645
+ $X2=2.625 $Y2=2.675
cc_178 N_VDD_M1009_b N_A_27_115#_c_303_n 0.00167153f $X=-0.045 $Y=2.645
+ $X2=3.055 $Y2=2.675
cc_179 N_VDD_M1009_b N_A_27_115#_c_305_n 0.00167153f $X=-0.045 $Y=2.645
+ $X2=3.485 $Y2=2.675
cc_180 N_VDD_M1009_b N_A_27_115#_c_309_n 0.0103979f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.205
cc_181 N_VDD_c_124_p N_A_27_115#_c_309_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.205
cc_182 N_VDD_c_126_p N_A_27_115#_c_309_n 0.00435496f $X=3.74 $Y=5.36 $X2=0.26
+ $Y2=3.205
cc_183 N_VDD_M1009_b N_Y_c_523_n 0.00333732f $X=-0.045 $Y=2.645 $X2=1.12 $Y2=2.7
cc_184 N_VDD_c_134_p N_Y_c_523_n 0.0045126f $X=1.465 $Y=5.397 $X2=1.12 $Y2=2.7
cc_185 N_VDD_c_126_p N_Y_c_523_n 0.00434939f $X=3.74 $Y=5.36 $X2=1.12 $Y2=2.7
cc_186 N_VDD_M1009_b N_Y_c_526_n 0.00381442f $X=-0.045 $Y=2.645 $X2=1.98 $Y2=2.7
cc_187 N_VDD_c_146_p N_Y_c_526_n 0.00474282f $X=2.325 $Y=5.397 $X2=1.98 $Y2=2.7
cc_188 N_VDD_c_126_p N_Y_c_526_n 0.00434939f $X=3.74 $Y=5.36 $X2=1.98 $Y2=2.7
cc_189 N_VDD_M1009_b N_Y_c_529_n 0.00381442f $X=-0.045 $Y=2.645 $X2=2.84 $Y2=2.7
cc_190 N_VDD_c_157_p N_Y_c_529_n 0.00465594f $X=3.185 $Y=5.397 $X2=2.84 $Y2=2.7
cc_191 N_VDD_c_126_p N_Y_c_529_n 0.00434939f $X=3.74 $Y=5.36 $X2=2.84 $Y2=2.7
cc_192 N_VDD_M1009_b N_Y_c_532_n 0.00381442f $X=-0.045 $Y=2.645 $X2=3.7 $Y2=2.7
cc_193 N_VDD_c_168_p N_Y_c_532_n 0.0045126f $X=4.045 $Y=5.397 $X2=3.7 $Y2=2.7
cc_194 N_VDD_c_126_p N_Y_c_532_n 0.00434939f $X=3.74 $Y=5.36 $X2=3.7 $Y2=2.7
cc_195 N_VDD_M1009_b N_Y_c_498_n 0.00409378f $X=-0.045 $Y=2.645 $X2=1.12
+ $Y2=2.585
cc_196 N_VDD_M1009_b N_Y_c_536_n 0.00520877f $X=-0.045 $Y=2.645 $X2=1.835
+ $Y2=2.7
cc_197 N_VDD_c_139_p N_Y_c_536_n 0.0090257f $X=1.55 $Y=3.205 $X2=1.835 $Y2=2.7
cc_198 N_VDD_M1009_b N_Y_c_538_n 0.00520877f $X=-0.045 $Y=2.645 $X2=2.695
+ $Y2=2.7
cc_199 N_VDD_c_151_p N_Y_c_538_n 0.0090257f $X=2.41 $Y=3.205 $X2=2.695 $Y2=2.7
cc_200 N_VDD_M1009_b N_Y_c_510_n 0.00409378f $X=-0.045 $Y=2.645 $X2=2.125
+ $Y2=2.7
cc_201 N_VDD_M1009_b N_Y_c_541_n 0.00520877f $X=-0.045 $Y=2.645 $X2=3.555
+ $Y2=2.7
cc_202 N_VDD_c_162_p N_Y_c_541_n 0.0090257f $X=3.27 $Y=3.205 $X2=3.555 $Y2=2.7
cc_203 N_VDD_M1009_b N_Y_c_518_n 0.00409378f $X=-0.045 $Y=2.645 $X2=2.985
+ $Y2=2.7
cc_204 N_VDD_M1009_b N_Y_c_522_n 0.00409378f $X=-0.045 $Y=2.645 $X2=3.7
+ $Y2=2.585
cc_205 A N_A_27_115#_M1009_s 0.00414531f $X=0.635 $Y=3.07 $X2=0.135 $Y2=2.825
cc_206 N_A_M1007_g N_A_27_115#_M1002_g 0.0415224f $X=0.475 $Y=0.895 $X2=0.905
+ $Y2=0.895
cc_207 A N_A_27_115#_c_314_n 0.00419145f $X=0.635 $Y=3.07 $X2=0.905 $Y2=2.75
cc_208 N_A_M1007_g N_A_27_115#_c_249_n 0.00260138f $X=0.475 $Y=0.895 $X2=1.18
+ $Y2=2.6
cc_209 N_A_M1009_g N_A_27_115#_c_249_n 0.00209773f $X=0.475 $Y=3.825 $X2=1.18
+ $Y2=2.6
cc_210 N_A_c_210_n N_A_27_115#_c_249_n 0.0139096f $X=0.635 $Y=2.22 $X2=1.18
+ $Y2=2.6
cc_211 N_A_c_211_n N_A_27_115#_c_249_n 0.00361737f $X=0.635 $Y=2.22 $X2=1.18
+ $Y2=2.6
cc_212 N_A_M1009_g N_A_27_115#_c_258_n 0.0506363f $X=0.475 $Y=3.825 $X2=1.41
+ $Y2=2.675
cc_213 N_A_c_211_n N_A_27_115#_c_258_n 0.00477416f $X=0.635 $Y=2.22 $X2=1.41
+ $Y2=2.675
cc_214 N_A_M1007_g N_A_27_115#_c_306_n 0.0183389f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=0.865
cc_215 N_A_M1007_g N_A_27_115#_c_309_n 0.0341146f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=3.205
cc_216 N_A_c_211_n N_A_27_115#_c_309_n 0.0548951f $X=0.635 $Y=2.22 $X2=0.26
+ $Y2=3.205
cc_217 A N_A_27_115#_c_309_n 0.0155137f $X=0.635 $Y=3.07 $X2=0.26 $Y2=3.205
cc_218 N_A_M1007_g N_A_27_115#_c_310_n 0.0207696f $X=0.475 $Y=0.895 $X2=0.88
+ $Y2=1.675
cc_219 N_A_c_210_n N_A_27_115#_c_310_n 0.00273049f $X=0.635 $Y=2.22 $X2=0.88
+ $Y2=1.675
cc_220 N_A_c_211_n N_A_27_115#_c_310_n 0.00886797f $X=0.635 $Y=2.22 $X2=0.88
+ $Y2=1.675
cc_221 N_A_M1007_g N_A_27_115#_c_313_n 6.59135e-19 $X=0.475 $Y=0.895 $X2=0.965
+ $Y2=1.675
cc_222 N_A_c_211_n N_Y_c_523_n 0.0135622f $X=0.635 $Y=2.22 $X2=1.12 $Y2=2.7
cc_223 A N_Y_c_523_n 0.00731851f $X=0.635 $Y=3.07 $X2=1.12 $Y2=2.7
cc_224 N_A_M1007_g N_Y_c_495_n 8.23842e-19 $X=0.475 $Y=0.895 $X2=1.12 $Y2=1.335
cc_225 N_A_c_211_n N_Y_c_498_n 0.00677552f $X=0.635 $Y=2.22 $X2=1.12 $Y2=2.585
cc_226 N_A_M1007_g Y 0.00310306f $X=0.475 $Y=0.895 $X2=1.055 $Y2=2.01
cc_227 N_A_c_210_n Y 0.00441844f $X=0.635 $Y=2.22 $X2=1.055 $Y2=2.01
cc_228 N_A_c_211_n Y 0.0200396f $X=0.635 $Y=2.22 $X2=1.055 $Y2=2.01
cc_229 N_A_27_115#_M1002_g N_Y_c_477_n 0.00339663f $X=0.905 $Y=0.895 $X2=1.12
+ $Y2=0.865
cc_230 N_A_27_115#_M1004_g N_Y_c_477_n 0.00339663f $X=1.335 $Y=0.895 $X2=1.12
+ $Y2=0.865
cc_231 N_A_27_115#_c_256_n N_Y_c_477_n 0.0030245f $X=1.41 $Y=1.585 $X2=1.12
+ $Y2=0.865
cc_232 N_A_27_115#_c_313_n N_Y_c_477_n 7.50437e-19 $X=0.965 $Y=1.675 $X2=1.12
+ $Y2=0.865
cc_233 N_A_27_115#_c_314_n N_Y_c_523_n 0.00163525f $X=0.905 $Y=2.75 $X2=1.12
+ $Y2=2.7
cc_234 N_A_27_115#_c_318_n N_Y_c_523_n 0.00258898f $X=1.335 $Y=2.75 $X2=1.12
+ $Y2=2.7
cc_235 N_A_27_115#_c_258_n N_Y_c_523_n 0.0126676f $X=1.41 $Y=2.675 $X2=1.12
+ $Y2=2.7
cc_236 N_A_27_115#_M1008_g N_Y_c_481_n 0.00339663f $X=1.765 $Y=0.895 $X2=1.98
+ $Y2=0.865
cc_237 N_A_27_115#_c_263_n N_Y_c_481_n 0.00280419f $X=2.12 $Y=1.585 $X2=1.98
+ $Y2=0.865
cc_238 N_A_27_115#_M1011_g N_Y_c_481_n 0.00339663f $X=2.195 $Y=0.895 $X2=1.98
+ $Y2=0.865
cc_239 N_A_27_115#_c_326_n N_Y_c_526_n 0.00258898f $X=1.765 $Y=2.75 $X2=1.98
+ $Y2=2.7
cc_240 N_A_27_115#_c_264_n N_Y_c_526_n 0.0138847f $X=2.12 $Y=2.675 $X2=1.98
+ $Y2=2.7
cc_241 N_A_27_115#_c_331_n N_Y_c_526_n 0.00258898f $X=2.195 $Y=2.75 $X2=1.98
+ $Y2=2.7
cc_242 N_A_27_115#_M1012_g N_Y_c_486_n 0.00339663f $X=2.625 $Y=0.895 $X2=2.84
+ $Y2=0.865
cc_243 N_A_27_115#_c_277_n N_Y_c_486_n 0.00280419f $X=2.98 $Y=1.585 $X2=2.84
+ $Y2=0.865
cc_244 N_A_27_115#_M1013_g N_Y_c_486_n 0.00339663f $X=3.055 $Y=0.895 $X2=2.84
+ $Y2=0.865
cc_245 N_A_27_115#_c_337_n N_Y_c_529_n 0.00258898f $X=2.625 $Y=2.75 $X2=2.84
+ $Y2=2.7
cc_246 N_A_27_115#_c_278_n N_Y_c_529_n 0.0138847f $X=2.98 $Y=2.675 $X2=2.84
+ $Y2=2.7
cc_247 N_A_27_115#_c_342_n N_Y_c_529_n 0.00258898f $X=3.055 $Y=2.75 $X2=2.84
+ $Y2=2.7
cc_248 N_A_27_115#_M1014_g N_Y_c_491_n 0.00339663f $X=3.485 $Y=0.895 $X2=3.7
+ $Y2=0.865
cc_249 N_A_27_115#_c_290_n N_Y_c_491_n 0.00280419f $X=3.84 $Y=1.585 $X2=3.7
+ $Y2=0.865
cc_250 N_A_27_115#_M1015_g N_Y_c_491_n 0.00339663f $X=3.915 $Y=0.895 $X2=3.7
+ $Y2=0.865
cc_251 N_A_27_115#_c_348_n N_Y_c_532_n 0.00258898f $X=3.485 $Y=2.75 $X2=3.7
+ $Y2=2.7
cc_252 N_A_27_115#_c_291_n N_Y_c_532_n 0.013404f $X=3.84 $Y=2.675 $X2=3.7
+ $Y2=2.7
cc_253 N_A_27_115#_c_353_n N_Y_c_532_n 0.00258898f $X=3.915 $Y=2.75 $X2=3.7
+ $Y2=2.7
cc_254 N_A_27_115#_M1002_g N_Y_c_495_n 0.00541983f $X=0.905 $Y=0.895 $X2=1.12
+ $Y2=1.335
cc_255 N_A_27_115#_M1004_g N_Y_c_495_n 0.00262362f $X=1.335 $Y=0.895 $X2=1.12
+ $Y2=1.335
cc_256 N_A_27_115#_c_313_n N_Y_c_495_n 0.00278861f $X=0.965 $Y=1.675 $X2=1.12
+ $Y2=1.335
cc_257 N_A_27_115#_c_314_n N_Y_c_498_n 0.00120715f $X=0.905 $Y=2.75 $X2=1.12
+ $Y2=2.585
cc_258 N_A_27_115#_c_249_n N_Y_c_498_n 0.00215118f $X=1.18 $Y=2.6 $X2=1.12
+ $Y2=2.585
cc_259 N_A_27_115#_c_318_n N_Y_c_498_n 0.00113627f $X=1.335 $Y=2.75 $X2=1.12
+ $Y2=2.585
cc_260 N_A_27_115#_c_258_n N_Y_c_498_n 0.00372325f $X=1.41 $Y=2.675 $X2=1.12
+ $Y2=2.585
cc_261 N_A_27_115#_M1002_g Y 0.00251111f $X=0.905 $Y=0.895 $X2=1.055 $Y2=2.01
cc_262 N_A_27_115#_c_249_n Y 0.0314621f $X=1.18 $Y=2.6 $X2=1.055 $Y2=2.01
cc_263 N_A_27_115#_M1004_g Y 0.00251111f $X=1.335 $Y=0.895 $X2=1.055 $Y2=2.01
cc_264 N_A_27_115#_c_256_n Y 0.0166018f $X=1.41 $Y=1.585 $X2=1.055 $Y2=2.01
cc_265 N_A_27_115#_c_310_n Y 8.73078e-19 $X=0.88 $Y=1.675 $X2=1.055 $Y2=2.01
cc_266 N_A_27_115#_c_313_n Y 0.0121742f $X=0.965 $Y=1.675 $X2=1.055 $Y2=2.01
cc_267 N_A_27_115#_M1004_g N_Y_c_500_n 0.0133661f $X=1.335 $Y=0.895 $X2=1.835
+ $Y2=1.22
cc_268 N_A_27_115#_c_254_n N_Y_c_500_n 0.00213861f $X=1.69 $Y=1.585 $X2=1.835
+ $Y2=1.22
cc_269 N_A_27_115#_M1008_g N_Y_c_500_n 0.0130095f $X=1.765 $Y=0.895 $X2=1.835
+ $Y2=1.22
cc_270 N_A_27_115#_c_318_n N_Y_c_536_n 0.00639369f $X=1.335 $Y=2.75 $X2=1.835
+ $Y2=2.7
cc_271 N_A_27_115#_c_257_n N_Y_c_536_n 0.0125005f $X=1.69 $Y=2.675 $X2=1.835
+ $Y2=2.7
cc_272 N_A_27_115#_c_258_n N_Y_c_536_n 0.00627763f $X=1.41 $Y=2.675 $X2=1.835
+ $Y2=2.7
cc_273 N_A_27_115#_c_326_n N_Y_c_536_n 0.00639369f $X=1.765 $Y=2.75 $X2=1.835
+ $Y2=2.7
cc_274 N_A_27_115#_c_297_n N_Y_c_536_n 0.00580646f $X=1.765 $Y=2.675 $X2=1.835
+ $Y2=2.7
cc_275 N_A_27_115#_c_256_n N_Y_c_503_n 0.013329f $X=1.41 $Y=1.585 $X2=1.98
+ $Y2=2.585
cc_276 N_A_27_115#_M1008_g N_Y_c_503_n 0.00251111f $X=1.765 $Y=0.895 $X2=1.98
+ $Y2=2.585
cc_277 N_A_27_115#_c_263_n N_Y_c_503_n 0.0178059f $X=2.12 $Y=1.585 $X2=1.98
+ $Y2=2.585
cc_278 N_A_27_115#_M1011_g N_Y_c_503_n 0.00251111f $X=2.195 $Y=0.895 $X2=1.98
+ $Y2=2.585
cc_279 N_A_27_115#_c_276_n N_Y_c_503_n 0.0137936f $X=2.625 $Y=2.6 $X2=1.98
+ $Y2=2.585
cc_280 N_A_27_115#_M1011_g N_Y_c_504_n 0.0130095f $X=2.195 $Y=0.895 $X2=2.695
+ $Y2=1.22
cc_281 N_A_27_115#_c_269_n N_Y_c_504_n 0.00213861f $X=2.55 $Y=1.585 $X2=2.695
+ $Y2=1.22
cc_282 N_A_27_115#_M1012_g N_Y_c_504_n 0.0136594f $X=2.625 $Y=0.895 $X2=2.695
+ $Y2=1.22
cc_283 N_A_27_115#_M1008_g N_Y_c_507_n 0.00259902f $X=1.765 $Y=0.895 $X2=2.125
+ $Y2=1.22
cc_284 N_A_27_115#_M1011_g N_Y_c_507_n 0.00259902f $X=2.195 $Y=0.895 $X2=2.125
+ $Y2=1.22
cc_285 N_A_27_115#_c_331_n N_Y_c_538_n 0.00639369f $X=2.195 $Y=2.75 $X2=2.695
+ $Y2=2.7
cc_286 N_A_27_115#_c_271_n N_Y_c_538_n 0.0130313f $X=2.55 $Y=2.675 $X2=2.695
+ $Y2=2.7
cc_287 N_A_27_115#_c_337_n N_Y_c_538_n 0.00639369f $X=2.625 $Y=2.75 $X2=2.695
+ $Y2=2.7
cc_288 N_A_27_115#_c_299_n N_Y_c_538_n 0.00580646f $X=2.195 $Y=2.675 $X2=2.695
+ $Y2=2.7
cc_289 N_A_27_115#_c_301_n N_Y_c_538_n 0.00666531f $X=2.625 $Y=2.675 $X2=2.695
+ $Y2=2.7
cc_290 N_A_27_115#_c_326_n N_Y_c_510_n 0.00113627f $X=1.765 $Y=2.75 $X2=2.125
+ $Y2=2.7
cc_291 N_A_27_115#_c_264_n N_Y_c_510_n 0.00364679f $X=2.12 $Y=2.675 $X2=2.125
+ $Y2=2.7
cc_292 N_A_27_115#_c_331_n N_Y_c_510_n 0.00113627f $X=2.195 $Y=2.75 $X2=2.125
+ $Y2=2.7
cc_293 N_A_27_115#_c_297_n N_Y_c_510_n 6.99501e-19 $X=1.765 $Y=2.675 $X2=2.125
+ $Y2=2.7
cc_294 N_A_27_115#_c_299_n N_Y_c_510_n 6.99501e-19 $X=2.195 $Y=2.675 $X2=2.125
+ $Y2=2.7
cc_295 N_A_27_115#_M1012_g N_Y_c_511_n 0.00251111f $X=2.625 $Y=0.895 $X2=2.84
+ $Y2=2.585
cc_296 N_A_27_115#_c_276_n N_Y_c_511_n 0.017762f $X=2.625 $Y=2.6 $X2=2.84
+ $Y2=2.585
cc_297 N_A_27_115#_c_277_n N_Y_c_511_n 0.0178059f $X=2.98 $Y=1.585 $X2=2.84
+ $Y2=2.585
cc_298 N_A_27_115#_M1013_g N_Y_c_511_n 0.00251111f $X=3.055 $Y=0.895 $X2=2.84
+ $Y2=2.585
cc_299 N_A_27_115#_M1013_g N_Y_c_512_n 0.0130095f $X=3.055 $Y=0.895 $X2=3.555
+ $Y2=1.22
cc_300 N_A_27_115#_c_283_n N_Y_c_512_n 0.00213861f $X=3.41 $Y=1.585 $X2=3.555
+ $Y2=1.22
cc_301 N_A_27_115#_M1014_g N_Y_c_512_n 0.0130095f $X=3.485 $Y=0.895 $X2=3.555
+ $Y2=1.22
cc_302 N_A_27_115#_M1012_g N_Y_c_515_n 0.00262362f $X=2.625 $Y=0.895 $X2=2.985
+ $Y2=1.22
cc_303 N_A_27_115#_M1013_g N_Y_c_515_n 0.00259902f $X=3.055 $Y=0.895 $X2=2.985
+ $Y2=1.22
cc_304 N_A_27_115#_c_342_n N_Y_c_541_n 0.00639369f $X=3.055 $Y=2.75 $X2=3.555
+ $Y2=2.7
cc_305 N_A_27_115#_c_285_n N_Y_c_541_n 0.0125005f $X=3.41 $Y=2.675 $X2=3.555
+ $Y2=2.7
cc_306 N_A_27_115#_c_348_n N_Y_c_541_n 0.00639369f $X=3.485 $Y=2.75 $X2=3.555
+ $Y2=2.7
cc_307 N_A_27_115#_c_303_n N_Y_c_541_n 0.00580646f $X=3.055 $Y=2.675 $X2=3.555
+ $Y2=2.7
cc_308 N_A_27_115#_c_305_n N_Y_c_541_n 0.00580646f $X=3.485 $Y=2.675 $X2=3.555
+ $Y2=2.7
cc_309 N_A_27_115#_c_276_n N_Y_c_518_n 8.30534e-19 $X=2.625 $Y=2.6 $X2=2.985
+ $Y2=2.7
cc_310 N_A_27_115#_c_337_n N_Y_c_518_n 0.00113627f $X=2.625 $Y=2.75 $X2=2.985
+ $Y2=2.7
cc_311 N_A_27_115#_c_278_n N_Y_c_518_n 0.00364679f $X=2.98 $Y=2.675 $X2=2.985
+ $Y2=2.7
cc_312 N_A_27_115#_c_342_n N_Y_c_518_n 0.00113627f $X=3.055 $Y=2.75 $X2=2.985
+ $Y2=2.7
cc_313 N_A_27_115#_c_301_n N_Y_c_518_n 6.59375e-19 $X=2.625 $Y=2.675 $X2=2.985
+ $Y2=2.7
cc_314 N_A_27_115#_c_303_n N_Y_c_518_n 6.99501e-19 $X=3.055 $Y=2.675 $X2=2.985
+ $Y2=2.7
cc_315 N_A_27_115#_M1014_g N_Y_c_519_n 0.00259902f $X=3.485 $Y=0.895 $X2=3.7
+ $Y2=1.335
cc_316 N_A_27_115#_M1015_g N_Y_c_519_n 0.00939545f $X=3.915 $Y=0.895 $X2=3.7
+ $Y2=1.335
cc_317 N_A_27_115#_M1014_g N_Y_c_522_n 0.00251111f $X=3.485 $Y=0.895 $X2=3.7
+ $Y2=2.585
cc_318 N_A_27_115#_c_348_n N_Y_c_522_n 0.00113627f $X=3.485 $Y=2.75 $X2=3.7
+ $Y2=2.585
cc_319 N_A_27_115#_c_290_n N_Y_c_522_n 0.0170354f $X=3.84 $Y=1.585 $X2=3.7
+ $Y2=2.585
cc_320 N_A_27_115#_c_291_n N_Y_c_522_n 0.00966211f $X=3.84 $Y=2.675 $X2=3.7
+ $Y2=2.585
cc_321 N_A_27_115#_M1015_g N_Y_c_522_n 0.00251111f $X=3.915 $Y=0.895 $X2=3.7
+ $Y2=2.585
cc_322 N_A_27_115#_c_353_n N_Y_c_522_n 0.0031083f $X=3.915 $Y=2.75 $X2=3.7
+ $Y2=2.585
cc_323 N_A_27_115#_c_305_n N_Y_c_522_n 6.99501e-19 $X=3.485 $Y=2.675 $X2=3.7
+ $Y2=2.585
