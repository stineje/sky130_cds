* File: sky130_osu_sc_12T_ms__nor2_l.pxi.spice
* Created: Fri Nov 12 15:25:37 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__NOR2_L%GND N_GND_M1003_s N_GND_M1001_d N_GND_M1003_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_12_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_MS__NOR2_L%GND
x_PM_SKY130_OSU_SC_12T_MS__NOR2_L%VDD N_VDD_M1000_d N_VDD_M1002_b N_VDD_c_28_p
+ N_VDD_c_34_p VDD N_VDD_c_29_p PM_SKY130_OSU_SC_12T_MS__NOR2_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__NOR2_L%B N_B_M1003_g N_B_M1002_g N_B_c_49_n
+ N_B_c_50_n N_B_c_51_n B PM_SKY130_OSU_SC_12T_MS__NOR2_L%B
x_PM_SKY130_OSU_SC_12T_MS__NOR2_L%A N_A_M1000_g N_A_M1001_g N_A_c_95_n
+ N_A_c_96_n A PM_SKY130_OSU_SC_12T_MS__NOR2_L%A
x_PM_SKY130_OSU_SC_12T_MS__NOR2_L%Y N_Y_M1003_d N_Y_M1002_s N_Y_c_122_n
+ N_Y_c_123_n Y N_Y_c_127_n N_Y_c_129_n N_Y_c_130_n N_Y_c_131_n
+ PM_SKY130_OSU_SC_12T_MS__NOR2_L%Y
cc_1 N_GND_M1003_b N_B_M1003_g 0.0747024f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.755
cc_2 N_GND_c_2_p N_B_M1003_g 0.00502587f $X=0.26 $Y=0.74 $X2=0.475 $Y2=0.755
cc_3 N_GND_c_3_p N_B_M1003_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.755
cc_4 N_GND_c_4_p N_B_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.755
cc_5 N_GND_M1003_b N_B_M1002_g 0.0410185f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.445
cc_6 N_GND_M1003_b N_B_c_49_n 0.0335172f $X=-0.045 $Y=0 $X2=0.415 $Y2=1.98
cc_7 N_GND_M1003_b N_B_c_50_n 0.00746714f $X=-0.045 $Y=0 $X2=0.565 $Y2=1.98
cc_8 N_GND_M1003_b N_B_c_51_n 0.0109743f $X=-0.045 $Y=0 $X2=0.65 $Y2=2.85
cc_9 N_GND_M1003_b B 0.00104324f $X=-0.045 $Y=0 $X2=0.65 $Y2=2.85
cc_10 N_GND_M1003_b N_A_M1001_g 0.134163f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.755
cc_11 N_GND_c_3_p N_A_M1001_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.755
cc_12 N_GND_c_12_p N_A_M1001_g 0.00502587f $X=1.12 $Y=0.74 $X2=0.905 $Y2=0.755
cc_13 N_GND_c_4_p N_A_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=0.755
cc_14 N_GND_M1003_b N_A_c_95_n 0.0375985f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.645
cc_15 N_GND_M1003_b N_A_c_96_n 0.00230061f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.48
cc_16 N_GND_M1003_b A 0.0185053f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.48
cc_17 N_GND_M1003_b N_Y_c_122_n 0.0154673f $X=-0.045 $Y=0 $X2=0.26 $Y2=2.48
cc_18 N_GND_M1003_b N_Y_c_123_n 0.0171459f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.74
cc_19 N_GND_c_3_p N_Y_c_123_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.74
cc_20 N_GND_c_4_p N_Y_c_123_n 0.00475776f $X=1.02 $Y=0.19 $X2=0.69 $Y2=0.74
cc_21 N_GND_M1003_b Y 0.040849f $X=-0.045 $Y=0 $X2=0.24 $Y2=1.685
cc_22 N_GND_M1003_b N_Y_c_127_n 0.00938169f $X=-0.045 $Y=0 $X2=0.345 $Y2=1.367
cc_23 N_GND_c_2_p N_Y_c_127_n 0.00832556f $X=0.26 $Y=0.74 $X2=0.345 $Y2=1.367
cc_24 N_GND_M1003_b N_Y_c_129_n 0.0154549f $X=-0.045 $Y=0 $X2=0.26 $Y2=2.48
cc_25 N_GND_M1003_b N_Y_c_130_n 0.0094923f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.37
cc_26 N_GND_M1003_b N_Y_c_131_n 0.00248521f $X=-0.045 $Y=0 $X2=0.545 $Y2=1.37
cc_27 N_VDD_M1002_b N_B_M1002_g 0.0273074f $X=-0.045 $Y=2.795 $X2=0.475
+ $Y2=3.445
cc_28 N_VDD_c_28_p N_B_M1002_g 0.00606474f $X=0.965 $Y=4.287 $X2=0.475 $Y2=3.445
cc_29 N_VDD_c_29_p N_B_M1002_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.445
cc_30 N_VDD_M1002_b N_B_c_51_n 0.00525583f $X=-0.045 $Y=2.795 $X2=0.65 $Y2=2.85
cc_31 N_VDD_M1002_b B 0.00896612f $X=-0.045 $Y=2.795 $X2=0.65 $Y2=2.85
cc_32 N_VDD_M1002_b N_A_M1000_g 0.0269579f $X=-0.045 $Y=2.795 $X2=0.835
+ $Y2=3.445
cc_33 N_VDD_c_28_p N_A_M1000_g 0.00606474f $X=0.965 $Y=4.287 $X2=0.835 $Y2=3.445
cc_34 N_VDD_c_34_p N_A_M1000_g 0.00713292f $X=1.05 $Y=3.275 $X2=0.835 $Y2=3.445
cc_35 N_VDD_c_29_p N_A_M1000_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.835 $Y2=3.445
cc_36 N_VDD_M1002_b N_A_c_95_n 0.00746821f $X=-0.045 $Y=2.795 $X2=0.99 $Y2=2.645
cc_37 N_VDD_c_34_p N_A_c_95_n 0.00298495f $X=1.05 $Y=3.275 $X2=0.99 $Y2=2.645
cc_38 N_VDD_M1002_b N_A_c_96_n 0.00323928f $X=-0.045 $Y=2.795 $X2=0.99 $Y2=2.48
cc_39 N_VDD_c_34_p N_A_c_96_n 0.00695908f $X=1.05 $Y=3.275 $X2=0.99 $Y2=2.48
cc_40 N_VDD_c_34_p A 0.0029636f $X=1.05 $Y=3.275 $X2=0.99 $Y2=2.48
cc_41 N_VDD_M1002_b N_Y_c_122_n 0.0121889f $X=-0.045 $Y=2.795 $X2=0.26 $Y2=2.48
cc_42 N_VDD_c_28_p N_Y_c_122_n 0.00736239f $X=0.965 $Y=4.287 $X2=0.26 $Y2=2.48
cc_43 N_VDD_c_29_p N_Y_c_122_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26 $Y2=2.48
cc_44 B N_A_M1000_g 0.00821593f $X=0.65 $Y=2.85 $X2=0.835 $Y2=3.445
cc_45 N_B_M1003_g N_A_M1001_g 0.0706022f $X=0.475 $Y=0.755 $X2=0.905 $Y2=0.755
cc_46 N_B_c_50_n N_A_M1001_g 0.00474266f $X=0.565 $Y=1.98 $X2=0.905 $Y2=0.755
cc_47 N_B_c_51_n N_A_M1001_g 0.00792155f $X=0.65 $Y=2.85 $X2=0.905 $Y2=0.755
cc_48 N_B_M1002_g N_A_c_95_n 0.0913308f $X=0.475 $Y=3.445 $X2=0.99 $Y2=2.645
cc_49 N_B_c_51_n N_A_c_95_n 0.00475824f $X=0.65 $Y=2.85 $X2=0.99 $Y2=2.645
cc_50 B N_A_c_95_n 0.00131279f $X=0.65 $Y=2.85 $X2=0.99 $Y2=2.645
cc_51 N_B_c_51_n N_A_c_96_n 0.0280464f $X=0.65 $Y=2.85 $X2=0.99 $Y2=2.48
cc_52 B N_A_c_96_n 0.00204062f $X=0.65 $Y=2.85 $X2=0.99 $Y2=2.48
cc_53 N_B_c_51_n A 0.00542135f $X=0.65 $Y=2.85 $X2=0.99 $Y2=2.48
cc_54 B A 0.00596751f $X=0.65 $Y=2.85 $X2=0.99 $Y2=2.48
cc_55 N_B_M1002_g N_Y_c_122_n 0.0167239f $X=0.475 $Y=3.445 $X2=0.26 $Y2=2.48
cc_56 N_B_c_49_n N_Y_c_122_n 0.00102058f $X=0.415 $Y=1.98 $X2=0.26 $Y2=2.48
cc_57 N_B_c_50_n N_Y_c_122_n 0.00330615f $X=0.565 $Y=1.98 $X2=0.26 $Y2=2.48
cc_58 N_B_c_51_n N_Y_c_122_n 0.0286186f $X=0.65 $Y=2.85 $X2=0.26 $Y2=2.48
cc_59 B N_Y_c_122_n 0.00819421f $X=0.65 $Y=2.85 $X2=0.26 $Y2=2.48
cc_60 N_B_M1003_g N_Y_c_123_n 0.0116832f $X=0.475 $Y=0.755 $X2=0.69 $Y2=0.74
cc_61 N_B_c_50_n N_Y_c_123_n 0.00364841f $X=0.565 $Y=1.98 $X2=0.69 $Y2=0.74
cc_62 N_B_M1003_g Y 0.00813678f $X=0.475 $Y=0.755 $X2=0.24 $Y2=1.685
cc_63 N_B_M1002_g Y 0.00514172f $X=0.475 $Y=3.445 $X2=0.24 $Y2=1.685
cc_64 N_B_c_49_n Y 0.00548589f $X=0.415 $Y=1.98 $X2=0.24 $Y2=1.685
cc_65 N_B_c_50_n Y 0.0141817f $X=0.565 $Y=1.98 $X2=0.24 $Y2=1.685
cc_66 N_B_c_51_n Y 0.0129003f $X=0.65 $Y=2.85 $X2=0.24 $Y2=1.685
cc_67 N_B_M1002_g N_Y_c_129_n 0.00399338f $X=0.475 $Y=3.445 $X2=0.26 $Y2=2.48
cc_68 N_B_c_49_n N_Y_c_129_n 0.00138163f $X=0.415 $Y=1.98 $X2=0.26 $Y2=2.48
cc_69 N_B_c_50_n N_Y_c_129_n 0.00227834f $X=0.565 $Y=1.98 $X2=0.26 $Y2=2.48
cc_70 N_B_c_51_n N_Y_c_129_n 0.00269535f $X=0.65 $Y=2.85 $X2=0.26 $Y2=2.48
cc_71 B N_Y_c_129_n 9.25684e-19 $X=0.65 $Y=2.85 $X2=0.26 $Y2=2.48
cc_72 N_B_M1003_g N_Y_c_130_n 0.0028533f $X=0.475 $Y=0.755 $X2=0.69 $Y2=1.37
cc_73 N_B_c_50_n N_Y_c_130_n 0.0057569f $X=0.565 $Y=1.98 $X2=0.69 $Y2=1.37
cc_74 N_B_M1003_g N_Y_c_131_n 0.010737f $X=0.475 $Y=0.755 $X2=0.545 $Y2=1.37
cc_75 N_B_c_49_n N_Y_c_131_n 0.00121385f $X=0.415 $Y=1.98 $X2=0.545 $Y2=1.37
cc_76 N_B_c_50_n N_Y_c_131_n 0.00589915f $X=0.565 $Y=1.98 $X2=0.545 $Y2=1.37
cc_77 N_A_M1001_g N_Y_c_123_n 0.0116832f $X=0.905 $Y=0.755 $X2=0.69 $Y2=0.74
cc_78 N_A_M1001_g Y 3.32097e-19 $X=0.905 $Y=0.755 $X2=0.24 $Y2=1.685
cc_79 A N_Y_c_129_n 0.0146886f $X=0.99 $Y=2.48 $X2=0.26 $Y2=2.48
cc_80 N_A_M1001_g N_Y_c_130_n 0.0110755f $X=0.905 $Y=0.755 $X2=0.69 $Y2=1.37
