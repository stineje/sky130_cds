magic
tech sky130A
magscale 1 2
timestamp 1606864609
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 375 1341
<< nmos >>
rect 80 115 110 263
rect 166 115 196 263
rect 238 115 268 263
<< pmos >>
rect 80 817 110 1217
rect 166 817 196 1217
rect 238 817 268 1217
<< ndiff >>
rect 27 199 80 263
rect 27 131 35 199
rect 69 131 80 199
rect 27 115 80 131
rect 110 199 166 263
rect 110 131 121 199
rect 155 131 166 199
rect 110 115 166 131
rect 196 115 238 263
rect 268 199 321 263
rect 268 131 279 199
rect 313 131 321 199
rect 268 115 321 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 861 35 1201
rect 69 861 80 1201
rect 27 817 80 861
rect 110 1201 166 1217
rect 110 861 121 1201
rect 155 861 166 1201
rect 110 817 166 861
rect 196 817 238 1217
rect 268 1201 321 1217
rect 268 861 279 1201
rect 313 861 321 1201
rect 268 817 321 861
<< ndiffc >>
rect 35 131 69 199
rect 121 131 155 199
rect 279 131 313 199
<< pdiffc >>
rect 35 861 69 1201
rect 121 861 155 1201
rect 279 861 313 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 238 1217 268 1243
rect 80 602 110 817
rect 39 572 110 602
rect 39 360 69 572
rect 166 529 196 817
rect 133 513 196 529
rect 133 479 143 513
rect 177 479 196 513
rect 133 463 196 479
rect 238 451 268 817
rect 238 435 292 451
rect 111 387 165 403
rect 111 360 121 387
rect 39 353 121 360
rect 155 360 165 387
rect 238 401 248 435
rect 282 401 292 435
rect 238 385 292 401
rect 155 353 196 360
rect 39 330 196 353
rect 80 263 110 330
rect 166 263 196 330
rect 238 263 268 385
rect 80 89 110 115
rect 166 89 196 115
rect 238 89 268 115
<< polycont >>
rect 143 479 177 513
rect 121 353 155 387
rect 248 401 282 435
<< locali >>
rect 0 1311 374 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 374 1311
rect 35 1201 69 1217
rect 35 513 69 861
rect 121 1201 155 1271
rect 121 845 155 861
rect 279 1201 313 1217
rect 143 513 177 529
rect 35 479 143 513
rect 35 199 69 479
rect 143 463 177 479
rect 211 435 245 649
rect 279 535 313 861
rect 211 401 248 435
rect 282 401 298 435
rect 103 353 121 387
rect 155 353 171 387
rect 35 115 69 131
rect 121 199 155 215
rect 121 61 155 131
rect 279 199 313 279
rect 279 115 313 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 211 649 245 683
rect 279 501 313 535
rect 121 353 155 387
rect 279 279 313 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 374 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 374 1311
rect 0 1271 374 1277
rect 199 683 257 689
rect 177 649 211 683
rect 245 649 257 683
rect 199 643 257 649
rect 109 609 167 615
rect 109 575 189 609
rect 109 569 167 575
rect 121 393 155 569
rect 267 535 325 541
rect 267 501 279 535
rect 313 501 325 535
rect 267 495 325 501
rect 109 387 167 393
rect 109 353 121 387
rect 155 353 167 387
rect 109 347 167 353
rect 279 319 313 495
rect 267 313 325 319
rect 267 279 279 313
rect 313 279 325 313
rect 267 273 325 279
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 305 364 305 364 1 Y
port 1 n
rlabel metal1 228 666 228 666 1 A
port 2 n
rlabel metal1 138 592 138 592 1 OE
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
