magic
tech sky130A
magscale 1 2
timestamp 1604007754
<< checkpaint >>
rect -1267 2461 1310 2601
rect -1760 -1129 6260 2461
rect -1267 -1260 1310 -1129
<< error_p >>
rect 0 1271 44 1332
rect 50 581 161 1341
rect 0 0 44 61
<< nwell >>
rect -7 529 50 1119
<< locali >>
rect 0 1049 44 1110
rect 0 0 44 61
<< metal1 >>
rect 0 1049 44 1110
rect 0 0 44 61
<< labels >>
rlabel metal1 23 28 23 28 1 gnd
rlabel metal1 22 1078 22 1078 1 vdd
<< end >>
