* File: sky130_osu_sc_12T_ls__aoi22_l.spice
* Created: Fri Nov 12 15:34:49 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__aoi22_l.pex.spice"
.subckt sky130_osu_sc_12T_ls__aoi22_l  GND VDD A0 A1 B0 B1 Y
* 
* Y	Y
* B1	B1
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1005 A_110_115# N_A0_M1005_g N_GND_M1005_s N_GND_M1005_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_110_115# N_GND_M1005_b NSHORT L=0.15 W=0.52
+ AD=0.091 AS=0.0546 PD=0.87 PS=0.73 NRD=8.076 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75001 A=0.078 P=1.34 MULT=1
MM1000 A_282_115# N_B0_M1000_g N_Y_M1001_d N_GND_M1005_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.091 PD=0.73 PS=0.87 NRD=11.532 NRS=8.076 M=1 R=3.46667 SA=75001
+ SB=75000.5 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_B1_M1007_g A_282_115# N_GND_M1005_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0546 PD=1.57 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1003 N_VDD_M1003_d N_A0_M1003_g N_A_27_521#_M1003_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_27_521#_M1006_d N_A1_M1006_g N_VDD_M1003_d N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_B0_M1004_g N_A_27_521#_M1006_d N_VDD_M1003_b PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1002 N_A_27_521#_M1002_d N_B1_M1002_g N_Y_M1004_d N_VDD_M1003_b PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1005_b N_VDD_M1003_b NWDIODE A=4.8513 P=8.83
pX9_noxref noxref_11 A0 A0 PROBETYPE=1
pX10_noxref noxref_12 A1 A1 PROBETYPE=1
pX11_noxref noxref_13 B0 B0 PROBETYPE=1
pX12_noxref noxref_14 Y Y PROBETYPE=1
pX13_noxref noxref_15 B1 B1 PROBETYPE=1
c_287 A_282_115# 0 5.84789e-20 $X=1.41 $Y=0.575
*
.include "sky130_osu_sc_12T_ls__aoi22_l.pxi.spice"
*
.ends
*
*
