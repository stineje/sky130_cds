* File: sky130_osu_sc_18T_ms__inv_6.pex.spice
* Created: Fri Nov 12 14:04:38 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__INV_6%GND 1 2 3 4 41 45 47 54 56 63 65 73 84 86
r82 84 86 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r83 71 73 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.825
r84 66 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r85 65 71 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.305
r86 61 80 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r87 61 63 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r88 57 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r89 56 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r90 52 79 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r91 52 54 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r92 47 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r93 43 45 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r94 41 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r95 41 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r96 41 43 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r97 41 48 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r98 41 65 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r99 41 66 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r100 41 56 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r101 41 57 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r102 41 47 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r103 41 48 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r104 4 73 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r105 3 63 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r106 2 54 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r107 1 45 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_6%VDD 1 2 3 4 33 37 41 47 51 57 61 68 78 82
r58 78 82 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=2.38 $Y2=6.507
r59 73 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r60 68 71 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r61 66 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.84 $Y2=5.835
r62 64 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=6.47
+ $X2=2.38 $Y2=6.47
r63 62 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=1.98 $Y2=6.507
r64 62 64 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=2.38 $Y2=6.507
r65 61 66 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.84 $Y2=6.355
r66 61 64 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.38 $Y2=6.507
r67 57 60 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r68 55 76 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=6.507
r69 55 60 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r70 52 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r71 52 54 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r72 51 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.98 $Y2=6.507
r73 51 54 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r74 47 50 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r75 45 75 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r76 45 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r77 42 73 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r78 42 44 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r79 41 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r80 41 44 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r81 37 40 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r82 35 73 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r83 35 40 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r84 33 64 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r85 33 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r86 33 44 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r87 33 73 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r88 4 71 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r89 4 68 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r90 3 60 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r91 3 57 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r92 2 50 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r93 2 47 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r94 1 40 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r95 1 37 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_6%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 45 47 49 50 52 53 55 57 59 60 62 63 65 66 68
+ 69 70 71 72 73 74 75 76 79 81 83 86
c179 50 0 1.33323e-19 $X=2.195 $Y=2.96
c180 45 0 1.33323e-19 $X=2.195 $Y=1.7
c181 38 0 1.33323e-19 $X=1.765 $Y=2.96
c182 35 0 1.33323e-19 $X=1.765 $Y=1.7
c183 28 0 1.33323e-19 $X=1.335 $Y=2.96
c184 25 0 1.33323e-19 $X=1.335 $Y=1.7
c185 18 0 1.33323e-19 $X=0.905 $Y=2.96
c186 15 0 1.33323e-19 $X=0.905 $Y=1.7
r187 86 89 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=3.325
+ $X2=0.405 $Y2=3.33
r188 81 83 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.305
+ $X2=0.535 $Y2=2.305
r189 79 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r190 77 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=2.39
+ $X2=0.405 $Y2=2.305
r191 77 79 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.39
+ $X2=0.32 $Y2=3.33
r192 65 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.305 $X2=0.535 $Y2=2.305
r193 65 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.47
r194 65 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.14
r195 60 62 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.625 $Y=2.96
+ $X2=2.625 $Y2=4.585
r196 57 59 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.625 $Y=1.7
+ $X2=2.625 $Y2=1.075
r197 56 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.885
+ $X2=2.195 $Y2=2.885
r198 55 60 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.625 $Y2=2.96
r199 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.27 $Y2=2.885
r200 54 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.775
+ $X2=2.195 $Y2=1.775
r201 53 57 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=1.775
+ $X2=2.625 $Y2=1.7
r202 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.775
+ $X2=2.27 $Y2=1.775
r203 50 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=2.885
r204 50 52 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=4.585
r205 49 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.81
+ $X2=2.195 $Y2=2.885
r206 48 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.85
+ $X2=2.195 $Y2=1.775
r207 48 49 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.85
+ $X2=2.195 $Y2=2.81
r208 45 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.7 $X2=2.195
+ $Y2=1.775
r209 45 47 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.195 $Y=1.7
+ $X2=2.195 $Y2=1.075
r210 44 74 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.885
+ $X2=1.765 $Y2=2.885
r211 43 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=2.195 $Y2=2.885
r212 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=1.84 $Y2=2.885
r213 42 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.775
+ $X2=1.765 $Y2=1.775
r214 41 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.775
+ $X2=2.195 $Y2=1.775
r215 41 42 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.775
+ $X2=1.84 $Y2=1.775
r216 38 74 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=2.885
r217 38 40 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r218 35 73 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.7
+ $X2=1.765 $Y2=1.775
r219 35 37 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.765 $Y=1.7
+ $X2=1.765 $Y2=1.075
r220 34 72 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.885
+ $X2=1.335 $Y2=2.885
r221 33 74 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.885
r222 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.41 $Y2=2.885
r223 32 71 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.775
+ $X2=1.335 $Y2=1.775
r224 31 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.775
+ $X2=1.765 $Y2=1.775
r225 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.775
+ $X2=1.41 $Y2=1.775
r226 28 72 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=2.885
r227 28 30 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r228 25 71 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.7
+ $X2=1.335 $Y2=1.775
r229 25 27 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.335 $Y=1.7
+ $X2=1.335 $Y2=1.075
r230 24 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.885
+ $X2=0.905 $Y2=2.885
r231 23 72 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=1.335 $Y2=2.885
r232 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=0.98 $Y2=2.885
r233 22 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.775
+ $X2=0.905 $Y2=1.775
r234 21 71 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=1.335 $Y2=1.775
r235 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=0.98 $Y2=1.775
r236 18 70 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=2.885
r237 18 20 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=4.585
r238 15 69 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.775
r239 15 17 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.075
r240 14 68 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.885
+ $X2=0.475 $Y2=2.885
r241 13 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.905 $Y2=2.885
r242 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.55 $Y2=2.885
r243 12 63 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.775
+ $X2=0.475 $Y2=1.775
r244 11 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.905 $Y2=1.775
r245 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.55 $Y2=1.775
r246 8 68 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=2.885
r247 8 10 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=4.585
r248 7 68 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.885
r249 7 67 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.47
r250 4 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=1.775
r251 4 66 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=2.14
r252 1 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.775
r253 1 3 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_6%Y 1 2 3 7 8 9 26 32 40 46 54 60 67 68 70
+ 72 74 77 78 79 80 81 82 83
c129 83 0 1.33323e-19 $X=2.41 $Y=2.845
c130 82 0 1.33323e-19 $X=2.41 $Y=1.595
c131 81 0 2.66647e-19 $X=1.695 $Y=2.96
c132 79 0 2.66647e-19 $X=1.695 $Y=1.48
c133 68 0 1.33323e-19 $X=0.69 $Y=2.845
c134 67 0 1.33323e-19 $X=0.69 $Y=1.595
r135 83 95 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.845
+ $X2=2.41 $Y2=2.96
r136 82 93 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=1.48
r137 82 83 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=2.845
r138 81 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.96
+ $X2=1.55 $Y2=2.96
r139 80 95 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.96
+ $X2=2.41 $Y2=2.96
r140 80 81 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.96
+ $X2=1.695 $Y2=2.96
r141 79 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.48
+ $X2=1.55 $Y2=1.48
r142 78 93 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=2.41 $Y2=1.48
r143 78 79 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=1.695 $Y2=1.48
r144 77 91 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.845
+ $X2=1.55 $Y2=2.96
r145 76 89 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r146 76 77 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.845
r147 75 87 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.96
+ $X2=0.69 $Y2=2.96
r148 74 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=1.55 $Y2=2.96
r149 74 75 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=0.835 $Y2=2.96
r150 73 85 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.48
+ $X2=0.69 $Y2=1.48
r151 72 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=1.55 $Y2=1.48
r152 72 73 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=0.835 $Y2=1.48
r153 68 87 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.96
r154 68 70 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.2
r155 67 85 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.48
r156 67 70 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=2.2
r157 63 65 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r158 60 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.96
+ $X2=2.41 $Y2=2.96
r159 60 63 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.41 $Y=2.96
+ $X2=2.41 $Y2=3.455
r160 57 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.48
+ $X2=2.41 $Y2=1.48
r161 54 57 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.41 $Y=0.825
+ $X2=2.41 $Y2=1.48
r162 49 51 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r163 46 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=2.96
r164 46 49 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=3.455
r165 43 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r166 40 43 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r167 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r168 32 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=2.96
r169 32 35 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=3.455
r170 29 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.48
r171 26 29 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.69 $Y=0.825
+ $X2=0.69 $Y2=1.48
r172 9 65 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r173 9 63 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r174 8 51 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r175 8 49 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r176 7 37 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r177 7 35 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r178 3 54 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r179 2 40 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r180 1 26 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

