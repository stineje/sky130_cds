* File: sky130_osu_sc_12T_hs__and2_2.pex.spice
* Created: Fri Nov 12 15:06:52 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__AND2_2%GND 1 2 27 29 37 39 47 55 57
r44 55 57 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r45 45 47 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r46 39 45 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.305
r47 35 37 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.755
r48 27 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r49 27 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r50 27 35 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r51 27 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r52 27 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r53 27 39 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r54 27 40 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r55 27 29 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r56 2 47 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84 $Y=0.575
+ $X2=1.98 $Y2=0.755
r57 1 37 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.91 $Y=0.575
+ $X2=1.05 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__AND2_2%VDD 1 2 3 25 29 31 37 39 46 55 59
r36 55 59 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.7 $Y2=4.287
r37 51 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r38 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r39 44 49 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135 $X2=1.98
+ $Y2=3.635
r40 42 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=4.25 $X2=1.7
+ $Y2=4.25
r41 40 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r42 40 42 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r43 39 44 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.135
r44 39 42 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r45 35 53 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r46 35 37 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.295
r47 32 51 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r48 32 34 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r49 31 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r50 31 34 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r51 27 51 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r52 27 29 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135 $X2=0.26
+ $Y2=3.635
r53 25 42 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r54 25 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r55 25 51 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r56 3 49 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r57 3 46 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r58 2 37 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.295
r59 1 29 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__AND2_2%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=2.85
+ $X2=0.275 $Y2=2.85
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.85
+ $X2=0.27 $Y2=2.85
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.285
+ $X2=0.27 $Y2=2.85
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.285 $X2=0.27 $Y2=2.285
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.285
+ $X2=0.475 $Y2=2.285
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.45
+ $X2=0.475 $Y2=2.285
r38 5 7 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.475 $Y=2.45
+ $X2=0.475 $Y2=3.235
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=2.285
r40 1 3 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=0.85
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__AND2_2%B 3 7 10 14 22
c41 7 0 1.37149e-19 $X=0.905 $Y=3.235
r42 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.48
+ $X2=0.955 $Y2=2.48
r43 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.48
+ $X2=0.95 $Y2=2.48
r44 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=1.945
+ $X2=0.95 $Y2=2.48
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.945 $X2=0.95 $Y2=1.945
r46 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=1.945
+ $X2=0.922 $Y2=2.11
r47 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=1.945
+ $X2=0.922 $Y2=1.78
r48 7 12 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.11
r49 3 11 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.835 $Y=0.85
+ $X2=0.835 $Y2=1.78
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__AND2_2%A_27_115# 1 3 11 13 15 17 18 22 24 26 27
+ 31 35 37 38 43 47 49 50 51
r87 50 51 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.065
+ $X2=0.65 $Y2=3.235
r88 45 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.455
+ $X2=0.61 $Y2=1.455
r89 45 47 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.455
+ $X2=1.43 $Y2=1.455
r90 43 51 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.69 $Y=3.295 $X2=0.69
+ $Y2=3.235
r91 39 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.54 $X2=0.61
+ $Y2=1.455
r92 39 50 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=3.065
r93 37 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.455
+ $X2=0.61 $Y2=1.455
r94 37 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.455
+ $X2=0.345 $Y2=1.455
r95 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.345 $Y2=1.455
r96 33 35 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r97 31 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.455 $X2=1.43 $Y2=1.455
r98 29 31 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.455 $X2=1.43
+ $Y2=1.455
r99 28 29 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.455
+ $X2=1.37 $Y2=1.455
r100 24 26 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r101 20 31 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.43 $Y2=1.455
r102 20 22 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=0.85
r103 19 27 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.405
+ $X2=1.352 $Y2=2.405
r104 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.48
r105 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.445 $Y2=2.405
r106 17 27 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.33
+ $X2=1.352 $Y2=2.405
r107 16 29 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=1.455
r108 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=2.33
r109 13 27 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.352 $Y2=2.405
r110 13 15 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r111 9 28 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=1.455
r112 9 11 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.85
r113 3 43 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.295
r114 1 35 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__AND2_2%Y 1 3 10 16 26 29 32
c42 16 0 1.37149e-19 $X=1.55 $Y=2.11
r43 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=2.11
r44 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=1.74
r45 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r46 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.74
r47 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r48 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.11
r49 16 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.955
r50 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r51 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r52 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r53 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r54 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41 $Y=0.575
+ $X2=1.55 $Y2=0.755
.ends

