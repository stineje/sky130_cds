magic
tech sky130A
magscale 1 2
timestamp 1606864598
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 374 1341
<< nmos >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
<< pmoshvt >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 166 315
rect 110 131 121 267
rect 155 131 166 267
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 267 335 315
rect 282 131 293 267
rect 327 131 335 267
rect 282 115 335 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 725 35 1201
rect 69 725 80 1201
rect 27 617 80 725
rect 110 617 166 1217
rect 196 1201 252 1217
rect 196 793 207 1201
rect 241 793 252 1201
rect 196 617 252 793
rect 282 1201 335 1217
rect 282 657 293 1201
rect 327 657 335 1201
rect 282 617 335 657
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 207 131 241 267
rect 293 131 327 267
<< pdiffc >>
rect 35 725 69 1201
rect 207 793 241 1201
rect 293 657 327 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 80 568 110 617
rect 27 552 110 568
rect 27 518 37 552
rect 71 518 110 552
rect 27 502 110 518
rect 166 510 196 617
rect 252 592 282 617
rect 252 562 289 592
rect 80 315 110 502
rect 163 494 217 510
rect 163 460 173 494
rect 207 460 217 494
rect 163 444 217 460
rect 166 315 196 444
rect 259 420 289 562
rect 259 404 313 420
rect 259 384 269 404
rect 252 370 269 384
rect 303 370 313 404
rect 252 354 313 370
rect 252 315 282 354
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
<< polycont >>
rect 37 518 71 552
rect 173 460 207 494
rect 269 370 303 404
<< locali >>
rect 0 1311 374 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 374 1311
rect 35 1201 69 1217
rect 207 1201 241 1271
rect 207 777 241 793
rect 293 1201 327 1217
rect 69 725 139 743
rect 35 709 139 725
rect 37 552 71 575
rect 37 502 71 518
rect 105 404 139 709
rect 173 494 207 649
rect 293 535 327 657
rect 173 444 207 460
rect 105 370 269 404
rect 303 370 319 404
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 370
rect 121 115 155 131
rect 207 267 241 283
rect 207 61 241 131
rect 293 267 327 279
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 37 575 71 609
rect 173 649 207 683
rect 293 501 327 535
rect 293 279 327 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 374 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 374 1311
rect 0 1271 374 1277
rect 161 683 219 689
rect 140 649 173 683
rect 207 649 219 683
rect 161 643 219 649
rect 25 609 83 615
rect 25 575 37 609
rect 71 575 105 609
rect 25 569 83 575
rect 281 535 339 541
rect 281 501 293 535
rect 327 501 339 535
rect 281 495 339 501
rect 293 319 327 495
rect 281 313 339 319
rect 281 279 293 313
rect 327 279 339 313
rect 281 273 339 279
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 311 444 311 444 1 Y
port 1 n
rlabel metal1 190 666 190 666 1 A
port 2 n
rlabel metal1 54 592 54 592 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
