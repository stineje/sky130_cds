* File: sky130_osu_sc_18T_ls__xnor2_l.pex.spice
* Created: Fri Nov 12 14:20:42 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%GND 1 2 33 35 43 45 55 67 69
r69 67 69 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r70 53 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.825
r71 46 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r72 41 59 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r73 41 43 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r74 35 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r75 33 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r76 33 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r77 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r78 33 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r79 33 45 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r80 33 46 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r81 33 35 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r82 2 55 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.575 $X2=2.44 $Y2=0.825
r83 1 43 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%VDD 1 2 25 27 34 38 46 54 57 61
c40 34 0 1.59951e-19 $X=0.69 $Y=3.455
r41 57 61 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=2.38 $Y2=6.507
r42 54 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=6.47
+ $X2=2.38 $Y2=6.47
r43 46 49 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.44 $Y=3.455
+ $X2=2.44 $Y2=5.835
r44 44 54 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=6.355
+ $X2=2.44 $Y2=6.507
r45 44 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.44 $Y=6.355
+ $X2=2.44 $Y2=5.835
r46 41 43 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r47 39 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r48 39 41 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r49 38 54 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=6.507
+ $X2=2.44 $Y2=6.507
r50 38 43 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=6.507
+ $X2=1.7 $Y2=6.507
r51 34 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r52 32 52 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r53 32 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r54 29 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r55 27 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r56 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r57 25 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r58 25 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r59 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r60 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r61 2 49 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.3
+ $Y=3.085 $X2=2.44 $Y2=5.835
r62 2 46 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.3
+ $Y=3.085 $X2=2.44 $Y2=3.455
r63 1 37 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r64 1 34 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%A 3 5 8 9 13 16 18 19 20 21 22 26 30 37
+ 42 44 45 50 53
r114 47 50 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=0.845 $Y=1.48
+ $X2=0.85 $Y2=1.48
r115 45 50 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=0.99 $Y=1.48
+ $X2=0.85 $Y2=1.48
r116 44 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2 $Y=1.48
+ $X2=2.145 $Y2=1.48
r117 44 45 0.972511 $w=1.7e-07 $l=1.01e-06 $layer=MET1_cond $X=2 $Y=1.48
+ $X2=0.99 $Y2=1.48
r118 39 42 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.145 $Y=2.39
+ $X2=2.225 $Y2=2.39
r119 37 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=1.48
+ $X2=2.145 $Y2=1.48
r120 35 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.305
+ $X2=2.145 $Y2=2.39
r121 35 37 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.145 $Y=2.305
+ $X2=2.145 $Y2=1.48
r122 30 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.845 $Y=1.48
+ $X2=0.845 $Y2=1.48
r123 30 33 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.845 $Y=1.48
+ $X2=0.845 $Y2=1.85
r124 28 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=2.39 $X2=2.225 $Y2=2.39
r125 26 28 73.8383 $w=2.35e-07 $l=3.6e-07 $layer=POLY_cond $X=1.865 $Y=2.405
+ $X2=2.225 $Y2=2.405
r126 24 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.85 $X2=0.845 $Y2=1.85
r127 21 24 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=0.845 $Y=1.725
+ $X2=0.845 $Y2=1.85
r128 21 22 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.725
+ $X2=0.845 $Y2=1.65
r129 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.45 $Y=2.86 $X2=0.45
+ $Y2=3.01
r130 14 26 13.2911 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.865 $Y=2.555
+ $X2=1.865 $Y2=2.405
r131 14 16 1040.91 $w=1.5e-07 $l=2.03e-06 $layer=POLY_cond $X=1.865 $Y=2.555
+ $X2=1.865 $Y2=4.585
r132 13 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=1.65
r133 10 18 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=1.725
+ $X2=0.45 $Y2=1.725
r134 9 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=1.725
+ $X2=0.845 $Y2=1.725
r135 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=1.725
+ $X2=0.55 $Y2=1.725
r136 8 20 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=3.01
r137 3 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.45 $Y2=1.725
r138 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.65
+ $X2=0.475 $Y2=1.075
r139 1 18 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=1.8
+ $X2=0.45 $Y2=1.725
r140 1 19 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.425 $Y=1.8
+ $X2=0.425 $Y2=2.86
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%A_27_115# 1 3 11 13 15 17 21 25 29 33
+ 39 41
c78 39 0 1.07013e-19 $X=1.765 $Y=1.85
r79 37 39 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.765 $Y=2.305
+ $X2=1.765 $Y2=1.85
r80 34 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.39
+ $X2=0.26 $Y2=2.39
r81 34 36 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=2.39
+ $X2=0.845 $Y2=2.39
r82 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=2.39
+ $X2=1.765 $Y2=2.305
r83 33 36 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.68 $Y=2.39
+ $X2=0.845 $Y2=2.39
r84 29 31 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r85 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.475
+ $X2=0.26 $Y2=2.39
r86 27 29 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.26 $Y=2.475
+ $X2=0.26 $Y2=3.455
r87 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.305
+ $X2=0.26 $Y2=2.39
r88 23 25 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.26 $Y=2.305
+ $X2=0.26 $Y2=0.825
r89 21 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.85 $X2=1.765 $Y2=1.85
r90 21 22 15.9603 $w=3.02e-07 $l=1e-07 $layer=POLY_cond $X=1.765 $Y=1.85
+ $X2=1.865 $Y2=1.85
r91 17 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.39 $X2=0.845 $Y2=2.39
r92 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=2.39
+ $X2=0.845 $Y2=2.555
r93 13 22 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.685
+ $X2=1.865 $Y2=1.85
r94 13 15 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.865 $Y=1.685
+ $X2=1.865 $Y2=1.075
r95 11 19 1040.91 $w=1.5e-07 $l=2.03e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.555
r96 3 31 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r97 3 29 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r98 1 25 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%A_238_89# 1 3 11 15 18 21 27 31 35
r60 31 33 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.87 $Y=3.455
+ $X2=2.87 $Y2=5.835
r61 29 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.85 $X2=2.87
+ $Y2=2.765
r62 29 31 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.87 $Y=2.85
+ $X2=2.87 $Y2=3.455
r63 25 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.68 $X2=2.87
+ $Y2=2.765
r64 25 27 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=2.87 $Y=2.68
+ $X2=2.87 $Y2=0.825
r65 21 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=2.765
+ $X2=2.87 $Y2=2.765
r66 21 23 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=2.765
+ $X2=1.325 $Y2=2.765
r67 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.765 $X2=1.325 $Y2=2.765
r68 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.765
+ $X2=1.325 $Y2=2.93
r69 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.765
+ $X2=1.325 $Y2=2.6
r70 15 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.265 $Y=4.585
+ $X2=1.265 $Y2=2.93
r71 11 19 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=1.265 $Y=1.075
+ $X2=1.265 $Y2=2.6
r72 3 33 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.73
+ $Y=3.085 $X2=2.87 $Y2=5.835
r73 3 31 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.73
+ $Y=3.085 $X2=2.87 $Y2=3.455
r74 1 27 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.73
+ $Y=0.575 $X2=2.87 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 20 21 23 28
c56 20 0 1.07013e-19 $X=2.655 $Y=1.832
r57 23 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.85
+ $X2=2.53 $Y2=1.85
r58 19 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.85 $X2=2.53 $Y2=1.85
r59 19 20 21.9891 $w=2.74e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=1.832
+ $X2=2.655 $Y2=1.832
r60 14 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=3.01
+ $X2=2.655 $Y2=2.935
r61 14 16 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.655 $Y=3.01
+ $X2=2.655 $Y2=4.585
r62 13 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=2.86
+ $X2=2.655 $Y2=2.935
r63 12 20 16.847 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=2.655 $Y=2.015
+ $X2=2.655 $Y2=1.832
r64 12 13 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=2.655 $Y=2.015
+ $X2=2.655 $Y2=2.86
r65 9 20 16.847 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.832
r66 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.075
r67 7 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=2.935
+ $X2=2.655 $Y2=2.935
r68 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=2.935 $X2=2.3
+ $Y2=2.935
r69 4 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=3.01
+ $X2=2.3 $Y2=2.935
r70 4 6 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.225 $Y=3.01
+ $X2=2.225 $Y2=4.585
r71 1 19 53.6533 $w=2.74e-07 $l=3.85402e-07 $layer=POLY_cond $X=2.225 $Y=1.65
+ $X2=2.53 $Y2=1.832
r72 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.225 $Y=1.65
+ $X2=2.225 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XNOR2_L%Y 1 3 11 15 17 19 24 30 33 36
c56 30 0 1.59951e-19 $X=1.42 $Y=2.135
r57 28 36 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=3.215
+ $X2=1.425 $Y2=3.33
r58 28 30 1.03991 $w=1.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.425 $Y=3.215
+ $X2=1.425 $Y2=2.135
r59 27 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.965
+ $X2=1.425 $Y2=1.85
r60 27 30 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.425 $Y=1.965
+ $X2=1.425 $Y2=2.135
r61 26 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=3.33
+ $X2=1.425 $Y2=3.33
r62 23 24 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.537 $Y=1.245
+ $X2=1.537 $Y2=1.415
r63 19 21 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.565 $Y=3.455
+ $X2=1.565 $Y2=5.835
r64 17 26 3.84112 $w=3.85e-07 $l=1.28238e-07 $layer=LI1_cond $X=1.565 $Y=3.445
+ $X2=1.537 $Y2=3.33
r65 17 19 0.338954 $w=3.38e-07 $l=1e-08 $layer=LI1_cond $X=1.565 $Y=3.445
+ $X2=1.565 $Y2=3.455
r66 15 23 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.565 $Y=0.825
+ $X2=1.565 $Y2=1.245
r67 11 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=1.85
+ $X2=1.425 $Y2=1.85
r68 11 24 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.425 $Y=1.85
+ $X2=1.425 $Y2=1.415
r69 3 21 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.565 $Y2=5.835
r70 3 19 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.565 $Y2=3.455
r71 1 15 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.825
.ends

