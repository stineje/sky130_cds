magic
tech sky130A
magscale 1 2
timestamp 1612372309
<< nwell >>
rect -9 529 199 1119
<< nmoslvt >>
rect 80 115 110 243
<< pmos >>
rect 80 837 110 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 163 243
rect 110 131 121 215
rect 155 131 163 215
rect 110 115 163 131
<< pdiff >>
rect 27 949 80 965
rect 27 865 35 949
rect 69 865 80 949
rect 27 837 80 865
rect 110 949 163 965
rect 110 865 121 949
rect 155 865 163 949
rect 110 837 163 865
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
<< pdiffc >>
rect 35 865 69 949
rect 121 865 155 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1049 85 1083
<< poly >>
rect 80 965 110 991
rect 80 243 110 837
rect 80 80 110 115
<< locali >>
rect 0 1089 198 1110
rect 0 1049 51 1089
rect 85 1049 198 1089
rect 35 949 69 1049
rect 35 849 69 865
rect 121 949 155 1049
rect 121 849 155 865
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 231
rect 121 61 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1089 198 1110
rect 0 1055 51 1089
rect 85 1055 198 1089
rect 0 1049 198 1055
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
