* File: sky130_osu_sc_15T_hs__addf_1.spice
* Created: Fri Nov 12 14:26:08 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__addf_1.pex.spice"
.subckt sky130_osu_sc_15T_hs__addf_1  GND VDD A B CI CON S CO
* 
* CO	CO
* S	S
* CON	CON
* CI	CI
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1010 N_GND_M1010_d N_A_M1010_g N_A_27_115#_M1010_s N_GND_M1010_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005.3 A=0.096 P=1.58 MULT=1
MM1001 N_A_27_115#_M1001_d N_B_M1001_g N_GND_M1010_d N_GND_M1010_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75004.9 A=0.096 P=1.58 MULT=1
MM1003 N_CON_M1003_d N_CI_M1003_g N_A_27_115#_M1001_d N_GND_M1010_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75004.4 A=0.096 P=1.58 MULT=1
MM1023 A_368_115# N_B_M1023_g N_CON_M1003_d N_GND_M1010_b NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75004 A=0.096 P=1.58 MULT=1
MM1026 N_GND_M1026_d N_A_M1026_g A_368_115# N_GND_M1010_b NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75001.8
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1018 N_A_526_115#_M1018_d N_A_M1018_g N_GND_M1026_d N_GND_M1010_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1022 N_GND_M1022_d N_B_M1022_g N_A_526_115#_M1018_d N_GND_M1010_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.7 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1011 N_A_526_115#_M1011_d N_CI_M1011_g N_GND_M1022_d N_GND_M1010_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.1 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1012 N_A_784_115#_M1012_d N_CON_M1012_g N_A_526_115#_M1011_d N_GND_M1010_b
+ NLOWVT L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75003.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 A_870_115# N_B_M1013_g N_A_784_115#_M1012_d N_GND_M1010_b NLOWVT L=0.15
+ W=0.64 AD=0.0832 AS=0.0896 PD=0.9 PS=0.92 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75004 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 A_952_115# N_CI_M1005_g A_870_115# N_GND_M1010_b NLOWVT L=0.15 W=0.64
+ AD=0.0832 AS=0.0832 PD=0.9 PS=0.9 NRD=14.052 NRS=14.052 M=1 R=4.26667
+ SA=75004.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_GND_M1004_d N_A_M1004_g A_952_115# N_GND_M1010_b NLOWVT L=0.15 W=0.64
+ AD=0.1088 AS=0.0832 PD=0.98 PS=0.9 NRD=0 NRS=14.052 M=1 R=4.26667 SA=75004.8
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1014 N_S_M1014_d N_A_784_115#_M1014_g N_GND_M1004_d N_GND_M1010_b NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1088 PD=1.81 PS=0.98 NRD=0 NRS=11.244 M=1
+ R=4.26667 SA=75005.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 N_CO_M1019_d N_CON_M1019_g N_GND_M1019_s N_GND_M1010_b NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VDD_M1015_d N_A_M1015_g N_A_27_565#_M1015_s N_VDD_M1015_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75005.3 A=0.3 P=4.3 MULT=1
MM1006 N_A_27_565#_M1006_d N_B_M1006_g N_VDD_M1015_d N_VDD_M1015_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75004.9 A=0.3 P=4.3 MULT=1
MM1008 N_CON_M1008_d N_CI_M1008_g N_A_27_565#_M1006_d N_VDD_M1015_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75004.4 A=0.3 P=4.3 MULT=1
MM1000 A_368_565# N_B_M1000_g N_CON_M1008_d N_VDD_M1015_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75001.5
+ SB=75004 A=0.3 P=4.3 MULT=1
MM1002 N_VDD_M1002_d N_A_M1002_g A_368_565# N_VDD_M1015_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001.8
+ SB=75003.6 A=0.3 P=4.3 MULT=1
MM1024 N_A_526_565#_M1024_d N_A_M1024_g N_VDD_M1002_d N_VDD_M1015_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.3 SB=75003.2 A=0.3 P=4.3 MULT=1
MM1027 N_VDD_M1027_d N_B_M1027_g N_A_526_565#_M1024_d N_VDD_M1015_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.7 SB=75002.8 A=0.3 P=4.3 MULT=1
MM1016 N_A_526_565#_M1016_d N_CI_M1016_g N_VDD_M1027_d N_VDD_M1015_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.1 SB=75002.4 A=0.3 P=4.3 MULT=1
MM1017 N_A_784_115#_M1017_d N_CON_M1017_g N_A_526_565#_M1016_d N_VDD_M1015_b
+ PSHORT L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.6 SB=75001.9 A=0.3 P=4.3 MULT=1
MM1020 A_870_565# N_B_M1020_g N_A_784_115#_M1017_d N_VDD_M1015_b PSHORT L=0.15
+ W=2 AD=0.26 AS=0.28 PD=2.26 PS=2.28 NRD=7.3678 NRS=0 M=1 R=13.3333 SA=75004
+ SB=75001.5 A=0.3 P=4.3 MULT=1
MM1009 A_952_565# N_CI_M1009_g A_870_565# N_VDD_M1015_b PSHORT L=0.15 W=2
+ AD=0.26 AS=0.26 PD=2.26 PS=2.26 NRD=7.3678 NRS=7.3678 M=1 R=13.3333 SA=75004.4
+ SB=75001.1 A=0.3 P=4.3 MULT=1
MM1007 N_VDD_M1007_d N_A_M1007_g A_952_565# N_VDD_M1015_b PSHORT L=0.15 W=2
+ AD=0.34 AS=0.26 PD=2.34 PS=2.26 NRD=0 NRS=7.3678 M=1 R=13.3333 SA=75004.8
+ SB=75000.7 A=0.3 P=4.3 MULT=1
MM1021 N_S_M1021_d N_A_784_115#_M1021_g N_VDD_M1007_d N_VDD_M1015_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.34 PD=4.53 PS=2.34 NRD=0 NRS=5.8903 M=1 R=13.3333
+ SA=75005.3 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1025 N_CO_M1025_d N_CON_M1025_g N_VDD_M1025_s N_VDD_M1015_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX28_noxref N_GND_M1010_b N_VDD_M1015_b NWDIODE A=21.299 P=20.34
pX29_noxref noxref_20 A A PROBETYPE=1
pX30_noxref noxref_21 B B PROBETYPE=1
pX31_noxref noxref_22 CI CI PROBETYPE=1
pX32_noxref noxref_23 S S PROBETYPE=1
pX33_noxref noxref_24 CON CON PROBETYPE=1
pX34_noxref noxref_25 CO CO PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__addf_1.pxi.spice"
*
.ends
*
*
