magic
tech sky130A
magscale 1 2
timestamp 1606864594
<< checkpaint >>
rect -1210 -1243 2840 2575
<< nwell >>
rect -10 581 1741 1341
<< nmos >>
rect 80 115 110 263
rect 152 115 182 263
rect 356 115 386 315
rect 428 115 458 315
rect 548 115 578 315
rect 620 115 650 315
rect 706 115 736 315
rect 778 115 808 315
rect 898 115 928 315
rect 970 115 1000 315
rect 1056 115 1086 315
rect 1246 115 1276 263
rect 1318 115 1348 263
rect 1522 115 1552 263
rect 1608 115 1638 263
<< pmoshvt >>
rect 80 817 110 1217
rect 166 817 196 1217
rect 356 617 386 1217
rect 428 617 458 1217
rect 548 617 578 1217
rect 620 617 650 1217
rect 706 617 736 1217
rect 778 617 808 1217
rect 898 617 928 1217
rect 970 617 1000 1217
rect 1056 617 1086 1217
rect 1246 817 1276 1217
rect 1332 817 1362 1217
rect 1522 817 1552 1217
rect 1608 817 1638 1217
<< ndiff >>
rect 303 267 356 315
rect 27 199 80 263
rect 27 131 35 199
rect 69 131 80 199
rect 27 115 80 131
rect 110 115 152 263
rect 182 199 235 263
rect 182 131 193 199
rect 227 131 235 199
rect 182 115 235 131
rect 303 131 311 267
rect 345 131 356 267
rect 303 115 356 131
rect 386 115 428 315
rect 458 267 548 315
rect 458 131 469 267
rect 537 131 548 267
rect 458 115 548 131
rect 578 115 620 315
rect 650 199 706 315
rect 650 131 661 199
rect 695 131 706 199
rect 650 115 706 131
rect 736 115 778 315
rect 808 267 898 315
rect 808 131 819 267
rect 887 131 898 267
rect 808 115 898 131
rect 928 115 970 315
rect 1000 267 1056 315
rect 1000 131 1011 267
rect 1045 131 1056 267
rect 1000 115 1056 131
rect 1086 267 1139 315
rect 1086 131 1097 267
rect 1131 131 1139 267
rect 1086 115 1139 131
rect 1193 199 1246 263
rect 1193 131 1201 199
rect 1235 131 1246 199
rect 1193 115 1246 131
rect 1276 115 1318 263
rect 1348 199 1401 263
rect 1348 131 1359 199
rect 1393 131 1401 199
rect 1348 115 1401 131
rect 1469 199 1522 263
rect 1469 131 1477 199
rect 1511 131 1522 199
rect 1469 115 1522 131
rect 1552 199 1608 263
rect 1552 131 1563 199
rect 1597 131 1608 199
rect 1552 115 1608 131
rect 1638 199 1691 263
rect 1638 131 1649 199
rect 1683 131 1691 199
rect 1638 115 1691 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 929 35 1201
rect 69 929 80 1201
rect 27 817 80 929
rect 110 1201 166 1217
rect 110 929 121 1201
rect 155 929 166 1201
rect 110 817 166 929
rect 196 1201 249 1217
rect 196 929 207 1201
rect 241 929 249 1201
rect 196 817 249 929
rect 303 1201 356 1217
rect 303 725 311 1201
rect 345 725 356 1201
rect 303 617 356 725
rect 386 617 428 1217
rect 458 1201 548 1217
rect 458 657 469 1201
rect 537 657 548 1201
rect 458 617 548 657
rect 578 617 620 1217
rect 650 1201 706 1217
rect 650 725 661 1201
rect 695 725 706 1201
rect 650 617 706 725
rect 736 617 778 1217
rect 808 1201 898 1217
rect 808 725 819 1201
rect 887 725 898 1201
rect 808 617 898 725
rect 928 617 970 1217
rect 1000 1201 1056 1217
rect 1000 657 1011 1201
rect 1045 657 1056 1201
rect 1000 617 1056 657
rect 1086 1201 1139 1217
rect 1086 657 1097 1201
rect 1131 657 1139 1201
rect 1193 1201 1246 1217
rect 1193 929 1201 1201
rect 1235 929 1246 1201
rect 1193 817 1246 929
rect 1276 1201 1332 1217
rect 1276 929 1287 1201
rect 1321 929 1332 1201
rect 1276 817 1332 929
rect 1362 1201 1415 1217
rect 1362 929 1373 1201
rect 1407 929 1415 1201
rect 1362 817 1415 929
rect 1469 1201 1522 1217
rect 1469 861 1477 1201
rect 1511 861 1522 1201
rect 1469 817 1522 861
rect 1552 1201 1608 1217
rect 1552 861 1563 1201
rect 1597 861 1608 1201
rect 1552 817 1608 861
rect 1638 1201 1691 1217
rect 1638 861 1649 1201
rect 1683 861 1691 1201
rect 1638 817 1691 861
rect 1086 617 1139 657
<< ndiffc >>
rect 35 131 69 199
rect 193 131 227 199
rect 311 131 345 267
rect 469 131 537 267
rect 661 131 695 199
rect 819 131 887 267
rect 1011 131 1045 267
rect 1097 131 1131 267
rect 1201 131 1235 199
rect 1359 131 1393 199
rect 1477 131 1511 199
rect 1563 131 1597 199
rect 1649 131 1683 199
<< pdiffc >>
rect 35 929 69 1201
rect 121 929 155 1201
rect 207 929 241 1201
rect 311 725 345 1201
rect 469 657 537 1201
rect 661 725 695 1201
rect 819 725 887 1201
rect 1011 657 1045 1201
rect 1097 657 1131 1201
rect 1201 929 1235 1201
rect 1287 929 1321 1201
rect 1373 929 1407 1201
rect 1477 861 1511 1201
rect 1563 861 1597 1201
rect 1649 861 1683 1201
<< psubdiff >>
rect 26 27 50 61
rect 84 27 108 61
rect 162 27 186 61
rect 220 27 244 61
rect 298 27 322 61
rect 356 27 380 61
rect 434 27 458 61
rect 492 27 516 61
rect 570 27 594 61
rect 628 27 652 61
rect 706 27 730 61
rect 764 27 788 61
rect 842 27 866 61
rect 900 27 924 61
rect 978 27 1002 61
rect 1036 27 1060 61
rect 1114 27 1138 61
rect 1172 27 1196 61
rect 1250 27 1274 61
rect 1308 27 1332 61
rect 1386 27 1410 61
rect 1444 27 1468 61
rect 1522 27 1546 61
rect 1580 27 1604 61
<< nsubdiff >>
rect 26 1271 50 1305
rect 84 1271 108 1305
rect 162 1271 186 1305
rect 220 1271 244 1305
rect 298 1271 322 1305
rect 356 1271 380 1305
rect 434 1271 458 1305
rect 492 1271 516 1305
rect 570 1271 594 1305
rect 628 1271 652 1305
rect 706 1271 730 1305
rect 764 1271 788 1305
rect 842 1271 866 1305
rect 900 1271 924 1305
rect 978 1271 1002 1305
rect 1036 1271 1060 1305
rect 1114 1271 1138 1305
rect 1172 1271 1196 1305
rect 1250 1271 1274 1305
rect 1308 1271 1332 1305
rect 1386 1271 1410 1305
rect 1444 1271 1468 1305
rect 1522 1271 1546 1305
rect 1580 1271 1604 1305
<< psubdiffcont >>
rect 50 27 84 61
rect 186 27 220 61
rect 322 27 356 61
rect 458 27 492 61
rect 594 27 628 61
rect 730 27 764 61
rect 866 27 900 61
rect 1002 27 1036 61
rect 1138 27 1172 61
rect 1274 27 1308 61
rect 1410 27 1444 61
rect 1546 27 1580 61
<< nsubdiffcont >>
rect 50 1271 84 1305
rect 186 1271 220 1305
rect 322 1271 356 1305
rect 458 1271 492 1305
rect 594 1271 628 1305
rect 730 1271 764 1305
rect 866 1271 900 1305
rect 1002 1271 1036 1305
rect 1138 1271 1172 1305
rect 1274 1271 1308 1305
rect 1410 1271 1444 1305
rect 1546 1271 1580 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 356 1217 386 1243
rect 428 1217 458 1243
rect 548 1217 578 1243
rect 620 1217 650 1243
rect 706 1217 736 1243
rect 778 1217 808 1243
rect 898 1217 928 1243
rect 970 1217 1000 1243
rect 1056 1217 1086 1243
rect 1246 1217 1276 1243
rect 1332 1217 1362 1243
rect 1522 1217 1552 1243
rect 1608 1217 1638 1243
rect 80 403 110 817
rect 166 494 196 817
rect 37 387 110 403
rect 37 353 47 387
rect 81 353 110 387
rect 37 337 110 353
rect 80 263 110 337
rect 152 478 233 494
rect 152 444 189 478
rect 223 444 233 478
rect 152 428 233 444
rect 356 477 386 617
rect 428 586 458 617
rect 428 570 482 586
rect 428 536 438 570
rect 472 536 482 570
rect 428 520 482 536
rect 356 461 410 477
rect 548 475 578 617
rect 620 580 650 617
rect 706 580 736 617
rect 620 570 736 580
rect 620 536 652 570
rect 686 536 736 570
rect 620 526 736 536
rect 778 475 808 617
rect 898 586 928 617
rect 874 570 928 586
rect 874 536 884 570
rect 918 536 928 570
rect 874 520 928 536
rect 152 263 182 428
rect 356 427 366 461
rect 400 427 410 461
rect 356 411 410 427
rect 452 445 904 475
rect 356 315 386 411
rect 452 367 482 445
rect 874 403 904 445
rect 970 471 1000 617
rect 1056 586 1086 617
rect 1056 570 1127 586
rect 1056 556 1083 570
rect 1067 536 1083 556
rect 1117 536 1127 570
rect 1067 520 1127 536
rect 970 455 1024 471
rect 970 421 980 455
rect 1014 421 1024 455
rect 970 405 1024 421
rect 428 337 482 367
rect 524 387 578 403
rect 524 353 534 387
rect 568 353 578 387
rect 524 337 578 353
rect 428 315 458 337
rect 548 315 578 337
rect 620 387 736 397
rect 620 353 652 387
rect 686 353 736 387
rect 620 343 736 353
rect 620 315 650 343
rect 706 315 736 343
rect 778 387 832 403
rect 778 353 788 387
rect 822 353 832 387
rect 778 337 832 353
rect 874 387 928 403
rect 874 353 884 387
rect 918 353 928 387
rect 874 337 928 353
rect 778 315 808 337
rect 898 315 928 337
rect 970 315 1000 405
rect 1067 367 1097 520
rect 1246 403 1276 817
rect 1056 337 1097 367
rect 1193 387 1276 403
rect 1193 353 1203 387
rect 1237 353 1276 387
rect 1193 337 1276 353
rect 1056 315 1086 337
rect 1246 263 1276 337
rect 1332 351 1362 817
rect 1522 601 1552 817
rect 1512 571 1552 601
rect 1512 471 1542 571
rect 1608 512 1638 817
rect 1487 455 1542 471
rect 1487 421 1497 455
rect 1531 421 1542 455
rect 1584 496 1638 512
rect 1584 462 1594 496
rect 1628 462 1638 496
rect 1584 446 1638 462
rect 1487 405 1542 421
rect 1512 360 1542 405
rect 1332 335 1399 351
rect 1318 301 1355 335
rect 1389 301 1399 335
rect 1512 330 1552 360
rect 1318 285 1399 301
rect 1318 263 1348 285
rect 1522 263 1552 330
rect 1608 263 1638 446
rect 80 89 110 115
rect 152 89 182 115
rect 356 89 386 115
rect 428 89 458 115
rect 548 89 578 115
rect 620 89 650 115
rect 706 89 736 115
rect 778 89 808 115
rect 898 89 928 115
rect 970 89 1000 115
rect 1056 89 1086 115
rect 1246 89 1276 115
rect 1318 89 1348 115
rect 1522 89 1552 115
rect 1608 89 1638 115
<< polycont >>
rect 47 353 81 387
rect 189 444 223 478
rect 438 536 472 570
rect 652 536 686 570
rect 884 536 918 570
rect 366 427 400 461
rect 1083 536 1117 570
rect 980 421 1014 455
rect 534 353 568 387
rect 652 353 686 387
rect 788 353 822 387
rect 884 353 918 387
rect 1203 353 1237 387
rect 1497 421 1531 455
rect 1594 462 1628 496
rect 1355 301 1389 335
<< locali >>
rect 0 1311 1738 1332
rect 0 1271 50 1311
rect 84 1271 186 1311
rect 220 1271 322 1311
rect 356 1271 458 1311
rect 492 1271 594 1311
rect 628 1271 730 1311
rect 764 1271 866 1311
rect 900 1271 1002 1311
rect 1036 1271 1138 1311
rect 1172 1271 1274 1311
rect 1308 1271 1410 1311
rect 1444 1271 1546 1311
rect 1580 1271 1738 1311
rect 35 1201 69 1271
rect 35 913 69 929
rect 121 1201 155 1217
rect 47 387 81 403
rect 47 313 81 353
rect 121 387 155 929
rect 207 1201 241 1271
rect 207 913 241 929
rect 311 1201 345 1271
rect 311 709 345 725
rect 469 1201 537 1217
rect 661 1201 695 1271
rect 661 709 695 725
rect 819 1201 887 1217
rect 469 654 537 657
rect 819 654 887 725
rect 121 233 155 353
rect 189 620 537 654
rect 720 620 887 654
rect 1011 1201 1045 1271
rect 1011 641 1045 657
rect 1097 1201 1131 1217
rect 1201 1201 1235 1271
rect 1201 913 1235 929
rect 1287 1201 1321 1217
rect 1097 654 1131 657
rect 1097 620 1187 654
rect 189 478 223 620
rect 438 570 472 586
rect 438 535 472 536
rect 652 570 686 586
rect 472 501 568 535
rect 189 370 223 444
rect 366 461 400 477
rect 366 411 400 427
rect 534 387 568 501
rect 652 387 686 536
rect 189 336 500 370
rect 534 337 568 353
rect 652 337 686 353
rect 720 387 754 620
rect 884 570 918 586
rect 884 535 918 536
rect 466 283 500 336
rect 720 303 754 353
rect 788 501 884 535
rect 1083 570 1117 586
rect 1083 535 1117 536
rect 788 387 822 501
rect 1151 467 1187 620
rect 964 421 980 455
rect 1014 421 1030 455
rect 1097 433 1187 467
rect 1287 455 1321 929
rect 1373 1201 1407 1271
rect 1373 913 1407 929
rect 1477 1201 1511 1217
rect 1477 609 1511 861
rect 1563 1201 1597 1271
rect 1563 845 1597 861
rect 1649 1201 1683 1217
rect 1649 683 1683 861
rect 1682 666 1683 683
rect 1682 649 1706 666
rect 1649 632 1706 649
rect 1477 570 1511 575
rect 1477 536 1628 570
rect 1594 496 1628 536
rect 1097 387 1131 433
rect 1287 421 1497 455
rect 1531 421 1547 455
rect 868 353 884 387
rect 918 353 1131 387
rect 1187 353 1203 387
rect 1237 353 1253 387
rect 788 337 822 353
rect 35 199 155 233
rect 311 267 345 283
rect 193 199 227 215
rect 35 115 69 131
rect 193 61 227 131
rect 466 267 537 283
rect 720 269 887 303
rect 466 249 469 267
rect 311 61 345 131
rect 819 267 887 269
rect 469 115 537 131
rect 661 199 695 215
rect 661 61 695 131
rect 819 115 887 131
rect 1011 267 1045 283
rect 1011 61 1045 131
rect 1097 267 1131 353
rect 1287 233 1321 421
rect 1594 387 1628 462
rect 1477 353 1628 387
rect 1355 335 1389 351
rect 1097 115 1131 131
rect 1201 199 1321 233
rect 1359 199 1393 215
rect 1201 115 1235 131
rect 1359 61 1393 131
rect 1477 199 1511 353
rect 1672 320 1706 632
rect 1649 286 1706 320
rect 1477 115 1511 131
rect 1563 199 1597 215
rect 1563 61 1597 131
rect 1649 199 1683 286
rect 1649 115 1683 131
rect 0 21 50 61
rect 84 21 186 61
rect 220 21 322 61
rect 356 21 458 61
rect 492 21 594 61
rect 628 21 730 61
rect 764 21 866 61
rect 900 21 1002 61
rect 1036 21 1138 61
rect 1172 21 1274 61
rect 1308 21 1410 61
rect 1444 21 1546 61
rect 1580 21 1738 61
rect 0 0 1738 21
<< viali >>
rect 50 1305 84 1311
rect 50 1277 84 1305
rect 186 1305 220 1311
rect 186 1277 220 1305
rect 322 1305 356 1311
rect 322 1277 356 1305
rect 458 1305 492 1311
rect 458 1277 492 1305
rect 594 1305 628 1311
rect 594 1277 628 1305
rect 730 1305 764 1311
rect 730 1277 764 1305
rect 866 1305 900 1311
rect 866 1277 900 1305
rect 1002 1305 1036 1311
rect 1002 1277 1036 1305
rect 1138 1305 1172 1311
rect 1138 1277 1172 1305
rect 1274 1305 1308 1311
rect 1274 1277 1308 1305
rect 1410 1305 1444 1311
rect 1410 1277 1444 1305
rect 1546 1305 1580 1311
rect 1546 1277 1580 1305
rect 47 279 81 313
rect 121 353 155 387
rect 438 501 472 535
rect 366 427 400 461
rect 634 353 652 387
rect 652 353 668 387
rect 720 353 754 387
rect 884 501 918 535
rect 1083 501 1117 535
rect 980 421 1014 455
rect 1648 649 1682 683
rect 1477 575 1511 609
rect 1497 421 1531 455
rect 1203 353 1237 387
rect 1355 301 1389 313
rect 1355 279 1389 301
rect 50 27 84 55
rect 50 21 84 27
rect 186 27 220 55
rect 186 21 220 27
rect 322 27 356 55
rect 322 21 356 27
rect 458 27 492 55
rect 458 21 492 27
rect 594 27 628 55
rect 594 21 628 27
rect 730 27 764 55
rect 730 21 764 27
rect 866 27 900 55
rect 866 21 900 27
rect 1002 27 1036 55
rect 1002 21 1036 27
rect 1138 27 1172 55
rect 1138 21 1172 27
rect 1274 27 1308 55
rect 1274 21 1308 27
rect 1410 27 1444 55
rect 1410 21 1444 27
rect 1546 27 1580 55
rect 1546 21 1580 27
<< metal1 >>
rect 0 1311 1738 1332
rect 0 1277 50 1311
rect 84 1277 186 1311
rect 220 1277 322 1311
rect 356 1277 458 1311
rect 492 1277 594 1311
rect 628 1277 730 1311
rect 764 1277 866 1311
rect 900 1277 1002 1311
rect 1036 1277 1138 1311
rect 1172 1277 1274 1311
rect 1308 1277 1410 1311
rect 1444 1277 1546 1311
rect 1580 1277 1738 1311
rect 0 1271 1738 1277
rect 1636 683 1694 689
rect 1614 649 1648 683
rect 1682 649 1694 683
rect 1636 643 1694 649
rect 1465 609 1523 615
rect 1442 575 1477 609
rect 1511 575 1523 609
rect 1465 569 1523 575
rect 426 535 484 541
rect 872 535 930 541
rect 1071 535 1129 541
rect 426 501 438 535
rect 472 501 884 535
rect 918 501 1083 535
rect 1117 501 1129 535
rect 426 495 484 501
rect 872 495 930 501
rect 1071 495 1129 501
rect 354 461 412 467
rect 354 427 366 461
rect 400 427 434 461
rect 968 455 1026 461
rect 1485 455 1543 461
rect 354 421 412 427
rect 968 421 980 455
rect 1014 421 1497 455
rect 1531 421 1543 455
rect 968 415 1026 421
rect 1485 415 1543 421
rect 109 387 167 393
rect 622 387 680 393
rect 109 353 121 387
rect 155 353 634 387
rect 668 353 680 387
rect 109 347 167 353
rect 622 347 680 353
rect 708 387 766 393
rect 1191 387 1249 393
rect 708 353 720 387
rect 754 353 1203 387
rect 1237 353 1249 387
rect 708 347 766 353
rect 1191 347 1249 353
rect 35 313 93 319
rect 1343 313 1401 319
rect 35 279 47 313
rect 81 279 1355 313
rect 1389 279 1401 313
rect 35 273 93 279
rect 1343 273 1401 279
rect 0 55 1738 61
rect 0 21 50 55
rect 84 21 186 55
rect 220 21 322 55
rect 356 21 458 55
rect 492 21 594 55
rect 628 21 730 55
rect 764 21 866 55
rect 900 21 1002 55
rect 1036 21 1138 55
rect 1172 21 1274 55
rect 1308 21 1410 55
rect 1444 21 1546 55
rect 1580 21 1738 55
rect 0 0 1738 21
<< labels >>
rlabel viali 383 444 383 444 1 D
port 1 n
rlabel viali 1100 518 1100 518 1 CK
port 2 n
rlabel viali 1665 666 1665 666 1 Q
port 4 n
rlabel viali 1495 592 1495 592 1 QN
port 3 n
rlabel viali 64 296 64 296 1 SN
rlabel viali 67 48 67 48 1 gnd
rlabel viali 67 1284 67 1284 1 vdd
<< end >>
