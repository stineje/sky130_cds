* File: sky130_osu_sc_18T_hs__addh_1.pex.spice
* Created: Fri Nov 12 13:46:12 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%GND 1 2 45 47 55 57 70 86 88
r94 86 88 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r95 72 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r96 68 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r97 68 70 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.825
r98 58 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r99 57 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r100 53 81 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r101 53 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.825
r102 47 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r103 45 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r104 45 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r105 45 72 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r106 45 57 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r107 45 58 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r108 45 47 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r109 2 70 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.825
r110 1 55 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%VDD 1 2 3 37 39 46 50 56 60 68 74 82 86
r57 82 86 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.74 $Y2=6.507
r58 74 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=6.47
+ $X2=3.74 $Y2=6.47
r59 72 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.05 $Y2=6.507
r60 72 74 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.74 $Y2=6.507
r61 68 71 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.05 $Y=3.455
+ $X2=3.05 $Y2=5.835
r62 66 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=6.507
r63 66 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=5.835
r64 63 65 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=6.507
+ $X2=2.38 $Y2=6.507
r65 61 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.61 $Y2=6.507
r66 61 63 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.7 $Y2=6.507
r67 60 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=3.05 $Y2=6.507
r68 60 65 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=2.38 $Y2=6.507
r69 56 59 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.61 $Y=3.795
+ $X2=1.61 $Y2=5.835
r70 54 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=6.507
r71 54 59 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=5.835
r72 51 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=0.75 $Y2=6.507
r73 51 53 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=1.02 $Y2=6.507
r74 50 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.61 $Y2=6.507
r75 50 53 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.02 $Y2=6.507
r76 46 49 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.75 $Y=3.455
+ $X2=0.75 $Y2=5.835
r77 44 77 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=6.507
r78 44 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=5.835
r79 41 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r80 39 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.75 $Y2=6.507
r81 39 41 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.34 $Y2=6.507
r82 37 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r83 37 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r84 37 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r85 37 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r86 37 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r87 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r88 3 71 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=5.835
r89 3 68 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=3.455
r90 2 59 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=5.835
r91 2 56 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=3.795
r92 1 49 150 $w=1.7e-07 $l=2.84825e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.75 $Y2=5.835
r93 1 46 150 $w=1.7e-07 $l=4.59238e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.75 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%CON 1 3 4 15 18 21 22 28 30 31 34 38 40
+ 42 44 48 54 57 58 63 66
c128 66 0 2.7119e-19 $X=3.42 $Y=1.85
c129 58 0 1.57622e-19 $X=0.78 $Y=1.85
c130 42 0 1.92558e-19 $X=3.42 $Y=1.765
r131 58 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.85
+ $X2=0.635 $Y2=1.85
r132 57 63 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=2.62 $Y2=1.85
r133 57 58 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=0.78 $Y2=1.85
r134 56 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.85
+ $X2=3.42 $Y2=1.85
r135 53 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.85
+ $X2=2.62 $Y2=1.85
r136 48 50 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.84 $Y=3.455
+ $X2=3.84 $Y2=5.835
r137 46 48 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.84 $Y=3.035
+ $X2=3.84 $Y2=3.455
r138 42 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.85
r139 42 44 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.165
r140 41 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.95
+ $X2=2.62 $Y2=2.95
r141 40 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=3.84 $Y2=3.035
r142 40 41 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=2.705 $Y2=2.95
r143 39 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.85
+ $X2=2.62 $Y2=1.85
r144 38 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=3.42 $Y2=1.85
r145 38 39 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=2.705 $Y2=1.85
r146 34 36 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.62 $Y=3.455
+ $X2=2.62 $Y2=5.835
r147 32 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=2.95
r148 32 34 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=3.455
r149 31 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.865
+ $X2=2.62 $Y2=2.95
r150 30 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=1.85
r151 30 31 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=2.865
r152 28 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.85
+ $X2=0.635 $Y2=1.85
r153 25 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.35 $Y=1.85
+ $X2=0.635 $Y2=1.85
r154 21 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.85 $X2=0.35 $Y2=1.85
r155 21 23 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=2.015
r156 21 22 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=1.685
r157 18 23 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.015
r158 15 22 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=1.685
r159 4 50 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=5.835
r160 4 48 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=3.455
r161 3 36 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=5.835
r162 3 34 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=3.455
r163 1 44 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=1.165
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%B 3 7 11 15 18 22 25 30 39 42 44
c101 44 0 4.99902e-20 $X=3.21 $Y=2.22
c102 22 0 1.42567e-19 $X=3.205 $Y=2.22
c103 18 0 1.57622e-19 $X=0.905 $Y=2.22
r104 41 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=3.205 $Y=2.22
+ $X2=3.21 $Y2=2.22
r105 41 42 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.205 $Y=2.22
+ $X2=3.06 $Y2=2.22
r106 39 42 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=2.222
+ $X2=3.06 $Y2=2.222
r107 37 39 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=2.22
+ $X2=1.05 $Y2=2.22
r108 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.22
r109 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.22
r110 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=2.22 $X2=3.205 $Y2=2.22
r111 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.385
r112 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=2.22 $X2=0.905 $Y2=2.22
r113 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.385
r114 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.055
r115 15 23 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=3.265 $Y=4.585
+ $X2=3.265 $Y2=2.385
r116 9 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=2.22
r117 9 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=1.075
r118 7 20 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.965 $Y=4.585
+ $X2=0.965 $Y2=2.385
r119 3 19 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.965 $Y=1.075
+ $X2=0.965 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%A 3 7 11 15 18 22 26 31 40 42 43
c87 22 0 1.74252e-19 $X=3.685 $Y=2.59
r88 42 43 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.59
+ $X2=3.54 $Y2=2.59
r89 40 43 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.587
+ $X2=3.54 $Y2=2.587
r90 38 40 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.59
+ $X2=1.53 $Y2=2.59
r91 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.59
r92 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.59
r93 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.59 $X2=3.685 $Y2=2.59
r94 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.755
r95 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.425
r96 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.59 $X2=1.385 $Y2=2.59
r97 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.755
r98 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.425
r99 15 23 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=3.635 $Y=1.075
+ $X2=3.635 $Y2=2.425
r100 11 24 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.625 $Y=4.585
+ $X2=3.625 $Y2=2.755
r101 7 20 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=1.395 $Y=4.585
+ $X2=1.395 $Y2=2.755
r102 3 19 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=1.325 $Y=1.075
+ $X2=1.325 $Y2=2.425
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%A_208_617# 1 3 10 13 15 17 21 23 27 31
+ 33 38 39 42 46 47 50 53 55
c113 31 0 2.52869e-20 $X=2.835 $Y=4.585
c114 23 0 9.69384e-20 $X=2.7 $Y=1.8
r115 55 57 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.955
+ $X2=1.825 $Y2=1.955
r116 54 55 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.955
+ $X2=1.725 $Y2=1.955
r117 52 55 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=1.955
r118 52 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=2.925
r119 48 54 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=1.955
r120 48 50 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=0.825
r121 46 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.725 $Y2=2.925
r122 46 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.265 $Y2=3.01
r123 42 44 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.18 $Y=3.795
+ $X2=1.18 $Y2=5.835
r124 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.265 $Y2=3.01
r125 40 42 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.18 $Y2=3.795
r126 36 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.955 $X2=1.825 $Y2=1.955
r127 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.955
+ $X2=1.825 $Y2=2.12
r128 33 36 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.8
+ $X2=1.825 $Y2=1.955
r129 29 31 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=2.835 $Y=2.745
+ $X2=2.835 $Y2=4.585
r130 25 27 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=1.075
r131 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.8
+ $X2=2.285 $Y2=1.8
r132 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.8
+ $X2=2.775 $Y2=1.725
r133 23 24 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.8 $X2=2.36
+ $Y2=1.8
r134 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=1.8
r135 19 21 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=1.075
r136 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.67
+ $X2=1.885 $Y2=2.67
r137 17 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.67
+ $X2=2.835 $Y2=2.745
r138 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.67 $X2=1.96
+ $Y2=2.67
r139 16 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.8
+ $X2=1.825 $Y2=1.8
r140 15 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=2.285 $Y2=1.8
r141 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=1.96 $Y2=1.8
r142 11 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=2.67
r143 11 13 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=4.585
r144 10 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.67
r145 10 37 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.12
r146 3 44 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=5.835
r147 3 42 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=3.795
r148 1 50 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%S 1 3 10 16 26 29 32
r32 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=3.33
r33 24 26 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=2.385
r34 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=1.475
r35 23 26 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=2.385
r36 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r37 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=3.33
r38 16 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=3.455
r39 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.475
+ $X2=0.26 $Y2=1.475
r40 10 13 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.26 $Y=0.825
+ $X2=0.26 $Y2=1.475
r41 3 21 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r42 3 19 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r43 1 10 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%CO 1 3 11 15 23 26 27 30
c51 26 0 2.52869e-20 $X=2.175 $Y=2.96
r52 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.96
+ $X2=2.175 $Y2=2.96
r53 26 28 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=3.045
r54 26 27 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=2.875
r55 21 23 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.472
+ $X2=2.175 $Y2=1.472
r56 19 23 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=1.472
r57 19 27 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=2.875
r58 15 17 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.1 $Y=3.455
+ $X2=2.1 $Y2=5.835
r59 15 28 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.1 $Y=3.455 $X2=2.1
+ $Y2=3.045
r60 9 21 0.89264 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.07 $Y=1.385 $X2=2.07
+ $Y2=1.472
r61 9 11 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.07 $Y=1.385
+ $X2=2.07 $Y2=0.825
r62 3 17 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.96
+ $Y=3.085 $X2=2.1 $Y2=5.835
r63 3 15 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.96
+ $Y=3.085 $X2=2.1 $Y2=3.455
r64 1 11 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__ADDH_1%A_570_115# 1 2 11 13 14
r11 15 17 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.85 $Y=0.72
+ $X2=3.85 $Y2=0.825
r12 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.85 $Y2=0.72
r13 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.075 $Y2=0.635
r14 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.72
+ $X2=3.075 $Y2=0.635
r15 9 11 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.72
+ $X2=2.99 $Y2=0.825
r16 2 17 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.825
r17 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.825
.ends

