* File: sky130_osu_sc_12T_ms__inv_8.pex.spice
* Created: Fri Nov 12 15:24:47 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__INV_8%GND 1 2 3 4 5 51 55 57 64 66 73 75 82 84
+ 92 104 106
r120 104 106 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.06 $Y2=0.152
r121 90 92 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.755
r122 85 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r123 84 90 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=3.615 $Y=0.152
+ $X2=3.7 $Y2=0.305
r124 80 100 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r125 80 82 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.755
r126 76 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r127 75 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r128 71 99 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r129 71 73 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r130 67 98 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r131 66 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r132 62 98 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r133 62 64 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r134 57 98 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r135 53 55 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r136 51 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=0.19
+ $X2=3.06 $Y2=0.19
r137 51 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r138 51 53 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r139 51 58 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r140 51 84 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r141 51 85 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r142 51 75 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r143 51 76 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r144 51 66 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r145 51 67 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r146 51 57 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r147 51 58 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r148 5 92 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.755
r149 4 82 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.7 $Y=0.575
+ $X2=2.84 $Y2=0.755
r150 3 73 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.755
r151 2 64 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.755
r152 1 55 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__INV_8%VDD 1 2 3 4 5 41 45 47 53 57 63 67 73 77
+ 84 95 99
r77 95 99 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=3.06 $Y2=4.287
r78 89 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r79 84 87 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=2.955 $X2=3.7
+ $Y2=3.635
r80 82 87 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.7 $Y=4.135 $X2=3.7
+ $Y2=3.635
r81 80 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=4.25
+ $X2=3.06 $Y2=4.25
r82 78 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=4.287
+ $X2=2.84 $Y2=4.287
r83 78 80 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=4.287
+ $X2=3.06 $Y2=4.287
r84 77 82 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=3.615 $Y=4.287
+ $X2=3.7 $Y2=4.135
r85 77 80 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=4.287
+ $X2=3.06 $Y2=4.287
r86 73 76 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=2.955
+ $X2=2.84 $Y2=3.635
r87 71 93 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=4.135
+ $X2=2.84 $Y2=4.287
r88 71 76 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.84 $Y=4.135 $X2=2.84
+ $Y2=3.635
r89 68 92 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=1.98 $Y2=4.287
r90 68 70 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=2.38 $Y2=4.287
r91 67 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.84 $Y2=4.287
r92 67 70 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.38 $Y2=4.287
r93 63 66 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r94 61 92 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=4.287
r95 61 66 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135 $X2=1.98
+ $Y2=3.635
r96 58 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r97 58 60 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r98 57 92 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.287
r99 57 60 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r100 53 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r101 51 91 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r102 51 56 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.635
r103 48 89 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r104 48 50 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r105 47 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r106 47 50 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r107 43 89 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r108 43 45 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r109 41 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r110 41 70 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r111 41 60 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r112 41 50 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r113 41 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r114 5 87 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=3.635
r115 5 84 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=2.955
r116 4 76 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=3.635
r117 4 73 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=2.955
r118 3 66 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r119 3 63 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r120 2 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r121 2 53 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r122 1 45 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__INV_8%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 45 47 49 50 52 53 55 57 59 60 62 63 65 67 69
+ 70 72 73 75 77 79 80 82 83 85 86 88 89 90 91 92 93 94 95 96 97 98 99 100 103
+ 105 107 110
c234 70 0 1.33323e-19 $X=3.055 $Y=2.48
c235 67 0 1.33323e-19 $X=3.055 $Y=1.22
c236 60 0 1.33323e-19 $X=2.625 $Y=2.48
c237 57 0 1.33323e-19 $X=2.625 $Y=1.22
c238 50 0 1.33323e-19 $X=2.195 $Y=2.48
c239 45 0 1.33323e-19 $X=2.195 $Y=1.22
c240 38 0 1.33323e-19 $X=1.765 $Y=2.48
c241 35 0 1.33323e-19 $X=1.765 $Y=1.22
c242 28 0 1.33323e-19 $X=1.335 $Y=2.48
c243 25 0 1.33323e-19 $X=1.335 $Y=1.22
c244 18 0 1.33323e-19 $X=0.905 $Y=2.48
c245 15 0 1.33323e-19 $X=0.905 $Y=1.22
r246 110 113 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=2.845
+ $X2=0.405 $Y2=2.85
r247 105 107 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=1.825
+ $X2=0.535 $Y2=1.825
r248 103 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r249 101 105 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.405 $Y2=1.825
r250 101 103 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.32 $Y2=2.85
r251 85 107 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.825 $X2=0.535 $Y2=1.825
r252 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.99
r253 85 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.66
r254 80 82 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.485 $Y=2.48
+ $X2=3.485 $Y2=3.235
r255 77 79 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.485 $Y=1.22
+ $X2=3.485 $Y2=0.835
r256 76 100 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.405
+ $X2=3.055 $Y2=2.405
r257 75 80 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=2.405
+ $X2=3.485 $Y2=2.48
r258 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.405
+ $X2=3.13 $Y2=2.405
r259 74 99 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.295
+ $X2=3.055 $Y2=1.295
r260 73 77 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.485 $Y2=1.22
r261 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.13 $Y2=1.295
r262 70 100 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.48
+ $X2=3.055 $Y2=2.405
r263 70 72 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.055 $Y=2.48
+ $X2=3.055 $Y2=3.235
r264 67 99 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.22
+ $X2=3.055 $Y2=1.295
r265 67 69 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.055 $Y=1.22
+ $X2=3.055 $Y2=0.835
r266 66 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.405
+ $X2=2.625 $Y2=2.405
r267 65 100 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.405
+ $X2=3.055 $Y2=2.405
r268 65 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.405
+ $X2=2.7 $Y2=2.405
r269 64 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.295
+ $X2=2.625 $Y2=1.295
r270 63 99 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.295
+ $X2=3.055 $Y2=1.295
r271 63 64 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.295
+ $X2=2.7 $Y2=1.295
r272 60 98 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=2.405
r273 60 62 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=3.235
r274 57 97 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.22
+ $X2=2.625 $Y2=1.295
r275 57 59 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.625 $Y=1.22
+ $X2=2.625 $Y2=0.835
r276 56 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.405
+ $X2=2.195 $Y2=2.405
r277 55 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.625 $Y2=2.405
r278 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.27 $Y2=2.405
r279 54 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.295
+ $X2=2.195 $Y2=1.295
r280 53 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.295
+ $X2=2.625 $Y2=1.295
r281 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.295
+ $X2=2.27 $Y2=1.295
r282 50 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=2.405
r283 50 52 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=3.235
r284 49 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.33
+ $X2=2.195 $Y2=2.405
r285 48 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.37
+ $X2=2.195 $Y2=1.295
r286 48 49 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.37
+ $X2=2.195 $Y2=2.33
r287 45 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.22
+ $X2=2.195 $Y2=1.295
r288 45 47 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.195 $Y=1.22
+ $X2=2.195 $Y2=0.835
r289 44 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.405
+ $X2=1.765 $Y2=2.405
r290 43 96 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=2.195 $Y2=2.405
r291 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=1.84 $Y2=2.405
r292 42 93 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.295
+ $X2=1.765 $Y2=1.295
r293 41 95 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.295
+ $X2=2.195 $Y2=1.295
r294 41 42 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.295
+ $X2=1.84 $Y2=1.295
r295 38 94 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=2.405
r296 38 40 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r297 35 93 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.22
+ $X2=1.765 $Y2=1.295
r298 35 37 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.765 $Y=1.22
+ $X2=1.765 $Y2=0.835
r299 34 92 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.405
+ $X2=1.335 $Y2=2.405
r300 33 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.405
r301 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.41 $Y2=2.405
r302 32 91 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.335 $Y2=1.295
r303 31 93 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.295
+ $X2=1.765 $Y2=1.295
r304 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.295
+ $X2=1.41 $Y2=1.295
r305 28 92 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=2.405
r306 28 30 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r307 25 91 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=1.295
r308 25 27 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=0.835
r309 24 90 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.405
+ $X2=0.905 $Y2=2.405
r310 23 92 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=1.335 $Y2=2.405
r311 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=0.98 $Y2=2.405
r312 22 89 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.295
+ $X2=0.905 $Y2=1.295
r313 21 91 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=1.335 $Y2=1.295
r314 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=0.98 $Y2=1.295
r315 18 90 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=2.405
r316 18 20 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=3.235
r317 15 89 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=1.295
r318 15 17 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=0.835
r319 14 88 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.405
+ $X2=0.475 $Y2=2.405
r320 13 90 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.905 $Y2=2.405
r321 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.55 $Y2=2.405
r322 12 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.475 $Y2=1.295
r323 11 89 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.905 $Y2=1.295
r324 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.55 $Y2=1.295
r325 8 88 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=2.405
r326 8 10 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=3.235
r327 7 88 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=2.405
r328 7 87 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=1.99
r329 4 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.295
r330 4 86 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.66
r331 1 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=1.295
r332 1 3 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__INV_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68 76
+ 82 89 90 92 94 96 99 100 101 102 103 105 106 107 108 109 110 111
c181 111 0 1.33323e-19 $X=3.27 $Y=2.365
c182 110 0 1.33323e-19 $X=3.27 $Y=1.115
c183 109 0 2.66647e-19 $X=2.555 $Y=2.48
c184 107 0 2.66647e-19 $X=2.555 $Y=1
c185 103 0 2.66647e-19 $X=1.695 $Y=2.48
c186 101 0 2.66647e-19 $X=1.695 $Y=1
c187 90 0 1.33323e-19 $X=0.69 $Y=2.365
c188 89 0 1.33323e-19 $X=0.69 $Y=1.115
r189 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.365
+ $X2=3.27 $Y2=2.48
r190 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.115
+ $X2=3.27 $Y2=1
r191 110 111 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.27 $Y=1.115
+ $X2=3.27 $Y2=2.365
r192 109 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.48
+ $X2=2.41 $Y2=2.48
r193 108 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.48
+ $X2=3.27 $Y2=2.48
r194 108 109 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.48
+ $X2=2.555 $Y2=2.48
r195 107 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1
+ $X2=2.41 $Y2=1
r196 106 125 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1
+ $X2=3.27 $Y2=1
r197 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1
+ $X2=2.555 $Y2=1
r198 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.365
+ $X2=2.41 $Y2=2.48
r199 104 121 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=1
r200 104 105 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=2.365
r201 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.48
+ $X2=1.55 $Y2=2.48
r202 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.48
+ $X2=2.41 $Y2=2.48
r203 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.48
+ $X2=1.695 $Y2=2.48
r204 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1
+ $X2=1.55 $Y2=1
r205 100 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=2.41 $Y2=1
r206 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=1.695 $Y2=1
r207 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.48
r208 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r209 98 99 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=2.365
r210 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.48
+ $X2=0.69 $Y2=2.48
r211 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=1.55 $Y2=2.48
r212 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=0.835 $Y2=2.48
r213 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1
+ $X2=0.69 $Y2=1
r214 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=1.55 $Y2=1
r215 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=0.835 $Y2=1
r216 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.48
r217 90 92 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=1.72
r218 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1
r219 89 92 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1.72
r220 85 87 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=2.955
+ $X2=3.27 $Y2=3.635
r221 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.48
+ $X2=3.27 $Y2=2.48
r222 82 85 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.27 $Y=2.48
+ $X2=3.27 $Y2=2.955
r223 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1 $X2=3.27
+ $Y2=1
r224 76 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.27 $Y=0.755
+ $X2=3.27 $Y2=1
r225 71 73 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=2.955
+ $X2=2.41 $Y2=3.635
r226 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.48
+ $X2=2.41 $Y2=2.48
r227 68 71 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.41 $Y=2.48
+ $X2=2.41 $Y2=2.955
r228 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1 $X2=2.41
+ $Y2=1
r229 62 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.41 $Y=0.755
+ $X2=2.41 $Y2=1
r230 57 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r231 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.48
r232 54 57 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.955
r233 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r234 48 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r235 43 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r236 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r237 40 43 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.955
r238 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1 $X2=0.69
+ $Y2=1
r239 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0.755
+ $X2=0.69 $Y2=1
r240 12 87 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=3.635
r241 12 85 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=2.955
r242 11 73 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=3.635
r243 11 71 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=2.955
r244 10 59 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r245 10 57 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r246 9 45 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r247 9 43 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r248 4 76 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.755
r249 3 62 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.755
r250 2 48 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
r251 1 34 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

