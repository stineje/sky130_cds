* File: sky130_osu_sc_15T_ls__addh_l.pex.spice
* Created: Fri Nov 12 14:53:15 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%GND 1 2 45 47 55 57 70 86 88
r96 86 88 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r97 72 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r98 68 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r99 68 70 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.74
r100 58 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r101 57 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r102 53 81 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r103 53 55 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.74
r104 47 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r105 45 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r106 45 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r107 45 72 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r108 45 57 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r109 45 58 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r110 45 47 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r111 2 70 91 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.74
r112 1 55 91 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%VDD 1 2 3 37 39 46 50 56 60 68 74 82 86
r57 82 86 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=3.74 $Y2=5.397
r58 74 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=5.36
+ $X2=3.74 $Y2=5.36
r59 72 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=5.397
+ $X2=3.05 $Y2=5.397
r60 72 74 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=5.397
+ $X2=3.74 $Y2=5.397
r61 68 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.05 $Y=3.215
+ $X2=3.05 $Y2=4.575
r62 66 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=5.245
+ $X2=3.05 $Y2=5.397
r63 66 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=5.245
+ $X2=3.05 $Y2=4.575
r64 63 65 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=5.397
+ $X2=2.38 $Y2=5.397
r65 61 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=5.397
+ $X2=1.61 $Y2=5.397
r66 61 63 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=5.397
+ $X2=1.7 $Y2=5.397
r67 60 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=5.397
+ $X2=3.05 $Y2=5.397
r68 60 65 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=5.397
+ $X2=2.38 $Y2=5.397
r69 56 59 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.61 $Y=3.555
+ $X2=1.61 $Y2=4.575
r70 54 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=5.245
+ $X2=1.61 $Y2=5.397
r71 54 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.61 $Y=5.245
+ $X2=1.61 $Y2=4.575
r72 51 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=5.397
+ $X2=0.75 $Y2=5.397
r73 51 53 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=5.397
+ $X2=1.02 $Y2=5.397
r74 50 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=5.397
+ $X2=1.61 $Y2=5.397
r75 50 53 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=5.397
+ $X2=1.02 $Y2=5.397
r76 46 49 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.75 $Y=3.215
+ $X2=0.75 $Y2=4.575
r77 44 77 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=5.245
+ $X2=0.75 $Y2=5.397
r78 44 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.75 $Y=5.245
+ $X2=0.75 $Y2=4.575
r79 41 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r80 39 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=5.397
+ $X2=0.75 $Y2=5.397
r81 39 41 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=5.397
+ $X2=0.34 $Y2=5.397
r82 37 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r83 37 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r84 37 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r85 37 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r86 37 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r87 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r88 3 59 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.825 $X2=1.61 $Y2=4.575
r89 3 56 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.825 $X2=1.61 $Y2=3.555
r90 2 49 240 $w=1.7e-07 $l=1.10549e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.565 $X2=0.75 $Y2=4.575
r91 2 46 240 $w=1.7e-07 $l=4.38748e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.565 $X2=0.75 $Y2=3.215
r92 1 71 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=2.825 $X2=3.05 $Y2=4.575
r93 1 68 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=2.825 $X2=3.05 $Y2=3.215
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%CON 1 3 4 15 19 22 29 31 32 35 39 41 43
+ 45 49 55 58 59 64 67
c128 67 0 2.7119e-19 $X=3.42 $Y=1.59
c129 59 0 1.57622e-19 $X=0.78 $Y=1.59
c130 43 0 1.92558e-19 $X=3.42 $Y=1.505
r131 59 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.59
+ $X2=0.635 $Y2=1.59
r132 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.59
+ $X2=2.62 $Y2=1.59
r133 58 59 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.59
+ $X2=0.78 $Y2=1.59
r134 57 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.59
+ $X2=3.42 $Y2=1.59
r135 54 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.59
+ $X2=2.62 $Y2=1.59
r136 49 51 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.84 $Y=3.215
+ $X2=3.84 $Y2=4.575
r137 47 49 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.84 $Y=2.775
+ $X2=3.84 $Y2=3.215
r138 43 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.505
+ $X2=3.42 $Y2=1.59
r139 43 45 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.42 $Y=1.505
+ $X2=3.42 $Y2=1.065
r140 42 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.69
+ $X2=2.62 $Y2=2.69
r141 41 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.69
+ $X2=3.84 $Y2=2.775
r142 41 42 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.69
+ $X2=2.705 $Y2=2.69
r143 40 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.59
+ $X2=2.62 $Y2=1.59
r144 39 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.59
+ $X2=3.42 $Y2=1.59
r145 39 40 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.59
+ $X2=2.705 $Y2=1.59
r146 35 37 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.62 $Y=3.215
+ $X2=2.62 $Y2=4.575
r147 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.775
+ $X2=2.62 $Y2=2.69
r148 33 35 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.62 $Y=2.775
+ $X2=2.62 $Y2=3.215
r149 32 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.605
+ $X2=2.62 $Y2=2.69
r150 31 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.675
+ $X2=2.62 $Y2=1.59
r151 31 32 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.675
+ $X2=2.62 $Y2=2.605
r152 29 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.59
+ $X2=0.635 $Y2=1.59
r153 26 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.35 $Y=1.59
+ $X2=0.635 $Y2=1.59
r154 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.59 $X2=0.35 $Y2=1.59
r155 22 24 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.59
+ $X2=0.382 $Y2=1.755
r156 22 23 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.59
+ $X2=0.382 $Y2=1.425
r157 19 24 1251.15 $w=1.5e-07 $l=2.44e-06 $layer=POLY_cond $X=0.475 $Y=4.195
+ $X2=0.475 $Y2=1.755
r158 15 23 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.425
r159 4 51 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=2.825 $X2=3.84 $Y2=4.575
r160 4 49 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=2.825 $X2=3.84 $Y2=3.215
r161 3 37 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=2.825 $X2=2.62 $Y2=4.575
r162 3 35 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=2.825 $X2=2.62 $Y2=3.215
r163 1 45 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=1.065
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%B 3 7 11 15 18 22 25 30 39 42 44
c102 44 0 4.99902e-20 $X=3.21 $Y=1.96
c103 22 0 1.42567e-19 $X=3.205 $Y=1.96
c104 18 0 1.57622e-19 $X=0.905 $Y=1.96
c105 7 0 4.43035e-20 $X=0.965 $Y=3.825
r106 41 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=3.205 $Y=1.96
+ $X2=3.21 $Y2=1.96
r107 41 42 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.205 $Y=1.96
+ $X2=3.06 $Y2=1.96
r108 39 42 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=1.962
+ $X2=3.06 $Y2=1.962
r109 37 39 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=1.96
+ $X2=1.05 $Y2=1.96
r110 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=1.96
+ $X2=3.205 $Y2=1.96
r111 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=1.96
r112 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.96 $X2=3.205 $Y2=1.96
r113 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.96
+ $X2=3.205 $Y2=2.125
r114 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.96 $X2=0.905 $Y2=1.96
r115 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=2.125
r116 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=1.795
r117 15 23 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=3.265 $Y=3.825
+ $X2=3.265 $Y2=2.125
r118 9 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.795
+ $X2=3.205 $Y2=1.96
r119 9 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.205 $Y=1.795
+ $X2=3.205 $Y2=0.945
r120 7 20 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=0.965 $Y=3.825
+ $X2=0.965 $Y2=2.125
r121 3 19 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.965 $Y=0.945
+ $X2=0.965 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%A 3 7 11 15 18 22 26 31 40 42 43
c87 22 0 1.74252e-19 $X=3.685 $Y=2.33
r88 42 43 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.33
+ $X2=3.54 $Y2=2.33
r89 40 43 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.327
+ $X2=3.54 $Y2=2.327
r90 38 40 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.33
+ $X2=1.53 $Y2=2.33
r91 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.33
+ $X2=3.685 $Y2=2.33
r92 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.33
+ $X2=1.385 $Y2=2.33
r93 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.33 $X2=3.685 $Y2=2.33
r94 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.33
+ $X2=3.685 $Y2=2.495
r95 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.33
+ $X2=3.685 $Y2=2.165
r96 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.33 $X2=1.385 $Y2=2.33
r97 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.33
+ $X2=1.385 $Y2=2.495
r98 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.33
+ $X2=1.385 $Y2=2.165
r99 15 23 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=3.635 $Y=0.945
+ $X2=3.635 $Y2=2.165
r100 11 24 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.625 $Y=3.825
+ $X2=3.625 $Y2=2.495
r101 7 20 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.395 $Y=3.825
+ $X2=1.395 $Y2=2.495
r102 3 19 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.325 $Y=0.945
+ $X2=1.325 $Y2=2.165
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%A_208_565# 1 3 10 13 15 17 21 23 27 31
+ 33 38 39 42 46 47 50 53 55
c113 31 0 2.52869e-20 $X=2.835 $Y=3.825
c114 23 0 9.69384e-20 $X=2.7 $Y=1.54
r115 55 57 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.695
+ $X2=1.825 $Y2=1.695
r116 54 55 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.695
+ $X2=1.725 $Y2=1.695
r117 52 55 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.86
+ $X2=1.725 $Y2=1.695
r118 52 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=1.86
+ $X2=1.725 $Y2=2.665
r119 48 54 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.53
+ $X2=1.54 $Y2=1.695
r120 48 50 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.54 $Y=1.53
+ $X2=1.54 $Y2=0.74
r121 46 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=2.75
+ $X2=1.725 $Y2=2.665
r122 46 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=2.75
+ $X2=1.265 $Y2=2.75
r123 42 44 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.18 $Y=3.555
+ $X2=1.18 $Y2=4.575
r124 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=2.835
+ $X2=1.265 $Y2=2.75
r125 40 42 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.18 $Y=2.835
+ $X2=1.18 $Y2=3.555
r126 36 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.695 $X2=1.825 $Y2=1.695
r127 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.695
+ $X2=1.825 $Y2=1.86
r128 33 36 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.54
+ $X2=1.825 $Y2=1.695
r129 29 31 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=2.835 $Y=2.485
+ $X2=2.835 $Y2=3.825
r130 25 27 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.775 $Y=1.465
+ $X2=2.775 $Y2=0.945
r131 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.54
+ $X2=2.285 $Y2=1.54
r132 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.54
+ $X2=2.775 $Y2=1.465
r133 23 24 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.54 $X2=2.36
+ $Y2=1.54
r134 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.465
+ $X2=2.285 $Y2=1.54
r135 19 21 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=2.285 $Y=1.465
+ $X2=2.285 $Y2=0.88
r136 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.41
+ $X2=1.885 $Y2=2.41
r137 17 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.41
+ $X2=2.835 $Y2=2.485
r138 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.41 $X2=1.96
+ $Y2=2.41
r139 16 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.54
+ $X2=1.825 $Y2=1.54
r140 15 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.54
+ $X2=2.285 $Y2=1.54
r141 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.54
+ $X2=1.96 $Y2=1.54
r142 11 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.485
+ $X2=1.885 $Y2=2.41
r143 11 13 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=1.885 $Y=2.485
+ $X2=1.885 $Y2=4.195
r144 10 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.335
+ $X2=1.885 $Y2=2.41
r145 10 37 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.335
+ $X2=1.885 $Y2=1.86
r146 3 44 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.825 $X2=1.18 $Y2=4.575
r147 3 42 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.825 $X2=1.18 $Y2=3.555
r148 1 50 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%S 1 3 10 16 26 29 32
c31 32 0 4.43035e-20 $X=0.26 $Y=3.07
r32 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.07
r33 24 26 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=2.125
r34 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.33
+ $X2=0.26 $Y2=1.215
r35 23 26 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.33
+ $X2=0.26 $Y2=2.125
r36 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.895
+ $X2=0.26 $Y2=4.575
r37 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.07
+ $X2=0.26 $Y2=3.07
r38 16 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.26 $Y=3.07
+ $X2=0.26 $Y2=3.895
r39 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.215
+ $X2=0.26 $Y2=1.215
r40 10 13 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.26 $Y=0.825
+ $X2=0.26 $Y2=1.215
r41 3 21 400 $w=1.7e-07 $l=1.07068e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.575
r42 3 19 400 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=3.895
r43 1 10 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%CO 1 3 11 15 23 26 27 30
c53 26 0 2.52869e-20 $X=2.175 $Y=2.7
r54 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.7
+ $X2=2.175 $Y2=2.7
r55 26 28 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.7
+ $X2=2.137 $Y2=2.785
r56 26 27 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.7
+ $X2=2.137 $Y2=2.615
r57 21 23 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.215
+ $X2=2.175 $Y2=1.215
r58 19 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=1.3
+ $X2=2.175 $Y2=1.215
r59 19 27 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.3
+ $X2=2.175 $Y2=2.615
r60 15 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.1 $Y=3.895 $X2=2.1
+ $Y2=4.575
r61 15 28 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.1 $Y=3.895
+ $X2=2.1 $Y2=2.785
r62 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.13 $X2=2.07
+ $Y2=1.215
r63 9 11 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.07 $Y=1.13
+ $X2=2.07 $Y2=0.825
r64 3 17 400 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=3.565 $X2=2.1 $Y2=4.575
r65 3 15 400 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=3.565 $X2=2.1 $Y2=3.895
r66 1 11 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ADDH_L%A_570_115# 1 2 11 13 14
r11 15 17 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.85 $Y=0.645
+ $X2=3.85 $Y2=0.74
r12 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.56
+ $X2=3.85 $Y2=0.645
r13 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.56
+ $X2=3.075 $Y2=0.56
r14 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.645
+ $X2=3.075 $Y2=0.56
r15 9 11 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.99 $Y=0.645
+ $X2=2.99 $Y2=0.74
r16 2 17 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.74
r17 1 11 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.74
.ends

