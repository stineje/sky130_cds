* File: sky130_osu_sc_12T_hs__oai22_l.pxi.spice
* Created: Fri Nov 12 15:12:26 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%GND N_GND_M1003_d N_GND_M1003_b N_GND_c_3_p
+ N_GND_c_4_p GND N_GND_c_5_p PM_SKY130_OSU_SC_12T_HS__OAI22_L%GND
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%VDD N_VDD_M1000_s N_VDD_M1004_d N_VDD_M1000_b
+ N_VDD_c_47_p N_VDD_c_48_p N_VDD_c_61_p VDD N_VDD_c_49_p
+ PM_SKY130_OSU_SC_12T_HS__OAI22_L%VDD
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%A0 N_A0_c_67_n N_A0_c_68_n N_A0_M1003_g
+ N_A0_c_72_n N_A0_M1000_g N_A0_c_73_n N_A0_c_80_n A0
+ PM_SKY130_OSU_SC_12T_HS__OAI22_L%A0
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%A1 N_A1_M1006_g N_A1_M1001_g N_A1_c_99_n
+ N_A1_c_100_n A1 PM_SKY130_OSU_SC_12T_HS__OAI22_L%A1
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%B0 N_B0_M1002_g N_B0_M1005_g N_B0_c_141_n
+ N_B0_c_142_n N_B0_c_143_n B0 PM_SKY130_OSU_SC_12T_HS__OAI22_L%B0
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%B1 N_B1_c_193_n N_B1_M1004_g N_B1_M1007_g
+ N_B1_c_196_n B1 PM_SKY130_OSU_SC_12T_HS__OAI22_L%B1
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%Y N_Y_M1002_d N_Y_M1006_d N_Y_c_220_n
+ N_Y_c_228_n N_Y_c_224_n N_Y_c_217_n N_Y_c_218_n Y
+ PM_SKY130_OSU_SC_12T_HS__OAI22_L%Y
x_PM_SKY130_OSU_SC_12T_HS__OAI22_L%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1001_d N_A_27_115#_M1007_d N_A_27_115#_c_259_n
+ N_A_27_115#_c_262_n N_A_27_115#_c_265_n N_A_27_115#_c_266_n
+ N_A_27_115#_c_268_n N_A_27_115#_c_271_n
+ PM_SKY130_OSU_SC_12T_HS__OAI22_L%A_27_115#
cc_1 N_GND_M1003_b N_A0_c_67_n 0.0582151f $X=-0.045 $Y=0 $X2=0.345 $Y2=2.085
cc_2 N_GND_M1003_b N_A0_c_68_n 0.0204667f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.23
cc_3 N_GND_c_3_p N_A0_c_68_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.23
cc_4 N_GND_c_4_p N_A0_c_68_n 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=1.23
cc_5 N_GND_c_5_p N_A0_c_68_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=1.23
cc_6 N_GND_M1003_b N_A0_c_72_n 0.0357139f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.445
cc_7 N_GND_M1003_b N_A0_c_73_n 0.0236679f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.307
cc_8 N_GND_M1003_b A0 0.0213621f $X=-0.045 $Y=0 $X2=0.345 $Y2=2.11
cc_9 N_GND_M1003_b N_A1_M1006_g 0.0298922f $X=-0.045 $Y=0 $X2=0.835 $Y2=3.235
cc_10 N_GND_M1003_b N_A1_M1001_g 0.0422444f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.85
cc_11 N_GND_c_4_p N_A1_M1001_g 0.00263049f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.85
cc_12 N_GND_c_5_p N_A1_M1001_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.905 $Y2=0.85
cc_13 N_GND_M1003_b N_A1_c_99_n 0.0311068f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.74
cc_14 N_GND_M1003_b N_A1_c_100_n 0.00291407f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.74
cc_15 N_GND_M1003_b A1 0.00481617f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.74
cc_16 N_GND_M1003_b N_B0_M1002_g 0.0440457f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.85
cc_17 N_GND_c_5_p N_B0_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335 $Y2=0.85
cc_18 N_GND_M1003_b N_B0_M1005_g 0.0202068f $X=-0.045 $Y=0 $X2=1.335 $Y2=3.235
cc_19 N_GND_M1003_b N_B0_c_141_n 0.0276507f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.85
cc_20 N_GND_M1003_b N_B0_c_142_n 0.00340289f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.48
cc_21 N_GND_M1003_b N_B0_c_143_n 0.00354178f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.85
cc_22 N_GND_M1003_b B0 0.00578565f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.48
cc_23 N_GND_M1003_b N_B1_c_193_n 0.0700015f $X=-0.045 $Y=0 $X2=1.695 $Y2=2.52
cc_24 N_GND_M1003_b N_B1_M1007_g 0.0802435f $X=-0.045 $Y=0 $X2=1.765 $Y2=0.85
cc_25 N_GND_c_5_p N_B1_M1007_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765 $Y2=0.85
cc_26 N_GND_M1003_b N_B1_c_196_n 0.0125315f $X=-0.045 $Y=0 $X2=2.005 $Y2=2.115
cc_27 N_GND_M1003_b B1 0.00895888f $X=-0.045 $Y=0 $X2=2.005 $Y2=2.115
cc_28 N_GND_M1003_b N_Y_c_217_n 0.00215516f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.235
cc_29 N_GND_M1003_b N_Y_c_218_n 0.00880857f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.74
cc_30 N_GND_M1003_b Y 0.00647907f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.74
cc_31 N_GND_M1003_b N_A_27_115#_c_259_n 0.0015601f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_32 N_GND_c_3_p N_A_27_115#_c_259_n 0.00735421f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_33 N_GND_c_5_p N_A_27_115#_c_259_n 0.00476028f $X=1.7 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_34 N_GND_M1003_d N_A_27_115#_c_262_n 0.00176461f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.16
cc_35 N_GND_M1003_b N_A_27_115#_c_262_n 0.0100074f $X=-0.045 $Y=0 $X2=1.035
+ $Y2=1.16
cc_36 N_GND_c_4_p N_A_27_115#_c_262_n 0.0135055f $X=0.69 $Y=0.74 $X2=1.035
+ $Y2=1.16
cc_37 N_GND_M1003_b N_A_27_115#_c_265_n 0.00830224f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.16
cc_38 N_GND_M1003_b N_A_27_115#_c_266_n 0.034563f $X=-0.045 $Y=0 $X2=1.895
+ $Y2=0.63
cc_39 N_GND_c_5_p N_A_27_115#_c_266_n 0.0189415f $X=1.7 $Y=0.19 $X2=1.895
+ $Y2=0.63
cc_40 N_GND_M1003_b N_A_27_115#_c_268_n 0.0104598f $X=-0.045 $Y=0 $X2=1.205
+ $Y2=0.63
cc_41 N_GND_c_4_p N_A_27_115#_c_268_n 0.00181622f $X=0.69 $Y=0.74 $X2=1.205
+ $Y2=0.63
cc_42 N_GND_c_5_p N_A_27_115#_c_268_n 0.00490588f $X=1.7 $Y=0.19 $X2=1.205
+ $Y2=0.63
cc_43 N_GND_M1003_b N_A_27_115#_c_271_n 0.0109759f $X=-0.045 $Y=0 $X2=1.98
+ $Y2=0.63
cc_44 N_GND_c_5_p N_A_27_115#_c_271_n 0.00475375f $X=1.7 $Y=0.19 $X2=1.98
+ $Y2=0.63
cc_45 N_VDD_M1000_b N_A0_c_72_n 0.00966186f $X=-0.045 $Y=2.415 $X2=0.475
+ $Y2=2.445
cc_46 N_VDD_M1000_b N_A0_M1000_g 0.0234447f $X=-0.045 $Y=2.415 $X2=0.475
+ $Y2=3.235
cc_47 N_VDD_c_47_p N_A0_M1000_g 0.00502587f $X=0.26 $Y=3.35 $X2=0.475 $Y2=3.235
cc_48 N_VDD_c_48_p N_A0_M1000_g 0.00606474f $X=1.825 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_49 N_VDD_c_49_p N_A0_M1000_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.475 $Y2=3.235
cc_50 N_VDD_M1000_b N_A0_c_80_n 0.00545313f $X=-0.045 $Y=2.415 $X2=0.345
+ $Y2=2.11
cc_51 N_VDD_M1000_b N_A1_M1006_g 0.0210839f $X=-0.045 $Y=2.415 $X2=0.835
+ $Y2=3.235
cc_52 N_VDD_c_48_p N_A1_M1006_g 0.00606474f $X=1.825 $Y=4.287 $X2=0.835
+ $Y2=3.235
cc_53 N_VDD_c_49_p N_A1_M1006_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.835 $Y2=3.235
cc_54 N_VDD_M1000_b N_B0_M1005_g 0.0200941f $X=-0.045 $Y=2.415 $X2=1.335
+ $Y2=3.235
cc_55 N_VDD_c_48_p N_B0_M1005_g 0.00606474f $X=1.825 $Y=4.287 $X2=1.335
+ $Y2=3.235
cc_56 N_VDD_c_49_p N_B0_M1005_g 0.00468827f $X=1.7 $Y=4.25 $X2=1.335 $Y2=3.235
cc_57 N_VDD_M1000_b N_B0_c_142_n 0.00243756f $X=-0.045 $Y=2.415 $X2=1.2 $Y2=2.48
cc_58 N_VDD_M1000_b B0 0.00672004f $X=-0.045 $Y=2.415 $X2=1.2 $Y2=2.48
cc_59 N_VDD_M1000_b N_B1_c_193_n 0.0292218f $X=-0.045 $Y=2.415 $X2=1.695
+ $Y2=2.52
cc_60 N_VDD_c_48_p N_B1_c_193_n 0.00606474f $X=1.825 $Y=4.287 $X2=1.695 $Y2=2.52
cc_61 N_VDD_c_61_p N_B1_c_193_n 0.00542179f $X=1.91 $Y=3.35 $X2=1.695 $Y2=2.52
cc_62 N_VDD_c_49_p N_B1_c_193_n 0.00468827f $X=1.7 $Y=4.25 $X2=1.695 $Y2=2.52
cc_63 N_VDD_M1000_b N_Y_c_220_n 0.00156987f $X=-0.045 $Y=2.415 $X2=1.085
+ $Y2=3.01
cc_64 N_VDD_c_48_p N_Y_c_220_n 0.00738471f $X=1.825 $Y=4.287 $X2=1.085 $Y2=3.01
cc_65 N_VDD_c_49_p N_Y_c_220_n 0.00476747f $X=1.7 $Y=4.25 $X2=1.085 $Y2=3.01
cc_66 N_VDD_M1000_b N_Y_c_218_n 0.00106911f $X=-0.045 $Y=2.415 $X2=1.665
+ $Y2=1.74
cc_67 N_A0_c_67_n N_A1_M1006_g 0.0076084f $X=0.345 $Y=2.085 $X2=0.835 $Y2=3.235
cc_68 N_A0_c_72_n N_A1_M1006_g 0.113499f $X=0.475 $Y=2.445 $X2=0.835 $Y2=3.235
cc_69 N_A0_c_80_n N_A1_M1006_g 0.003633f $X=0.345 $Y=2.11 $X2=0.835 $Y2=3.235
cc_70 A0 N_A1_M1006_g 0.00372502f $X=0.345 $Y=2.11 $X2=0.835 $Y2=3.235
cc_71 N_A0_c_67_n N_A1_M1001_g 0.00779003f $X=0.345 $Y=2.085 $X2=0.905 $Y2=0.85
cc_72 N_A0_c_68_n N_A1_M1001_g 0.0255439f $X=0.475 $Y=1.23 $X2=0.905 $Y2=0.85
cc_73 N_A0_c_67_n N_A1_c_99_n 0.0168667f $X=0.345 $Y=2.085 $X2=0.815 $Y2=1.74
cc_74 N_A0_c_67_n N_A1_c_100_n 0.00347363f $X=0.345 $Y=2.085 $X2=0.815 $Y2=1.74
cc_75 N_A0_c_67_n A1 0.0012072f $X=0.345 $Y=2.085 $X2=0.815 $Y2=1.74
cc_76 A0 N_B0_c_142_n 0.00617211f $X=0.345 $Y=2.11 $X2=1.2 $Y2=2.48
cc_77 N_A0_c_80_n B0 0.0016426f $X=0.345 $Y=2.11 $X2=1.2 $Y2=2.48
cc_78 N_A0_c_68_n N_A_27_115#_c_262_n 0.0132289f $X=0.475 $Y=1.23 $X2=1.035
+ $Y2=1.16
cc_79 N_A0_c_73_n N_A_27_115#_c_262_n 0.00968589f $X=0.475 $Y=1.307 $X2=1.035
+ $Y2=1.16
cc_80 N_A0_c_73_n N_A_27_115#_c_265_n 0.00669281f $X=0.475 $Y=1.307 $X2=0.345
+ $Y2=1.16
cc_81 N_A1_M1001_g N_B0_M1002_g 0.037162f $X=0.905 $Y=0.85 $X2=1.335 $Y2=0.85
cc_82 N_A1_c_100_n N_B0_M1002_g 7.86889e-19 $X=0.815 $Y=1.74 $X2=1.335 $Y2=0.85
cc_83 A1 N_B0_M1002_g 2.44378e-19 $X=0.815 $Y=1.74 $X2=1.335 $Y2=0.85
cc_84 N_A1_M1006_g N_B0_M1005_g 0.0307551f $X=0.835 $Y=3.235 $X2=1.335 $Y2=3.235
cc_85 N_A1_M1006_g N_B0_c_141_n 0.00572826f $X=0.835 $Y=3.235 $X2=1.325 $Y2=1.85
cc_86 N_A1_c_99_n N_B0_c_141_n 0.0126055f $X=0.815 $Y=1.74 $X2=1.325 $Y2=1.85
cc_87 N_A1_c_100_n N_B0_c_141_n 3.07574e-19 $X=0.815 $Y=1.74 $X2=1.325 $Y2=1.85
cc_88 N_A1_M1006_g N_B0_c_142_n 0.0105014f $X=0.835 $Y=3.235 $X2=1.2 $Y2=2.48
cc_89 N_A1_M1006_g N_B0_c_143_n 0.00258968f $X=0.835 $Y=3.235 $X2=1.325 $Y2=1.85
cc_90 N_A1_c_99_n N_B0_c_143_n 0.00113642f $X=0.815 $Y=1.74 $X2=1.325 $Y2=1.85
cc_91 N_A1_c_100_n N_B0_c_143_n 0.011508f $X=0.815 $Y=1.74 $X2=1.325 $Y2=1.85
cc_92 A1 N_B0_c_143_n 0.00222079f $X=0.815 $Y=1.74 $X2=1.325 $Y2=1.85
cc_93 N_A1_M1006_g B0 0.00416458f $X=0.835 $Y=3.235 $X2=1.2 $Y2=2.48
cc_94 N_A1_c_99_n B0 7.13593e-19 $X=0.815 $Y=1.74 $X2=1.2 $Y2=2.48
cc_95 A1 B0 0.001519f $X=0.815 $Y=1.74 $X2=1.2 $Y2=2.48
cc_96 N_A1_M1006_g N_Y_c_224_n 0.00482048f $X=0.835 $Y=3.235 $X2=1.17 $Y2=2.83
cc_97 A1 N_Y_c_218_n 2.09357e-19 $X=0.815 $Y=1.74 $X2=1.665 $Y2=1.74
cc_98 N_A1_c_100_n Y 5.04816e-19 $X=0.815 $Y=1.74 $X2=1.665 $Y2=1.74
cc_99 A1 Y 0.014403f $X=0.815 $Y=1.74 $X2=1.665 $Y2=1.74
cc_100 N_A1_M1001_g N_A_27_115#_c_262_n 0.0151241f $X=0.905 $Y=0.85 $X2=1.035
+ $Y2=1.16
cc_101 N_A1_c_99_n N_A_27_115#_c_262_n 0.00299395f $X=0.815 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_102 N_A1_c_100_n N_A_27_115#_c_262_n 0.00670548f $X=0.815 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_103 A1 N_A_27_115#_c_262_n 0.00917137f $X=0.815 $Y=1.74 $X2=1.035 $Y2=1.16
cc_104 N_A1_M1001_g N_A_27_115#_c_268_n 5.22852e-19 $X=0.905 $Y=0.85 $X2=1.205
+ $Y2=0.63
cc_105 N_B0_M1005_g N_B1_c_193_n 0.111794f $X=1.335 $Y=3.235 $X2=1.695 $Y2=2.52
cc_106 N_B0_c_142_n N_B1_c_193_n 6.45943e-19 $X=1.2 $Y=2.48 $X2=1.695 $Y2=2.52
cc_107 N_B0_M1002_g N_B1_M1007_g 0.0386549f $X=1.335 $Y=0.85 $X2=1.765 $Y2=0.85
cc_108 N_B0_c_141_n N_B1_M1007_g 0.0187771f $X=1.325 $Y=1.85 $X2=1.765 $Y2=0.85
cc_109 N_B0_c_143_n N_B1_M1007_g 3.80244e-19 $X=1.325 $Y=1.85 $X2=1.765 $Y2=0.85
cc_110 N_B0_M1005_g N_Y_c_228_n 0.0153691f $X=1.335 $Y=3.235 $X2=1.58 $Y2=2.83
cc_111 N_B0_c_142_n N_Y_c_228_n 0.00536561f $X=1.2 $Y=2.48 $X2=1.58 $Y2=2.83
cc_112 B0 N_Y_c_228_n 0.00561823f $X=1.2 $Y=2.48 $X2=1.58 $Y2=2.83
cc_113 N_B0_c_142_n N_Y_c_224_n 0.00372626f $X=1.2 $Y=2.48 $X2=1.17 $Y2=2.83
cc_114 B0 N_Y_c_224_n 0.00791606f $X=1.2 $Y=2.48 $X2=1.17 $Y2=2.83
cc_115 N_B0_M1002_g N_Y_c_217_n 0.00584345f $X=1.335 $Y=0.85 $X2=1.665 $Y2=1.235
cc_116 N_B0_c_141_n N_Y_c_217_n 0.0012173f $X=1.325 $Y=1.85 $X2=1.665 $Y2=1.235
cc_117 N_B0_c_143_n N_Y_c_217_n 8.58442e-19 $X=1.325 $Y=1.85 $X2=1.665 $Y2=1.235
cc_118 N_B0_M1002_g N_Y_c_218_n 0.0089275f $X=1.335 $Y=0.85 $X2=1.665 $Y2=1.74
cc_119 N_B0_M1005_g N_Y_c_218_n 0.00482513f $X=1.335 $Y=3.235 $X2=1.665 $Y2=1.74
cc_120 N_B0_c_141_n N_Y_c_218_n 0.0018033f $X=1.325 $Y=1.85 $X2=1.665 $Y2=1.74
cc_121 N_B0_c_142_n N_Y_c_218_n 0.0223282f $X=1.2 $Y=2.48 $X2=1.665 $Y2=1.74
cc_122 N_B0_c_143_n N_Y_c_218_n 0.0233023f $X=1.325 $Y=1.85 $X2=1.665 $Y2=1.74
cc_123 B0 N_Y_c_218_n 0.00640554f $X=1.2 $Y=2.48 $X2=1.665 $Y2=1.74
cc_124 N_B0_M1002_g Y 4.29441e-19 $X=1.335 $Y=0.85 $X2=1.665 $Y2=1.74
cc_125 N_B0_c_141_n Y 0.00355451f $X=1.325 $Y=1.85 $X2=1.665 $Y2=1.74
cc_126 N_B0_c_143_n Y 0.00220294f $X=1.325 $Y=1.85 $X2=1.665 $Y2=1.74
cc_127 N_B0_M1002_g N_A_27_115#_c_262_n 0.00123589f $X=1.335 $Y=0.85 $X2=1.035
+ $Y2=1.16
cc_128 N_B0_c_141_n N_A_27_115#_c_262_n 2.93581e-19 $X=1.325 $Y=1.85 $X2=1.035
+ $Y2=1.16
cc_129 N_B0_c_143_n N_A_27_115#_c_262_n 0.00406274f $X=1.325 $Y=1.85 $X2=1.035
+ $Y2=1.16
cc_130 N_B0_M1002_g N_A_27_115#_c_266_n 0.0123082f $X=1.335 $Y=0.85 $X2=1.895
+ $Y2=0.63
cc_131 N_B1_c_193_n N_Y_c_228_n 0.0176551f $X=1.695 $Y=2.52 $X2=1.58 $Y2=2.83
cc_132 N_B1_M1007_g N_Y_c_217_n 0.0175045f $X=1.765 $Y=0.85 $X2=1.665 $Y2=1.235
cc_133 N_B1_c_193_n N_Y_c_218_n 0.0336478f $X=1.695 $Y=2.52 $X2=1.665 $Y2=1.74
cc_134 N_B1_M1007_g N_Y_c_218_n 0.0306339f $X=1.765 $Y=0.85 $X2=1.665 $Y2=1.74
cc_135 N_B1_c_196_n N_Y_c_218_n 0.0203078f $X=2.005 $Y=2.115 $X2=1.665 $Y2=1.74
cc_136 B1 N_Y_c_218_n 0.00704472f $X=2.005 $Y=2.115 $X2=1.665 $Y2=1.74
cc_137 N_B1_M1007_g Y 0.0119786f $X=1.765 $Y=0.85 $X2=1.665 $Y2=1.74
cc_138 B1 Y 0.00540133f $X=2.005 $Y=2.115 $X2=1.665 $Y2=1.74
cc_139 N_B1_M1007_g N_A_27_115#_c_266_n 0.0111266f $X=1.765 $Y=0.85 $X2=1.895
+ $Y2=0.63
cc_140 N_B1_M1007_g N_A_27_115#_c_271_n 2.59689e-19 $X=1.765 $Y=0.85 $X2=1.98
+ $Y2=0.63
cc_141 N_Y_c_228_n A_282_521# 0.00732587f $X=1.58 $Y=2.83 $X2=1.41 $Y2=2.605
cc_142 N_Y_c_217_n N_A_27_115#_c_262_n 0.0107797f $X=1.665 $Y=1.235 $X2=1.035
+ $Y2=1.16
cc_143 N_Y_c_218_n N_A_27_115#_c_262_n 4.63961e-19 $X=1.665 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_144 N_Y_M1002_d N_A_27_115#_c_266_n 0.00176461f $X=1.41 $Y=0.575 $X2=1.895
+ $Y2=0.63
cc_145 N_Y_c_217_n N_A_27_115#_c_266_n 0.0176852f $X=1.665 $Y=1.235 $X2=1.895
+ $Y2=0.63
