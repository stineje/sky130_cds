* File: sky130_osu_sc_12T_hs__buf_8.pex.spice
* Created: Fri Nov 12 15:08:36 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__BUF_8%GND 1 2 3 4 5 57 59 67 69 76 78 85 87 94
+ 96 104 115 117
r125 115 117 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r126 102 104 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.13 $Y=0.305
+ $X2=4.13 $Y2=0.755
r127 97 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.152
+ $X2=3.27 $Y2=0.152
r128 96 102 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.045 $Y=0.152
+ $X2=4.13 $Y2=0.305
r129 92 111 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.152
r130 92 94 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.755
r131 87 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.152
+ $X2=3.27 $Y2=0.152
r132 83 85 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.755
r133 79 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0.152
+ $X2=1.55 $Y2=0.152
r134 74 107 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.152
r135 74 76 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.755
r136 70 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r137 69 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.152
r138 65 106 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r139 65 67 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r140 59 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r141 57 117 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r142 57 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r143 57 83 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.41 $Y2=0.305
r144 57 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.325 $Y2=0.152
r145 57 88 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.495 $Y2=0.152
r146 57 96 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.045 $Y2=0.152
r147 57 97 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.355 $Y2=0.152
r148 57 87 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.185 $Y2=0.152
r149 57 88 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.495 $Y2=0.152
r150 57 78 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r151 57 79 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r152 57 69 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r153 57 70 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r154 57 59 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r155 5 104 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.755
r156 4 94 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.755
r157 3 85 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.755
r158 2 76 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
r159 1 67 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_8%VDD 1 2 3 4 5 45 47 54 56 62 66 72 76 82
+ 86 93 103 107
r82 103 107 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=3.74 $Y2=4.287
r83 93 96 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.13 $Y=2.955
+ $X2=4.13 $Y2=3.635
r84 91 96 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.13 $Y=4.135 $X2=4.13
+ $Y2=3.635
r85 89 107 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=4.25
+ $X2=3.74 $Y2=4.25
r86 87 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=4.287
+ $X2=3.27 $Y2=4.287
r87 87 89 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=3.355 $Y=4.287
+ $X2=3.74 $Y2=4.287
r88 86 91 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.045 $Y=4.287
+ $X2=4.13 $Y2=4.135
r89 86 89 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.045 $Y=4.287
+ $X2=3.74 $Y2=4.287
r90 82 85 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=2.955
+ $X2=3.27 $Y2=3.635
r91 80 101 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.27 $Y=4.135
+ $X2=3.27 $Y2=4.287
r92 80 85 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.27 $Y=4.135 $X2=3.27
+ $Y2=3.635
r93 77 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=4.287
+ $X2=2.41 $Y2=4.287
r94 77 79 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=2.495 $Y=4.287
+ $X2=3.06 $Y2=4.287
r95 76 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=4.287
+ $X2=3.27 $Y2=4.287
r96 76 79 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=4.287
+ $X2=3.06 $Y2=4.287
r97 72 75 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=2.955
+ $X2=2.41 $Y2=3.635
r98 70 100 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.41 $Y=4.135
+ $X2=2.41 $Y2=4.287
r99 70 75 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.41 $Y=4.135 $X2=2.41
+ $Y2=3.635
r100 67 98 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=4.287
+ $X2=1.55 $Y2=4.287
r101 67 69 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=4.287
+ $X2=1.7 $Y2=4.287
r102 66 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=4.287
+ $X2=2.41 $Y2=4.287
r103 66 69 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=4.287
+ $X2=1.7 $Y2=4.287
r104 62 65 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r105 60 98 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=4.287
r106 60 65 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=3.635
r107 57 97 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r108 57 59 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r109 56 98 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=4.287
+ $X2=1.55 $Y2=4.287
r110 56 59 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=4.287
+ $X2=1.02 $Y2=4.287
r111 52 97 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r112 52 54 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.635
r113 49 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r114 47 97 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r115 47 49 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r116 45 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r117 45 79 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r118 45 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r119 45 69 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r120 45 59 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r121 45 49 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r122 5 96 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.605 $X2=4.13 $Y2=3.635
r123 5 93 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.605 $X2=4.13 $Y2=2.955
r124 4 85 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=3.635
r125 4 82 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=2.955
r126 3 75 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=3.635
r127 3 72 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=2.955
r128 2 65 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r129 2 62 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r130 1 54 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_8%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=2.85
+ $X2=0.635 $Y2=2.85
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2 $X2=0.635
+ $Y2=2.85
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635 $Y=2
+ $X2=0.635 $Y2=2
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=2.165
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=1.835
r45 7 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=2.165
r46 3 11 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=0.475 $Y=0.85
+ $X2=0.475 $Y2=1.835
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_8%A_27_115# 1 3 11 13 15 17 20 22 24 25 26
+ 27 28 31 33 35 36 38 42 44 46 47 49 53 56 57 59 60 62 66 68 70 71 73 77 79 81
+ 82 84 88 90 92 102 103 104 105 106 107 108 109 110 111 114 118 122 124 127
c232 79 0 1.33323e-19 $X=3.485 $Y=2.53
c233 77 0 1.33323e-19 $X=3.485 $Y=0.85
c234 68 0 1.33323e-19 $X=3.055 $Y=2.53
c235 66 0 1.33323e-19 $X=3.055 $Y=0.85
c236 57 0 1.33323e-19 $X=2.625 $Y=2.53
c237 53 0 1.33323e-19 $X=2.625 $Y=0.85
c238 44 0 1.33323e-19 $X=2.195 $Y=2.53
c239 42 0 1.33323e-19 $X=2.195 $Y=0.85
c240 33 0 1.33323e-19 $X=1.765 $Y=2.53
c241 31 0 1.33323e-19 $X=1.765 $Y=0.85
c242 22 0 1.33323e-19 $X=1.335 $Y=2.53
c243 20 0 1.33323e-19 $X=1.335 $Y=0.85
r244 123 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.455
+ $X2=0.26 $Y2=1.455
r245 122 127 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.965 $Y2=1.455
r246 122 123 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.345 $Y2=1.455
r247 118 120 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r248 116 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.54
+ $X2=0.26 $Y2=1.455
r249 116 118 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=0.26 $Y=1.54
+ $X2=0.26 $Y2=2.955
r250 112 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=1.455
r251 112 114 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r252 99 127 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.455 $X2=0.965 $Y2=1.455
r253 99 100 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.455
+ $X2=1.18 $Y2=1.455
r254 97 99 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.455
+ $X2=0.965 $Y2=1.455
r255 95 96 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.455
+ $X2=1.335 $Y2=2.455
r256 93 95 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.455
+ $X2=1.18 $Y2=2.455
r257 90 92 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.915 $Y=2.53
+ $X2=3.915 $Y2=3.235
r258 86 88 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.915 $Y=1.29
+ $X2=3.915 $Y2=0.85
r259 85 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.455
+ $X2=3.485 $Y2=2.455
r260 84 90 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=2.455
+ $X2=3.915 $Y2=2.53
r261 84 85 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.455
+ $X2=3.56 $Y2=2.455
r262 83 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.365
+ $X2=3.485 $Y2=1.365
r263 82 86 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=1.365
+ $X2=3.915 $Y2=1.29
r264 82 83 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.365
+ $X2=3.56 $Y2=1.365
r265 79 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.53
+ $X2=3.485 $Y2=2.455
r266 79 81 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.485 $Y=2.53
+ $X2=3.485 $Y2=3.235
r267 75 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.29
+ $X2=3.485 $Y2=1.365
r268 75 77 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.485 $Y=1.29
+ $X2=3.485 $Y2=0.85
r269 74 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.455
+ $X2=3.055 $Y2=2.455
r270 73 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.455
+ $X2=3.485 $Y2=2.455
r271 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.455
+ $X2=3.13 $Y2=2.455
r272 72 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.365
+ $X2=3.055 $Y2=1.365
r273 71 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.365
+ $X2=3.485 $Y2=1.365
r274 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.365
+ $X2=3.13 $Y2=1.365
r275 68 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.53
+ $X2=3.055 $Y2=2.455
r276 68 70 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.055 $Y=2.53
+ $X2=3.055 $Y2=3.235
r277 64 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.29
+ $X2=3.055 $Y2=1.365
r278 64 66 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.055 $Y=1.29
+ $X2=3.055 $Y2=0.85
r279 63 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.455
+ $X2=2.625 $Y2=2.455
r280 62 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.455
+ $X2=3.055 $Y2=2.455
r281 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.455
+ $X2=2.7 $Y2=2.455
r282 61 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.365
+ $X2=2.625 $Y2=1.365
r283 60 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.365
+ $X2=3.055 $Y2=1.365
r284 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.365
+ $X2=2.7 $Y2=1.365
r285 57 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.53
+ $X2=2.625 $Y2=2.455
r286 57 59 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.625 $Y=2.53
+ $X2=2.625 $Y2=3.235
r287 56 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.38
+ $X2=2.625 $Y2=2.455
r288 55 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=1.365
r289 55 56 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.625 $Y=1.44 $X2=2.625
+ $Y2=2.38
r290 51 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.29
+ $X2=2.625 $Y2=1.365
r291 51 53 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.625 $Y=1.29
+ $X2=2.625 $Y2=0.85
r292 50 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.455
+ $X2=2.195 $Y2=2.455
r293 49 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.455
+ $X2=2.625 $Y2=2.455
r294 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.455
+ $X2=2.27 $Y2=2.455
r295 48 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.365
+ $X2=2.195 $Y2=1.365
r296 47 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.365
+ $X2=2.625 $Y2=1.365
r297 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.365
+ $X2=2.27 $Y2=1.365
r298 44 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.53
+ $X2=2.195 $Y2=2.455
r299 44 46 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.195 $Y=2.53
+ $X2=2.195 $Y2=3.235
r300 40 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=1.365
r301 40 42 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=0.85
r302 39 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.455
+ $X2=1.765 $Y2=2.455
r303 38 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.455
+ $X2=2.195 $Y2=2.455
r304 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.455
+ $X2=1.84 $Y2=2.455
r305 37 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.365
+ $X2=1.765 $Y2=1.365
r306 36 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=2.195 $Y2=1.365
r307 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=1.84 $Y2=1.365
r308 33 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.53
+ $X2=1.765 $Y2=2.455
r309 33 35 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.765 $Y=2.53
+ $X2=1.765 $Y2=3.235
r310 29 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=1.365
r311 29 31 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=0.85
r312 28 96 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.455
+ $X2=1.335 $Y2=2.455
r313 27 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.455
+ $X2=1.765 $Y2=2.455
r314 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.455
+ $X2=1.41 $Y2=2.455
r315 25 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.365
+ $X2=1.765 $Y2=1.365
r316 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.365
+ $X2=1.41 $Y2=1.365
r317 22 96 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.53
+ $X2=1.335 $Y2=2.455
r318 22 24 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.335 $Y=2.53
+ $X2=1.335 $Y2=3.235
r319 18 26 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.41 $Y2=1.365
r320 18 100 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.18 $Y2=1.455
r321 18 20 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.85
r322 17 95 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.38
+ $X2=1.18 $Y2=2.455
r323 16 100 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=1.455
r324 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=2.38
r325 13 93 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=2.455
r326 13 15 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=3.235
r327 9 97 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=1.455
r328 9 11 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=0.85
r329 3 120 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r330 3 118 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r331 1 114 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__BUF_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68 76
+ 82 89 90 92 94 96 99 100 101 102 103 105 106 107 108 109 110 111
c173 111 0 1.33323e-19 $X=3.7 $Y=2.365
c174 110 0 1.33323e-19 $X=3.7 $Y=1.115
c175 109 0 2.66647e-19 $X=2.985 $Y=2.48
c176 107 0 2.66647e-19 $X=2.985 $Y=1
c177 103 0 2.66647e-19 $X=2.125 $Y=2.48
c178 101 0 2.66647e-19 $X=2.125 $Y=1
c179 90 0 1.33323e-19 $X=1.12 $Y=2.365
c180 89 0 1.33323e-19 $X=1.12 $Y=1.115
r181 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.7 $Y=2.365
+ $X2=3.7 $Y2=2.48
r182 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.7 $Y=1.115
+ $X2=3.7 $Y2=1
r183 110 111 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.7 $Y=1.115
+ $X2=3.7 $Y2=2.365
r184 109 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=2.48
+ $X2=2.84 $Y2=2.48
r185 108 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.555 $Y=2.48
+ $X2=3.7 $Y2=2.48
r186 108 109 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.555 $Y=2.48
+ $X2=2.985 $Y2=2.48
r187 107 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=1
+ $X2=2.84 $Y2=1
r188 106 125 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.555 $Y=1
+ $X2=3.7 $Y2=1
r189 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.555 $Y=1
+ $X2=2.985 $Y2=1
r190 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=2.365
+ $X2=2.84 $Y2=2.48
r191 104 121 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=1.115
+ $X2=2.84 $Y2=1
r192 104 105 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.84 $Y=1.115
+ $X2=2.84 $Y2=2.365
r193 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=2.48
+ $X2=1.98 $Y2=2.48
r194 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.48
+ $X2=2.84 $Y2=2.48
r195 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=2.48
+ $X2=2.125 $Y2=2.48
r196 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=1
+ $X2=1.98 $Y2=1
r197 100 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=1
+ $X2=2.84 $Y2=1
r198 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=1
+ $X2=2.125 $Y2=1
r199 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.365
+ $X2=1.98 $Y2=2.48
r200 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.115
+ $X2=1.98 $Y2=1
r201 98 99 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.115
+ $X2=1.98 $Y2=2.365
r202 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.48
+ $X2=1.12 $Y2=2.48
r203 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.48
+ $X2=1.98 $Y2=2.48
r204 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.48
+ $X2=1.265 $Y2=2.48
r205 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1
+ $X2=1.12 $Y2=1
r206 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1
+ $X2=1.98 $Y2=1
r207 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1
+ $X2=1.265 $Y2=1
r208 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=2.48
r209 90 92 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=1.79
r210 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1
r211 89 92 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1.79
r212 85 87 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=2.955
+ $X2=3.7 $Y2=3.635
r213 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=2.48
+ $X2=3.7 $Y2=2.48
r214 82 85 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.7 $Y=2.48
+ $X2=3.7 $Y2=2.955
r215 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=1 $X2=3.7
+ $Y2=1
r216 76 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.7 $Y=0.755
+ $X2=3.7 $Y2=1
r217 71 73 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=2.955
+ $X2=2.84 $Y2=3.635
r218 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=2.48
+ $X2=2.84 $Y2=2.48
r219 68 71 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.84 $Y=2.48
+ $X2=2.84 $Y2=2.955
r220 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=1 $X2=2.84
+ $Y2=1
r221 62 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.84 $Y=0.755
+ $X2=2.84 $Y2=1
r222 57 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r223 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.48
+ $X2=1.98 $Y2=2.48
r224 54 57 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.98 $Y=2.48
+ $X2=1.98 $Y2=2.955
r225 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1 $X2=1.98
+ $Y2=1
r226 48 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.98 $Y=0.755
+ $X2=1.98 $Y2=1
r227 43 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r228 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.48
r229 40 43 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.955
r230 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1 $X2=1.12
+ $Y2=1
r231 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.12 $Y=0.755
+ $X2=1.12 $Y2=1
r232 12 87 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=3.635
r233 12 85 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=2.955
r234 11 73 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=3.635
r235 11 71 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=2.955
r236 10 59 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r237 10 57 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r238 9 45 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r239 9 43 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r240 4 76 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.755
r241 3 62 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.7 $Y=0.575
+ $X2=2.84 $Y2=0.755
r242 2 48 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.755
r243 1 34 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.755
.ends

