* File: sky130_osu_sc_15T_ms__buf_4.spice
* Created: Fri Nov 12 14:41:38 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__buf_4.pex.spice"
.subckt sky130_osu_sc_15T_ms__buf_4  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_A_M1006_g N_A_27_115#_M1006_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1006_d N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1001_d N_A_27_115#_M1003_g N_GND_M1003_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_A_27_115#_M1008_g N_GND_M1003_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1008_d N_A_27_115#_M1009_g N_GND_M1009_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VDD_M1007_d N_A_M1007_g N_A_27_115#_M1007_s N_VDD_M1007_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001.9 A=0.3 P=4.3 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_VDD_M1007_d N_VDD_M1007_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75001.5 A=0.3 P=4.3 MULT=1
MM1002 N_Y_M1000_d N_A_27_115#_M1002_g N_VDD_M1002_s N_VDD_M1007_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1004 N_Y_M1004_d N_A_27_115#_M1004_g N_VDD_M1002_s N_VDD_M1007_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001.5
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1005 N_Y_M1004_d N_A_27_115#_M1005_g N_VDD_M1005_s N_VDD_M1007_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75001.9
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX10_noxref N_GND_M1006_b N_VDD_M1007_b NWDIODE A=8.27475 P=11.51
pX11_noxref noxref_6 A A PROBETYPE=1
pX12_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__buf_4.pxi.spice"
*
.ends
*
*
