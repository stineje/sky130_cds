* File: sky130_osu_sc_12T_ls__aoi22_l.pex.spice
* Created: Fri Nov 12 15:34:49 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%GND 1 2 27 31 33 44 56 58
c47 27 0 6.36774e-20 $X=-0.045 $Y=0
r48 56 58 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r49 42 52 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.152
r50 42 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.755
r51 33 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=0.152
+ $X2=1.91 $Y2=0.152
r52 29 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r53 27 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r54 27 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r55 27 29 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r56 27 34 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r57 27 33 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.825 $Y2=0.152
r58 27 34 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r59 2 44 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.77 $Y=0.575
+ $X2=1.91 $Y2=0.755
r60 1 31 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%VDD 1 17 19 26 32 37 41
r29 37 41 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.7 $Y2=4.287
r30 32 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=4.25 $X2=1.7
+ $Y2=4.25
r31 30 32 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r32 28 35 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r33 28 30 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r34 24 35 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r35 24 26 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.655
r36 21 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r37 19 35 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r38 19 21 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r39 17 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r40 17 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r41 17 21 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r42 1 26 600 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.655
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%A0 2 3 5 8 12 18 21 27
c33 21 0 1.36621e-19 $X=0.385 $Y=2.11
c34 8 0 6.36774e-20 $X=0.475 $Y=3.235
r35 21 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=2.11
+ $X2=0.385 $Y2=2.11
r36 21 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.385 $Y=2.11
+ $X2=0.385 $Y2=2.285
r37 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.285 $X2=0.385 $Y2=2.285
r38 17 18 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.285
+ $X2=0.475 $Y2=2.285
r39 14 17 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.285
+ $X2=0.385 $Y2=2.285
r40 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.29
+ $X2=0.475 $Y2=1.29
r41 6 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.42
+ $X2=0.475 $Y2=2.285
r42 6 8 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=0.475 $Y=2.42
+ $X2=0.475 $Y2=3.235
r43 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.21 $X2=0.475
+ $Y2=1.29
r44 3 5 120.5 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.475 $Y=1.21 $X2=0.475
+ $Y2=0.835
r45 2 14 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.15
+ $X2=0.295 $Y2=2.285
r46 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.37 $X2=0.295
+ $Y2=1.29
r47 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.37
+ $X2=0.295 $Y2=2.15
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%A1 3 5 7 12 18
c44 5 0 1.36621e-19 $X=0.905 $Y=2.09
r45 15 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.48
+ $X2=0.725 $Y2=2.48
r46 12 15 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.725 $Y=1.775
+ $X2=0.725 $Y2=2.48
r47 10 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.775 $X2=0.725 $Y2=1.775
r48 5 10 63.0864 $w=2.95e-07 $l=3.7229e-07 $layer=POLY_cond $X=0.905 $Y=2.09
+ $X2=0.78 $Y2=1.775
r49 5 7 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=0.905 $Y=2.09
+ $X2=0.905 $Y2=3.235
r50 1 10 38.578 $w=2.95e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.835 $Y=1.61
+ $X2=0.78 $Y2=1.775
r51 1 3 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=0.835 $Y=1.61
+ $X2=0.835 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%B0 3 7 10 15 17 21
c42 3 0 1.94783e-19 $X=1.335 $Y=0.835
r43 17 19 3.63576 $w=3.02e-07 $l=9e-08 $layer=LI1_cond $X=1.165 $Y=1.42
+ $X2=1.255 $Y2=1.42
r44 15 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.11
+ $X2=1.165 $Y2=2.11
r45 13 17 4.10007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=1.585
+ $X2=1.165 $Y2=1.42
r46 13 15 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.165 $Y=1.585
+ $X2=1.165 $Y2=2.11
r47 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.42 $X2=1.255 $Y2=1.42
r48 10 12 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.42
+ $X2=1.265 $Y2=1.585
r49 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.42
+ $X2=1.265 $Y2=1.255
r50 7 12 846.064 $w=1.5e-07 $l=1.65e-06 $layer=POLY_cond $X=1.335 $Y=3.235
+ $X2=1.335 $Y2=1.585
r51 3 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.335 $Y=0.835
+ $X2=1.335 $Y2=1.255
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%B1 3 7 10 14 19
r26 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.935 $Y=1.74
+ $X2=1.935 $Y2=1.74
r27 12 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.74 $X2=1.935 $Y2=1.74
r28 10 12 26.0955 $w=3.14e-07 $l=1.7e-07 $layer=POLY_cond $X=1.765 $Y=1.722
+ $X2=1.935 $Y2=1.722
r29 9 10 10.7452 $w=3.14e-07 $l=7e-08 $layer=POLY_cond $X=1.695 $Y=1.722
+ $X2=1.765 $Y2=1.722
r30 5 10 20.044 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=1.765 $Y=1.905
+ $X2=1.765 $Y2=1.722
r31 5 7 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.765 $Y=1.905
+ $X2=1.765 $Y2=3.235
r32 1 9 20.044 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=1.695 $Y=1.54
+ $X2=1.695 $Y2=1.722
r33 1 3 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.695 $Y=1.54 $X2=1.695
+ $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%A_27_521# 1 2 3 15 17 18 23 24
r23 25 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.98 $Y=3.74
+ $X2=1.98 $Y2=3.49
r24 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.895 $Y=3.825
+ $X2=1.98 $Y2=3.74
r25 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=3.825
+ $X2=1.205 $Y2=3.825
r26 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=3.74
+ $X2=1.205 $Y2=3.825
r27 20 22 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.12 $Y=3.74
+ $X2=1.12 $Y2=3.485
r28 19 22 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.12 $Y=3.23
+ $X2=1.12 $Y2=3.485
r29 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.145
+ $X2=1.12 $Y2=3.23
r30 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.145
+ $X2=0.345 $Y2=3.145
r31 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.23
+ $X2=0.345 $Y2=3.145
r32 13 15 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=3.23
+ $X2=0.26 $Y2=3.485
r33 3 27 600 $w=1.7e-07 $l=9.52431e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.49
r34 2 22 600 $w=1.7e-07 $l=9.47418e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.485
r35 1 15 600 $w=1.7e-07 $l=9.40425e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.485
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AOI22_L%Y 1 3 10 17 21 25 26 30 36
c41 30 0 5.84789e-20 $X=1.605 $Y=1.22
c42 26 0 1.94783e-19 $X=1.23 $Y=1
r43 36 37 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.595 $Y=1.37
+ $X2=1.595 $Y2=1.255
r44 30 37 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.605 $Y=1.22
+ $X2=1.605 $Y2=1.255
r45 27 30 0.129989 $w=1.7e-07 $l=1.35e-07 $layer=MET1_cond $X=1.605 $Y=1.085
+ $X2=1.605 $Y2=1.22
r46 26 33 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.23 $Y=1
+ $X2=1.085 $Y2=1
r47 25 27 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.52 $Y=1
+ $X2=1.605 $Y2=1.085
r48 25 26 0.279236 $w=1.7e-07 $l=2.9e-07 $layer=MET1_cond $X=1.52 $Y=1 $X2=1.23
+ $Y2=1
r49 23 24 9.11234 $w=2.13e-07 $l=1.7e-07 $layer=LI1_cond $X=1.572 $Y=2.68
+ $X2=1.572 $Y2=2.85
r50 21 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.595 $Y=1.37
+ $X2=1.595 $Y2=1.37
r51 21 23 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.595 $Y=1.37
+ $X2=1.595 $Y2=2.68
r52 17 24 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.55 $Y=3.315
+ $X2=1.55 $Y2=2.85
r53 13 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=1 $X2=1.085
+ $Y2=1
r54 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.085 $Y=0.755
+ $X2=1.085 $Y2=1
r55 3 17 600 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.315
r56 1 10 182 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.085 $Y2=0.755
.ends

