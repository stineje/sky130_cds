* File: sky130_osu_sc_15T_ls__oai22_l.spice
* Created: Fri Nov 12 14:59:03 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__oai22_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__oai22_l  GND VDD A0 A1 B0 B1 Y
* 
* Y	Y
* B1	B1
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1005 N_GND_M1005_d N_A0_M1005_g N_A_27_115#_M1005_s N_GND_M1005_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_115#_M1000_d N_A1_M1000_g N_GND_M1005_d N_GND_M1005_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_115#_M1000_d N_GND_M1005_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_115#_M1006_d N_B1_M1006_g N_Y_M1002_d N_GND_M1005_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_110_565# N_A0_M1001_g N_VDD_M1001_s N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001.4 A=0.3 P=4.3 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g A_110_565# N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.35 AS=0.21 PD=2.35 PS=2.21 NRD=3.4278 NRS=4.9053 M=1 R=13.3333 SA=75000.5
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1003 A_282_565# N_B0_M1003_g N_Y_M1007_d N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.21 AS=0.35 PD=2.21 PS=2.35 NRD=4.9053 NRS=3.4278 M=1 R=13.3333 SA=75001
+ SB=75000.5 A=0.3 P=4.3 MULT=1
MM1004 N_VDD_M1004_d N_B1_M1004_g A_282_565# N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.53 AS=0.21 PD=4.53 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001.4
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX8_noxref N_GND_M1005_b N_VDD_M1001_b NWDIODE A=6.94725 P=10.61
pX9_noxref noxref_11 A0 A0 PROBETYPE=1
pX10_noxref noxref_12 A1 A1 PROBETYPE=1
pX11_noxref noxref_13 B0 B0 PROBETYPE=1
pX12_noxref noxref_14 Y Y PROBETYPE=1
pX13_noxref noxref_15 B1 B1 PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__oai22_l.pxi.spice"
*
.ends
*
*
