magic
tech sky130A
magscale 1 2
timestamp 1612372967
<< nwell >>
rect -10 529 1917 1119
<< nmoslvt >>
rect 80 115 110 243
rect 270 115 300 199
rect 356 115 386 199
rect 546 115 576 243
rect 618 115 648 243
rect 738 115 768 243
rect 810 115 840 243
rect 896 115 926 243
rect 968 115 998 243
rect 1088 115 1118 243
rect 1160 115 1190 243
rect 1246 115 1276 243
rect 1436 115 1466 199
rect 1522 115 1552 199
rect 1712 115 1742 243
rect 1798 115 1828 243
<< pmos >>
rect 80 565 110 965
rect 270 713 300 965
rect 342 713 372 965
rect 546 565 576 965
rect 618 565 648 965
rect 738 565 768 965
rect 810 565 840 965
rect 896 565 926 965
rect 968 565 998 965
rect 1088 565 1118 965
rect 1160 565 1190 965
rect 1246 565 1276 965
rect 1436 713 1466 965
rect 1508 713 1538 965
rect 1712 565 1742 965
rect 1798 565 1828 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 163 243
rect 110 131 121 215
rect 155 131 163 215
rect 493 215 546 243
rect 110 115 163 131
rect 217 165 270 199
rect 217 131 225 165
rect 259 131 270 165
rect 217 115 270 131
rect 300 165 356 199
rect 300 131 311 165
rect 345 131 356 165
rect 300 115 356 131
rect 386 165 439 199
rect 386 131 397 165
rect 431 131 439 165
rect 386 115 439 131
rect 493 131 501 215
rect 535 131 546 215
rect 493 115 546 131
rect 576 115 618 243
rect 648 215 738 243
rect 648 131 659 215
rect 727 131 738 215
rect 648 115 738 131
rect 768 115 810 243
rect 840 165 896 243
rect 840 131 851 165
rect 885 131 896 165
rect 840 115 896 131
rect 926 115 968 243
rect 998 215 1088 243
rect 998 131 1009 215
rect 1077 131 1088 215
rect 998 115 1088 131
rect 1118 115 1160 243
rect 1190 215 1246 243
rect 1190 131 1201 215
rect 1235 131 1246 215
rect 1190 115 1246 131
rect 1276 215 1329 243
rect 1276 131 1287 215
rect 1321 131 1329 215
rect 1276 115 1329 131
rect 1383 165 1436 199
rect 1383 131 1391 165
rect 1425 131 1436 165
rect 1383 115 1436 131
rect 1466 165 1522 199
rect 1466 131 1477 165
rect 1511 131 1522 165
rect 1466 115 1522 131
rect 1552 165 1605 199
rect 1552 131 1563 165
rect 1597 131 1605 165
rect 1552 115 1605 131
rect 1659 165 1712 243
rect 1659 131 1667 165
rect 1701 131 1712 165
rect 1659 115 1712 131
rect 1742 165 1798 243
rect 1742 131 1753 165
rect 1787 131 1798 165
rect 1742 115 1798 131
rect 1828 165 1881 243
rect 1828 131 1839 165
rect 1873 131 1881 165
rect 1828 115 1881 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 949 163 965
rect 110 605 121 949
rect 155 605 163 949
rect 217 949 270 965
rect 217 809 225 949
rect 259 809 270 949
rect 217 713 270 809
rect 300 713 342 965
rect 372 949 425 965
rect 372 809 383 949
rect 417 809 425 949
rect 372 713 425 809
rect 493 949 546 965
rect 110 565 163 605
rect 493 673 501 949
rect 535 673 546 949
rect 493 565 546 673
rect 576 565 618 965
rect 648 949 738 965
rect 648 605 659 949
rect 727 605 738 949
rect 648 565 738 605
rect 768 565 810 965
rect 840 949 896 965
rect 840 673 851 949
rect 885 673 896 949
rect 840 565 896 673
rect 926 565 968 965
rect 998 949 1088 965
rect 998 673 1009 949
rect 1077 673 1088 949
rect 998 565 1088 673
rect 1118 565 1160 965
rect 1190 949 1246 965
rect 1190 605 1201 949
rect 1235 605 1246 949
rect 1190 565 1246 605
rect 1276 949 1329 965
rect 1276 605 1287 949
rect 1321 605 1329 949
rect 1383 949 1436 965
rect 1383 809 1391 949
rect 1425 809 1436 949
rect 1383 713 1436 809
rect 1466 713 1508 965
rect 1538 949 1591 965
rect 1538 809 1549 949
rect 1583 809 1591 949
rect 1538 713 1591 809
rect 1659 949 1712 965
rect 1659 809 1667 949
rect 1701 809 1712 949
rect 1276 565 1329 605
rect 1659 565 1712 809
rect 1742 949 1798 965
rect 1742 809 1753 949
rect 1787 809 1798 949
rect 1742 565 1798 809
rect 1828 949 1881 965
rect 1828 809 1839 949
rect 1873 809 1881 949
rect 1828 565 1881 809
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 225 131 259 165
rect 311 131 345 165
rect 397 131 431 165
rect 501 131 535 215
rect 659 131 727 215
rect 851 131 885 165
rect 1009 131 1077 215
rect 1201 131 1235 215
rect 1287 131 1321 215
rect 1391 131 1425 165
rect 1477 131 1511 165
rect 1563 131 1597 165
rect 1667 131 1701 165
rect 1753 131 1787 165
rect 1839 131 1873 165
<< pdiffc >>
rect 35 741 69 949
rect 121 605 155 949
rect 225 809 259 949
rect 383 809 417 949
rect 501 673 535 949
rect 659 605 727 949
rect 851 673 885 949
rect 1009 673 1077 949
rect 1201 605 1235 949
rect 1287 605 1321 949
rect 1391 809 1425 949
rect 1549 809 1583 949
rect 1667 809 1701 949
rect 1753 809 1787 949
rect 1839 809 1873 949
<< psubdiff >>
rect 26 27 50 61
rect 84 27 108 61
rect 162 27 186 61
rect 220 27 244 61
rect 298 27 322 61
rect 356 27 380 61
rect 434 27 458 61
rect 492 27 516 61
rect 570 27 594 61
rect 628 27 652 61
rect 706 27 730 61
rect 764 27 788 61
rect 842 27 866 61
rect 900 27 924 61
rect 978 27 1002 61
rect 1036 27 1060 61
rect 1114 27 1138 61
rect 1172 27 1196 61
rect 1250 27 1274 61
rect 1308 27 1332 61
rect 1386 27 1410 61
rect 1444 27 1468 61
rect 1522 27 1546 61
rect 1580 27 1604 61
rect 1658 27 1682 61
rect 1716 27 1740 61
rect 1794 27 1818 61
rect 1852 27 1876 61
<< nsubdiff >>
rect 26 1049 50 1083
rect 84 1049 108 1083
rect 162 1049 186 1083
rect 220 1049 244 1083
rect 298 1049 322 1083
rect 356 1049 380 1083
rect 434 1049 458 1083
rect 492 1049 516 1083
rect 570 1049 594 1083
rect 628 1049 652 1083
rect 706 1049 730 1083
rect 764 1049 788 1083
rect 842 1049 866 1083
rect 900 1049 924 1083
rect 978 1049 1002 1083
rect 1036 1049 1060 1083
rect 1114 1049 1138 1083
rect 1172 1049 1196 1083
rect 1250 1049 1274 1083
rect 1308 1049 1332 1083
rect 1386 1049 1410 1083
rect 1444 1049 1468 1083
rect 1522 1049 1546 1083
rect 1580 1049 1604 1083
rect 1658 1049 1682 1083
rect 1716 1049 1740 1083
rect 1794 1049 1818 1083
rect 1852 1049 1876 1083
<< psubdiffcont >>
rect 50 27 84 61
rect 186 27 220 61
rect 322 27 356 61
rect 458 27 492 61
rect 594 27 628 61
rect 730 27 764 61
rect 866 27 900 61
rect 1002 27 1036 61
rect 1138 27 1172 61
rect 1274 27 1308 61
rect 1410 27 1444 61
rect 1546 27 1580 61
rect 1682 27 1716 61
rect 1818 27 1852 61
<< nsubdiffcont >>
rect 50 1049 84 1083
rect 186 1049 220 1083
rect 322 1049 356 1083
rect 458 1049 492 1083
rect 594 1049 628 1083
rect 730 1049 764 1083
rect 866 1049 900 1083
rect 1002 1049 1036 1083
rect 1138 1049 1172 1083
rect 1274 1049 1308 1083
rect 1410 1049 1444 1083
rect 1546 1049 1580 1083
rect 1682 1049 1716 1083
rect 1818 1049 1852 1083
<< poly >>
rect 80 965 110 991
rect 270 965 300 991
rect 342 965 372 991
rect 546 965 576 991
rect 618 965 648 991
rect 738 965 768 991
rect 810 965 840 991
rect 896 965 926 991
rect 968 965 998 991
rect 1088 965 1118 991
rect 1160 965 1190 991
rect 1246 965 1276 991
rect 1436 965 1466 991
rect 1508 965 1538 991
rect 1712 965 1742 991
rect 1798 965 1828 991
rect 80 442 110 565
rect 79 426 133 442
rect 79 392 89 426
rect 123 392 133 426
rect 79 376 133 392
rect 79 375 110 376
rect 80 243 110 375
rect 270 307 300 713
rect 342 532 372 713
rect 342 516 415 532
rect 342 482 371 516
rect 405 482 415 516
rect 342 466 415 482
rect 219 291 300 307
rect 219 257 229 291
rect 263 257 300 291
rect 219 241 300 257
rect 270 199 300 241
rect 356 199 386 466
rect 546 425 576 565
rect 618 534 648 565
rect 618 518 672 534
rect 618 484 628 518
rect 662 484 672 518
rect 618 468 672 484
rect 546 409 600 425
rect 738 423 768 565
rect 810 528 840 565
rect 896 528 926 565
rect 810 518 926 528
rect 810 484 842 518
rect 876 484 926 518
rect 810 474 926 484
rect 968 423 998 565
rect 1088 534 1118 565
rect 1064 518 1118 534
rect 1064 484 1074 518
rect 1108 484 1118 518
rect 1064 468 1118 484
rect 546 375 556 409
rect 590 375 600 409
rect 546 359 600 375
rect 642 393 1094 423
rect 546 243 576 359
rect 642 315 672 393
rect 1064 351 1094 393
rect 1160 419 1190 565
rect 1246 534 1276 565
rect 1246 518 1317 534
rect 1246 504 1273 518
rect 1257 484 1273 504
rect 1307 484 1317 518
rect 1257 468 1317 484
rect 1160 403 1214 419
rect 1160 369 1170 403
rect 1204 369 1214 403
rect 1160 353 1214 369
rect 618 285 672 315
rect 714 335 768 351
rect 714 301 724 335
rect 758 301 768 335
rect 714 285 768 301
rect 618 243 648 285
rect 738 243 768 285
rect 810 335 926 345
rect 810 301 842 335
rect 876 301 926 335
rect 810 291 926 301
rect 810 243 840 291
rect 896 243 926 291
rect 968 335 1022 351
rect 968 301 978 335
rect 1012 301 1022 335
rect 968 285 1022 301
rect 1064 335 1118 351
rect 1064 301 1074 335
rect 1108 301 1118 335
rect 1064 285 1118 301
rect 968 243 998 285
rect 1088 243 1118 285
rect 1160 243 1190 353
rect 1257 315 1287 468
rect 1436 351 1466 713
rect 1246 285 1287 315
rect 1399 335 1466 351
rect 1399 301 1409 335
rect 1443 301 1466 335
rect 1399 285 1466 301
rect 1246 243 1276 285
rect 1423 284 1466 285
rect 1436 199 1466 284
rect 1508 307 1538 713
rect 1712 549 1742 565
rect 1702 519 1742 549
rect 1702 419 1732 519
rect 1798 460 1828 565
rect 1677 403 1732 419
rect 1677 369 1687 403
rect 1721 369 1732 403
rect 1774 444 1828 460
rect 1774 410 1784 444
rect 1818 410 1828 444
rect 1774 394 1828 410
rect 1677 353 1732 369
rect 1702 308 1732 353
rect 1508 291 1589 307
rect 1508 257 1545 291
rect 1579 257 1589 291
rect 1702 278 1742 308
rect 1508 241 1589 257
rect 1712 243 1742 278
rect 1798 243 1828 394
rect 1522 199 1552 241
rect 80 89 110 115
rect 270 89 300 115
rect 356 89 386 115
rect 546 89 576 115
rect 618 89 648 115
rect 738 89 768 115
rect 810 89 840 115
rect 896 89 926 115
rect 968 89 998 115
rect 1088 89 1118 115
rect 1160 89 1190 115
rect 1246 89 1276 115
rect 1436 89 1466 115
rect 1522 89 1552 115
rect 1712 89 1742 115
rect 1798 89 1828 115
<< polycont >>
rect 89 392 123 426
rect 371 482 405 516
rect 229 257 263 291
rect 628 484 662 518
rect 842 484 876 518
rect 1074 484 1108 518
rect 556 375 590 409
rect 1273 484 1307 518
rect 1170 369 1204 403
rect 724 301 758 335
rect 842 301 876 335
rect 978 301 1012 335
rect 1074 301 1108 335
rect 1409 301 1443 335
rect 1687 369 1721 403
rect 1784 410 1818 444
rect 1545 257 1579 291
<< locali >>
rect 0 1089 1914 1110
rect 0 1049 50 1089
rect 84 1049 186 1089
rect 220 1049 322 1089
rect 356 1049 458 1089
rect 492 1049 594 1089
rect 628 1049 730 1089
rect 764 1049 866 1089
rect 900 1049 1002 1089
rect 1036 1049 1138 1089
rect 1172 1049 1274 1089
rect 1308 1049 1410 1089
rect 1444 1049 1546 1089
rect 1580 1049 1682 1089
rect 1716 1049 1818 1089
rect 1852 1049 1914 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 121 949 155 965
rect 47 442 81 597
rect 121 513 155 605
rect 225 949 259 965
rect 121 479 191 513
rect 47 426 123 442
rect 47 392 89 426
rect 89 376 123 392
rect 157 291 191 479
rect 225 375 259 809
rect 383 949 417 1049
rect 383 793 417 809
rect 501 949 535 1049
rect 501 657 535 673
rect 659 949 727 965
rect 851 949 885 1049
rect 851 657 885 673
rect 1009 949 1077 965
rect 659 602 727 605
rect 1009 602 1077 673
rect 405 568 727 602
rect 910 568 1077 602
rect 1201 949 1235 1049
rect 1201 589 1235 605
rect 1287 949 1321 965
rect 1391 949 1425 965
rect 1391 721 1425 809
rect 1549 949 1583 1049
rect 1549 793 1583 809
rect 1667 949 1701 965
rect 1391 687 1511 721
rect 1287 602 1321 605
rect 1287 568 1377 602
rect 405 532 439 568
rect 371 516 439 532
rect 405 482 439 516
rect 371 466 439 482
rect 225 341 345 375
rect 311 335 345 341
rect 229 291 263 307
rect 121 257 229 291
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 257
rect 121 115 155 131
rect 225 165 259 181
rect 225 61 259 131
rect 311 165 345 301
rect 405 318 439 466
rect 628 518 662 534
rect 628 483 662 484
rect 842 518 876 534
rect 662 449 758 483
rect 556 409 590 425
rect 556 359 590 375
rect 724 335 758 449
rect 842 335 876 484
rect 405 284 690 318
rect 724 285 758 301
rect 842 285 876 301
rect 910 335 944 568
rect 1074 518 1108 534
rect 1074 483 1108 484
rect 656 231 690 284
rect 910 251 944 301
rect 978 449 1074 483
rect 1273 518 1307 534
rect 1273 483 1307 484
rect 978 335 1012 449
rect 1341 403 1377 568
rect 1154 369 1170 403
rect 1204 369 1220 403
rect 1287 369 1377 403
rect 1477 403 1511 687
rect 1667 557 1701 809
rect 1753 949 1787 1049
rect 1753 793 1787 809
rect 1839 949 1873 965
rect 1839 631 1873 809
rect 1872 614 1873 631
rect 1872 597 1896 614
rect 1839 580 1896 597
rect 1667 518 1701 523
rect 1667 484 1818 518
rect 1784 444 1818 484
rect 1477 369 1687 403
rect 1721 369 1737 403
rect 1287 335 1321 369
rect 1058 301 1074 335
rect 1108 301 1321 335
rect 978 285 1012 301
rect 501 215 535 231
rect 311 115 345 131
rect 397 165 431 181
rect 397 61 431 131
rect 656 215 727 231
rect 910 217 1077 251
rect 656 197 659 215
rect 501 61 535 131
rect 1009 215 1077 217
rect 659 115 727 131
rect 851 165 885 181
rect 851 61 885 131
rect 1009 115 1077 131
rect 1201 215 1235 231
rect 1201 61 1235 131
rect 1287 215 1321 301
rect 1409 335 1443 351
rect 1409 285 1443 301
rect 1287 115 1321 131
rect 1391 165 1425 181
rect 1391 61 1425 131
rect 1477 165 1511 369
rect 1784 335 1818 410
rect 1545 291 1579 307
rect 1667 301 1818 335
rect 1477 115 1511 131
rect 1563 165 1597 181
rect 1563 61 1597 131
rect 1667 165 1701 301
rect 1862 268 1896 580
rect 1839 234 1896 268
rect 1667 115 1701 131
rect 1753 165 1787 181
rect 1753 61 1787 131
rect 1839 165 1873 234
rect 1839 115 1873 131
rect 0 21 50 61
rect 84 21 186 61
rect 220 21 322 61
rect 356 21 458 61
rect 492 21 594 61
rect 628 21 730 61
rect 764 21 866 61
rect 900 21 1002 61
rect 1036 21 1138 61
rect 1172 21 1274 61
rect 1308 21 1410 61
rect 1444 21 1546 61
rect 1580 21 1682 61
rect 1716 21 1818 61
rect 1852 21 1914 61
rect 0 0 1914 21
<< viali >>
rect 50 1083 84 1089
rect 50 1055 84 1083
rect 186 1083 220 1089
rect 186 1055 220 1083
rect 322 1083 356 1089
rect 322 1055 356 1083
rect 458 1083 492 1089
rect 458 1055 492 1083
rect 594 1083 628 1089
rect 594 1055 628 1083
rect 730 1083 764 1089
rect 730 1055 764 1083
rect 866 1083 900 1089
rect 866 1055 900 1083
rect 1002 1083 1036 1089
rect 1002 1055 1036 1083
rect 1138 1083 1172 1089
rect 1138 1055 1172 1083
rect 1274 1083 1308 1089
rect 1274 1055 1308 1083
rect 1410 1083 1444 1089
rect 1410 1055 1444 1083
rect 1546 1083 1580 1089
rect 1546 1055 1580 1083
rect 1682 1083 1716 1089
rect 1682 1055 1716 1083
rect 1818 1083 1852 1089
rect 1818 1055 1852 1083
rect 47 597 81 631
rect 229 257 263 261
rect 229 227 263 257
rect 311 301 345 335
rect 628 449 662 483
rect 556 375 590 409
rect 824 301 842 335
rect 842 301 858 335
rect 910 301 944 335
rect 1074 449 1108 483
rect 1273 449 1307 483
rect 1170 369 1204 403
rect 1838 597 1872 631
rect 1667 523 1701 557
rect 1687 369 1721 403
rect 1409 301 1443 335
rect 1545 257 1579 261
rect 1545 227 1579 257
rect 50 27 84 55
rect 50 21 84 27
rect 186 27 220 55
rect 186 21 220 27
rect 322 27 356 55
rect 322 21 356 27
rect 458 27 492 55
rect 458 21 492 27
rect 594 27 628 55
rect 594 21 628 27
rect 730 27 764 55
rect 730 21 764 27
rect 866 27 900 55
rect 866 21 900 27
rect 1002 27 1036 55
rect 1002 21 1036 27
rect 1138 27 1172 55
rect 1138 21 1172 27
rect 1274 27 1308 55
rect 1274 21 1308 27
rect 1410 27 1444 55
rect 1410 21 1444 27
rect 1546 27 1580 55
rect 1546 21 1580 27
rect 1682 27 1716 55
rect 1682 21 1716 27
rect 1818 27 1852 55
rect 1818 21 1852 27
<< metal1 >>
rect 0 1089 1914 1110
rect 0 1055 50 1089
rect 84 1055 186 1089
rect 220 1055 322 1089
rect 356 1055 458 1089
rect 492 1055 594 1089
rect 628 1055 730 1089
rect 764 1055 866 1089
rect 900 1055 1002 1089
rect 1036 1055 1138 1089
rect 1172 1055 1274 1089
rect 1308 1055 1410 1089
rect 1444 1055 1546 1089
rect 1580 1055 1682 1089
rect 1716 1055 1818 1089
rect 1852 1055 1914 1089
rect 0 1049 1914 1055
rect 35 631 93 637
rect 1826 631 1884 637
rect 35 597 47 631
rect 81 597 127 631
rect 1804 597 1838 631
rect 1872 597 1884 631
rect 35 591 93 597
rect 1826 591 1884 597
rect 1655 557 1713 563
rect 1632 523 1667 557
rect 1701 523 1713 557
rect 1655 517 1713 523
rect 616 483 674 489
rect 1062 483 1120 489
rect 1261 483 1319 489
rect 616 449 628 483
rect 662 449 1074 483
rect 1108 449 1273 483
rect 1307 449 1319 483
rect 616 443 674 449
rect 1062 443 1120 449
rect 1261 443 1319 449
rect 544 409 602 415
rect 544 375 556 409
rect 590 375 624 409
rect 1158 403 1216 409
rect 1675 403 1733 409
rect 544 369 602 375
rect 1158 369 1170 403
rect 1204 369 1687 403
rect 1721 369 1733 403
rect 1158 363 1216 369
rect 1675 363 1733 369
rect 299 335 357 341
rect 812 335 870 341
rect 299 301 311 335
rect 345 301 824 335
rect 858 301 870 335
rect 299 295 357 301
rect 812 295 870 301
rect 898 335 956 341
rect 1397 335 1455 341
rect 898 301 910 335
rect 944 301 1409 335
rect 1443 301 1455 335
rect 898 295 956 301
rect 1397 295 1455 301
rect 217 261 275 267
rect 1533 261 1591 267
rect 217 227 229 261
rect 263 227 1545 261
rect 1579 227 1591 261
rect 217 221 275 227
rect 1533 221 1591 227
rect 0 55 1914 61
rect 0 21 50 55
rect 84 21 186 55
rect 220 21 322 55
rect 356 21 458 55
rect 492 21 594 55
rect 628 21 730 55
rect 764 21 866 55
rect 900 21 1002 55
rect 1036 21 1138 55
rect 1172 21 1274 55
rect 1308 21 1410 55
rect 1444 21 1546 55
rect 1580 21 1682 55
rect 1716 21 1818 55
rect 1852 21 1914 55
rect 0 0 1914 21
<< labels >>
rlabel viali 65 614 65 614 1 RN
port 1 n
rlabel viali 573 392 573 392 1 D
port 2 n
rlabel viali 1290 466 1290 466 1 CK
port 3 n
rlabel viali 1855 614 1855 614 1 Q
port 4 n
rlabel viali 1685 540 1685 540 1 QN
port 5 n
rlabel viali 67 48 67 48 1 gnd
rlabel viali 67 1062 67 1062 1 vdd
<< end >>
