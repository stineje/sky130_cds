* File: sky130_osu_sc_15T_ls__ant.pex.spice
* Created: Fri Nov 12 14:54:17 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__ANT%GND 7 10 17 20
r16 17 20 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=0.19
+ $X2=0.495 $Y2=0.24
r17 10 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r18 7 10 0.369697 $w=9.88e-07 $l=3e-08 $layer=LI1_cond $X=0.495 $Y=0.22
+ $X2=0.495 $Y2=0.19
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ANT%VDD 1 9 11 18 23
r7 23 26 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=5.31
+ $X2=0.495 $Y2=5.36
r8 18 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r9 16 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r10 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r11 11 16 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.245
r12 11 13 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r13 9 13 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r14 1 21 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r15 1 18 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__ANT%A 1 5 15 19 22 27 30 33 37 41 46 49 51
r23 46 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.33
+ $X2=0.32 $Y2=2.33
r24 43 46 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.26 $Y=2.33 $X2=0.32
+ $Y2=2.33
r25 39 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.69 $Y=1.655
+ $X2=0.69 $Y2=0.865
r26 38 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.74
+ $X2=0.26 $Y2=1.74
r27 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.74
+ $X2=0.69 $Y2=1.655
r28 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.74
+ $X2=0.345 $Y2=1.74
r29 33 35 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r30 31 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.415
+ $X2=0.26 $Y2=2.33
r31 31 33 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.26 $Y=2.415
+ $X2=0.26 $Y2=3.205
r32 30 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.245
+ $X2=0.26 $Y2=2.33
r33 29 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.825
+ $X2=0.26 $Y2=1.74
r34 29 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.26 $Y=1.825
+ $X2=0.26 $Y2=2.245
r35 25 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.655
+ $X2=0.26 $Y2=1.74
r36 25 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.26 $Y=1.655
+ $X2=0.26 $Y2=0.865
r37 22 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.33 $X2=0.32 $Y2=2.33
r38 22 24 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=2.33
+ $X2=0.362 $Y2=2.495
r39 22 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=2.33
+ $X2=0.362 $Y2=2.165
r40 19 24 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.495
r41 15 23 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=2.165
r42 5 35 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r43 5 33 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r44 1 41 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
r45 1 27 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

