* File: sky130_osu_sc_18T_hs__dlat_1.pex.spice
* Created: Fri Nov 12 13:49:50 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%GND 1 2 3 4 59 63 65 75 77 84 86 93 112
+ 114
r113 112 114 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r114 91 93 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.365 $Y=0.305
+ $X2=4.365 $Y2=0.825
r115 82 84 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.985 $Y=0.305
+ $X2=2.985 $Y2=0.825
r116 78 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.152
+ $X2=2.035 $Y2=0.152
r117 73 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.035 $Y=0.305
+ $X2=2.035 $Y2=0.152
r118 73 75 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.035 $Y=0.305
+ $X2=2.035 $Y2=0.825
r119 65 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.152
+ $X2=2.035 $Y2=0.152
r120 61 63 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.285 $Y=0.305
+ $X2=0.285 $Y2=0.825
r121 59 114 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r122 59 112 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r123 59 91 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.365 $Y2=0.305
r124 59 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.28 $Y2=0.152
r125 59 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.985 $Y=0.152
+ $X2=2.985 $Y2=0.305
r126 59 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.152
+ $X2=2.9 $Y2=0.152
r127 59 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.152
+ $X2=3.07 $Y2=0.152
r128 59 61 4.36583 $w=1.7e-07 $l=1.96746e-07 $layer=LI1_cond $X=0.185 $Y=0.152
+ $X2=0.285 $Y2=0.305
r129 59 66 3.19241 $w=3.05e-07 $l=1.85e-07 $layer=LI1_cond $X=0.185 $Y=0.152
+ $X2=0.37 $Y2=0.152
r130 59 86 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.28 $Y2=0.152
r131 59 87 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.07 $Y2=0.152
r132 59 77 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.9 $Y2=0.152
r133 59 78 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.12 $Y2=0.152
r134 59 65 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.95 $Y2=0.152
r135 59 66 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.37 $Y2=0.152
r136 4 93 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.225
+ $Y=0.575 $X2=4.365 $Y2=0.825
r137 3 84 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=2.86
+ $Y=0.575 $X2=2.985 $Y2=0.825
r138 2 75 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.895
+ $Y=0.575 $X2=2.035 $Y2=0.825
r139 1 63 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%VDD 1 2 3 4 45 49 53 61 65 71 75 81 94
+ 97 101
c61 81 0 1.98165e-19 $X=4.365 $Y=3.455
r62 97 101 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=4.42 $Y2=6.507
r63 94 101 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=6.47
+ $X2=4.42 $Y2=6.47
r64 88 97 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r65 81 84 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.365 $Y=3.455
+ $X2=4.365 $Y2=5.835
r66 79 94 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.365 $Y=6.355
+ $X2=4.365 $Y2=6.507
r67 79 84 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.365 $Y=6.355
+ $X2=4.365 $Y2=5.835
r68 76 92 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=6.507
+ $X2=2.985 $Y2=6.507
r69 76 78 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=3.07 $Y=6.507
+ $X2=3.74 $Y2=6.507
r70 75 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=6.507
+ $X2=4.365 $Y2=6.507
r71 75 78 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=4.28 $Y=6.507
+ $X2=3.74 $Y2=6.507
r72 71 74 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.985 $Y=3.795
+ $X2=2.985 $Y2=5.835
r73 69 92 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.985 $Y=6.355
+ $X2=2.985 $Y2=6.507
r74 69 74 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.985 $Y=6.355
+ $X2=2.985 $Y2=5.835
r75 66 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=6.507
+ $X2=2.035 $Y2=6.507
r76 66 68 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=2.12 $Y=6.507
+ $X2=2.38 $Y2=6.507
r77 65 92 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=6.507
+ $X2=2.985 $Y2=6.507
r78 65 68 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=2.9 $Y=6.507
+ $X2=2.38 $Y2=6.507
r79 61 64 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.035 $Y=3.455
+ $X2=2.035 $Y2=5.835
r80 59 90 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.035 $Y=6.355
+ $X2=2.035 $Y2=6.507
r81 59 64 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.035 $Y=6.355
+ $X2=2.035 $Y2=5.835
r82 56 58 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r83 54 88 3.19971 $w=3.05e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=6.507
+ $X2=0.185 $Y2=6.507
r84 54 56 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=0.37 $Y=6.507
+ $X2=1.02 $Y2=6.507
r85 53 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=6.507
+ $X2=2.035 $Y2=6.507
r86 53 58 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.95 $Y=6.507
+ $X2=1.7 $Y2=6.507
r87 49 52 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.285 $Y=3.795
+ $X2=0.285 $Y2=5.835
r88 47 88 4.35853 $w=1.7e-07 $l=1.95714e-07 $layer=LI1_cond $X=0.285 $Y=6.355
+ $X2=0.185 $Y2=6.507
r89 47 52 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.285 $Y=6.355
+ $X2=0.285 $Y2=5.835
r90 45 94 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r91 45 78 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r92 45 92 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r93 45 68 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r94 45 58 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r95 45 56 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r96 45 88 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r97 4 84 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.225
+ $Y=3.085 $X2=4.365 $Y2=5.835
r98 4 81 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.225
+ $Y=3.085 $X2=4.365 $Y2=3.455
r99 3 74 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=2.86
+ $Y=3.085 $X2=2.985 $Y2=5.835
r100 3 71 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=2.86
+ $Y=3.085 $X2=2.985 $Y2=3.795
r101 2 64 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.895
+ $Y=3.085 $X2=2.035 $Y2=5.835
r102 2 61 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.895
+ $Y=3.085 $X2=2.035 $Y2=3.455
r103 1 52 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.16
+ $Y=3.085 $X2=0.285 $Y2=5.835
r104 1 49 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=0.16
+ $Y=3.085 $X2=0.285 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%D 1 3 9 12 15 19 21 23 26 29 33 38 40 41
+ 42 43 44 47 51 56 61 65 66 71 75
c119 40 0 1.57671e-19 $X=0.58 $Y=3.1
c120 19 0 1.65121e-19 $X=0.5 $Y=4.585
r121 66 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.725 $Y=1.85
+ $X2=0.58 $Y2=1.85
r122 65 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.85 $Y=1.85
+ $X2=2.995 $Y2=1.85
r123 65 66 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=2.85 $Y=1.85
+ $X2=0.725 $Y2=1.85
r124 61 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.44 $Y=2.22
+ $X2=0.44 $Y2=2.22
r125 61 64 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.51 $Y=2.22
+ $X2=0.51 $Y2=2.385
r126 61 62 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.51 $Y=2.22
+ $X2=0.51 $Y2=2.055
r127 56 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.995 $Y=1.85
+ $X2=2.995 $Y2=1.85
r128 51 53 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.16 $Y=3.455
+ $X2=1.16 $Y2=5.835
r129 49 51 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=1.16 $Y=3.27
+ $X2=1.16 $Y2=3.455
r130 45 47 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=1.16 $Y=1.345
+ $X2=1.16 $Y2=0.825
r131 43 49 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.99 $Y=3.185
+ $X2=1.16 $Y2=3.27
r132 43 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.99 $Y=3.185
+ $X2=0.665 $Y2=3.185
r133 41 45 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.99 $Y=1.43
+ $X2=1.16 $Y2=1.345
r134 41 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.99 $Y=1.43
+ $X2=0.665 $Y2=1.43
r135 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.58 $Y=3.1
+ $X2=0.665 $Y2=3.185
r136 40 64 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.58 $Y=3.1
+ $X2=0.58 $Y2=2.385
r137 38 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.58 $Y=1.85
+ $X2=0.58 $Y2=1.85
r138 38 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.58 $Y=1.85
+ $X2=0.58 $Y2=2.055
r139 35 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.58 $Y=1.515
+ $X2=0.665 $Y2=1.43
r140 35 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.58 $Y=1.515
+ $X2=0.58 $Y2=1.85
r141 31 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=1.85 $X2=2.995 $Y2=1.85
r142 31 33 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.995 $Y=1.85
+ $X2=3.2 $Y2=1.85
r143 24 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=2.015
+ $X2=3.2 $Y2=1.85
r144 24 26 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=3.2 $Y=2.015
+ $X2=3.2 $Y2=4.585
r145 21 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.685
+ $X2=3.2 $Y2=1.85
r146 21 23 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.2 $Y=1.685
+ $X2=3.2 $Y2=1.075
r147 19 29 1112.7 $w=1.5e-07 $l=2.17e-06 $layer=POLY_cond $X=0.5 $Y=4.585
+ $X2=0.5 $Y2=2.415
r148 15 28 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.5 $Y=1.075
+ $X2=0.5 $Y2=2.005
r149 12 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.44
+ $Y=2.22 $X2=0.44 $Y2=2.22
r150 10 29 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.44 $Y=2.28
+ $X2=0.44 $Y2=2.415
r151 10 12 13.3304 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=0.44 $Y=2.28 $X2=0.44
+ $Y2=2.22
r152 9 28 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.44 $Y=2.14
+ $X2=0.44 $Y2=2.005
r153 9 12 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=0.44 $Y=2.14 $X2=0.44
+ $Y2=2.22
r154 3 53 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=0.935
+ $Y=3.085 $X2=1.16 $Y2=5.835
r155 3 51 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=0.935
+ $Y=3.085 $X2=1.16 $Y2=3.455
r156 1 47 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=0.575 $X2=1.16 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%CK 3 6 10 11 13 16 18 19 22 25 26 31 33
+ 34 36 43 47 48 53
c133 34 0 1.65121e-19 $X=1.005 $Y=2.59
r134 48 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.545 $Y=2.59
+ $X2=1.4 $Y2=2.59
r135 47 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.25 $Y=2.59
+ $X2=2.395 $Y2=2.59
r136 47 48 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=2.25 $Y=2.59
+ $X2=1.545 $Y2=2.59
r137 43 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.4 $Y=2.59 $X2=1.4
+ $Y2=2.59
r138 43 45 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.4 $Y=2.59
+ $X2=1.4 $Y2=2.765
r139 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.395 $Y=2.59
+ $X2=2.395 $Y2=2.59
r140 36 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.395 $Y=2.59
+ $X2=2.395 $Y2=2.765
r141 33 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.59
+ $X2=1.4 $Y2=2.59
r142 33 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.315 $Y=2.59
+ $X2=1.005 $Y2=2.59
r143 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.92 $Y=2.505
+ $X2=1.005 $Y2=2.59
r144 29 31 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.92 $Y=2.505
+ $X2=0.92 $Y2=1.85
r145 28 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=2.765 $X2=2.395 $Y2=2.765
r146 25 26 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.277 $Y=1.685
+ $X2=2.277 $Y2=1.835
r147 22 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=2.765 $X2=1.4 $Y2=2.765
r148 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=2.765
+ $X2=1.4 $Y2=2.93
r149 18 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.92
+ $Y=1.85 $X2=0.92 $Y2=1.85
r150 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.85
+ $X2=0.92 $Y2=1.685
r151 16 28 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=2.305 $Y=2.6
+ $X2=2.352 $Y2=2.765
r152 16 26 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.305 $Y=2.6
+ $X2=2.305 $Y2=1.835
r153 11 28 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=2.25 $Y=2.93
+ $X2=2.352 $Y2=2.765
r154 11 13 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.25 $Y=2.93
+ $X2=2.25 $Y2=4.585
r155 10 25 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.25 $Y=1.075
+ $X2=2.25 $Y2=1.685
r156 6 24 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.46 $Y=4.585
+ $X2=1.46 $Y2=2.93
r157 3 19 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.86 $Y=1.075
+ $X2=0.86 $Y2=1.685
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%A_157_445# 1 3 11 13 14 16 19 21 22 24
+ 30 33 36 41 42 45 49
r119 47 49 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.465 $Y=3.185
+ $X2=2.735 $Y2=3.185
r120 43 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.465 $Y=2.19
+ $X2=2.735 $Y2=2.19
r121 41 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=3.1
+ $X2=2.735 $Y2=3.185
r122 40 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=2.19
r123 40 41 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=3.1
r124 36 38 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.465 $Y=3.455
+ $X2=2.465 $Y2=5.835
r125 34 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.27
+ $X2=2.465 $Y2=3.185
r126 34 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.465 $Y=3.27
+ $X2=2.465 $Y2=3.455
r127 33 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=2.105
+ $X2=2.465 $Y2=2.19
r128 32 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.935
+ $X2=2.465 $Y2=1.85
r129 32 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.465 $Y=1.935
+ $X2=2.465 $Y2=2.105
r130 28 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.765
+ $X2=2.465 $Y2=1.85
r131 28 30 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.465 $Y=1.765
+ $X2=2.465 $Y2=0.825
r132 24 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=1.85
+ $X2=2.465 $Y2=1.85
r133 24 26 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.38 $Y=1.85
+ $X2=1.4 $Y2=1.85
r134 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=1.85 $X2=1.4 $Y2=1.85
r135 21 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.85
+ $X2=1.4 $Y2=2.015
r136 21 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.85
+ $X2=1.4 $Y2=1.685
r137 19 22 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.46 $Y=1.075
+ $X2=1.46 $Y2=1.685
r138 16 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.34 $Y=2.225
+ $X2=1.34 $Y2=2.015
r139 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.265 $Y=2.3
+ $X2=1.34 $Y2=2.225
r140 13 14 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.265 $Y=2.3
+ $X2=0.935 $Y2=2.3
r141 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.86 $Y=2.375
+ $X2=0.935 $Y2=2.3
r142 9 11 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=0.86 $Y=2.375
+ $X2=0.86 $Y2=4.585
r143 3 38 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.325
+ $Y=3.085 $X2=2.465 $Y2=5.835
r144 3 36 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.325
+ $Y=3.085 $X2=2.465 $Y2=3.455
r145 1 30 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%A_349_89# 1 3 11 15 23 26 28 32 33 35 36
+ 37 38 40 46 50 56 59 60 61 66
c131 37 0 8.77106e-20 $X=4.125 $Y=2.855
c132 32 0 2.20654e-19 $X=4.035 $Y=2.19
r133 61 63 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.025 $Y=2.19
+ $X2=1.88 $Y2=2.19
r134 60 66 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.89 $Y=2.19
+ $X2=4.035 $Y2=2.19
r135 60 61 1.79578 $w=1.7e-07 $l=1.865e-06 $layer=MET1_cond $X=3.89 $Y=2.19
+ $X2=2.025 $Y2=2.19
r136 56 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.035 $Y=2.19
+ $X2=4.035 $Y2=2.19
r137 54 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.19
+ $X2=3.415 $Y2=2.19
r138 54 56 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.5 $Y=2.19
+ $X2=4.035 $Y2=2.19
r139 50 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.415 $Y=3.455
+ $X2=3.415 $Y2=5.835
r140 48 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=2.275
+ $X2=3.415 $Y2=2.19
r141 48 50 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.415 $Y=2.275
+ $X2=3.415 $Y2=3.455
r142 44 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=2.105
+ $X2=3.415 $Y2=2.19
r143 44 46 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=3.415 $Y=2.105
+ $X2=3.415 $Y2=0.825
r144 40 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.88 $Y=2.19
+ $X2=1.88 $Y2=2.19
r145 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=2.855
+ $X2=4.125 $Y2=3.005
r146 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=1.65
+ $X2=4.125 $Y2=1.8
r147 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=4.1 $Y=2.355 $X2=4.1
+ $Y2=2.855
r148 33 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.1 $Y=2.025
+ $X2=4.1 $Y2=1.8
r149 32 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=2.19 $X2=4.035 $Y2=2.19
r150 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.037 $Y=2.19
+ $X2=4.037 $Y2=2.355
r151 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.037 $Y=2.19
+ $X2=4.037 $Y2=2.025
r152 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=2.19 $X2=1.88 $Y2=2.19
r153 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=2.19
+ $X2=1.88 $Y2=2.355
r154 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=2.19
+ $X2=1.88 $Y2=2.025
r155 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=4.15 $Y=4.585
+ $X2=4.15 $Y2=3.005
r156 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.15 $Y=1.075
+ $X2=4.15 $Y2=1.65
r157 15 30 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=1.82 $Y=4.585
+ $X2=1.82 $Y2=2.355
r158 11 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.82 $Y=1.075
+ $X2=1.82 $Y2=2.025
r159 3 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.275
+ $Y=3.085 $X2=3.415 $Y2=5.835
r160 3 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.275
+ $Y=3.085 $X2=3.415 $Y2=3.455
r161 1 46 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.275
+ $Y=0.575 $X2=3.415 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c74 44 0 8.77106e-20 $X=3.94 $Y=2.96
c75 35 0 9.99996e-20 $X=4.435 $Y=2.765
c76 33 0 1.20654e-19 $X=4.435 $Y=1.85
c77 18 0 1.98165e-19 $X=4.52 $Y=2.395
r78 42 44 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=3.935 $Y=2.96
+ $X2=3.94 $Y2=2.96
r79 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.52 $Y=2.68
+ $X2=4.52 $Y2=2.395
r80 37 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.52 $Y=1.935
+ $X2=4.52 $Y2=2.395
r81 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=2.765
+ $X2=4.52 $Y2=2.68
r82 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=2.765
+ $X2=4.02 $Y2=2.765
r83 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=1.85
+ $X2=4.52 $Y2=1.935
r84 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=1.85
+ $X2=4.02 $Y2=1.85
r85 29 31 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.935 $Y=3.455
+ $X2=3.935 $Y2=5.835
r86 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=2.96
+ $X2=3.935 $Y2=2.96
r87 27 29 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.935 $Y=2.96
+ $X2=3.935 $Y2=3.455
r88 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=2.85
+ $X2=4.02 $Y2=2.765
r89 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.935 $Y=2.85
+ $X2=3.935 $Y2=2.96
r90 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=1.765
+ $X2=4.02 $Y2=1.85
r91 21 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.935 $Y=1.765
+ $X2=3.935 $Y2=0.825
r92 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=2.395 $X2=4.52 $Y2=2.395
r93 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.395
+ $X2=4.52 $Y2=2.56
r94 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.395
+ $X2=4.52 $Y2=2.23
r95 15 20 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=4.58 $Y=4.585
+ $X2=4.58 $Y2=2.56
r96 11 19 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=4.58 $Y=1.075
+ $X2=4.58 $Y2=2.23
r97 3 31 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=3.81
+ $Y=3.085 $X2=3.935 $Y2=5.835
r98 3 29 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=3.81
+ $Y=3.085 $X2=3.935 $Y2=3.455
r99 1 23 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=3.81
+ $Y=0.575 $X2=3.935 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DLAT_1%Q 1 3 11 15 17 24 25 28
r19 24 25 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=4.86 $Y=1.61
+ $X2=4.86 $Y2=3.16
r20 23 24 8.82722 $w=2.33e-07 $l=1.8e-07 $layer=LI1_cond $X=4.827 $Y=1.43
+ $X2=4.827 $Y2=1.61
r21 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.795 $Y=3.455
+ $X2=4.795 $Y2=5.835
r22 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.795 $Y=3.33
+ $X2=4.795 $Y2=3.33
r23 15 25 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.827 $Y=3.33
+ $X2=4.827 $Y2=3.16
r24 15 17 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.795 $Y=3.33
+ $X2=4.795 $Y2=3.455
r25 11 23 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.795 $Y=0.825
+ $X2=4.795 $Y2=1.43
r26 3 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.655
+ $Y=3.085 $X2=4.795 $Y2=5.835
r27 3 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.655
+ $Y=3.085 $X2=4.795 $Y2=3.455
r28 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.655
+ $Y=0.575 $X2=4.795 $Y2=0.825
.ends

