* File: sky130_osu_sc_18T_ms__buf_l.pxi.spice
* Created: Thu Oct 29 17:28:39 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__BUF_L%GND N_GND_M1001_d N_GND_M1001_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_MS__BUF_L%GND
x_PM_SKY130_OSU_SC_18T_MS__BUF_L%VDD N_VDD_M1003_d N_VDD_M1003_b N_VDD_c_27_p
+ N_VDD_c_28_p VDD N_VDD_c_29_p N_VDD_c_35_p PM_SKY130_OSU_SC_18T_MS__BUF_L%VDD
x_PM_SKY130_OSU_SC_18T_MS__BUF_L%A N_A_M1001_g N_A_M1003_g A N_A_c_49_n
+ N_A_c_50_n PM_SKY130_OSU_SC_18T_MS__BUF_L%A
x_PM_SKY130_OSU_SC_18T_MS__BUF_L%A_27_115# N_A_27_115#_M1001_s
+ N_A_27_115#_M1003_s N_A_27_115#_M1000_g N_A_27_115#_M1002_g N_A_27_115#_c_83_n
+ N_A_27_115#_c_84_n N_A_27_115#_c_85_n N_A_27_115#_c_88_n N_A_27_115#_c_89_n
+ N_A_27_115#_c_90_n N_A_27_115#_c_91_n N_A_27_115#_c_92_n
+ PM_SKY130_OSU_SC_18T_MS__BUF_L%A_27_115#
x_PM_SKY130_OSU_SC_18T_MS__BUF_L%Y N_Y_M1000_d N_Y_M1002_d Y N_Y_c_134_n
+ N_Y_c_135_n N_Y_c_139_n N_Y_c_136_n PM_SKY130_OSU_SC_18T_MS__BUF_L%Y
cc_1 N_GND_M1001_b N_A_M1001_g 0.0735339f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1001_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_A_M1001_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=0.945
cc_4 N_GND_c_4_p N_A_M1001_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=0.945
cc_5 N_GND_M1001_b N_A_M1003_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=5.085
cc_6 N_GND_M1001_b N_A_c_49_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_7 N_GND_M1001_b N_A_c_50_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_8 N_GND_M1001_b N_A_27_115#_M1000_g 0.0510561f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.945
cc_9 N_GND_c_3_p N_A_27_115#_M1000_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=0.945
cc_10 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.905
+ $Y2=0.945
cc_11 N_GND_M1001_b N_A_27_115#_c_83_n 0.0597491f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.86
cc_12 N_GND_M1001_b N_A_27_115#_c_84_n 0.0168393f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.935
cc_13 N_GND_M1001_b N_A_27_115#_c_85_n 0.0271353f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_14 N_GND_c_2_p N_A_27_115#_c_85_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_15 N_GND_c_4_p N_A_27_115#_c_85_n 0.00476261f $X=1.02 $Y=0.17 $X2=0.26
+ $Y2=0.825
cc_16 N_GND_M1001_b N_A_27_115#_c_88_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=4.475
cc_17 N_GND_M1001_b N_A_27_115#_c_89_n 0.0172272f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.935
cc_18 N_GND_M1001_b N_A_27_115#_c_90_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.935
cc_19 N_GND_M1001_b N_A_27_115#_c_91_n 0.00663593f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.935
cc_20 N_GND_M1001_b N_A_27_115#_c_92_n 0.0562401f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=1.935
cc_21 N_GND_M1001_b Y 0.0164841f $X=-0.045 $Y=0 $X2=1.07 $Y2=2.26
cc_22 N_GND_M1001_b N_Y_c_134_n 0.014537f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.48
cc_23 N_GND_M1001_b N_Y_c_135_n 0.00501078f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.96
cc_24 N_GND_M1001_b N_Y_c_136_n 0.0198198f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.825
cc_25 N_GND_c_4_p N_Y_c_136_n 0.00476261f $X=1.02 $Y=0.17 $X2=1.12 $Y2=0.825
cc_26 N_VDD_M1003_b N_A_M1003_g 0.0817671f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_27 N_VDD_c_27_p N_A_M1003_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475 $Y2=5.085
cc_28 N_VDD_c_28_p N_A_M1003_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.475 $Y2=5.085
cc_29 N_VDD_c_29_p N_A_M1003_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=5.085
cc_30 N_VDD_M1003_b A 0.0157561f $X=-0.045 $Y=2.905 $X2=0.635 $Y2=3.33
cc_31 N_VDD_M1003_b N_A_c_49_n 0.011209f $X=-0.045 $Y=2.905 $X2=0.635 $Y2=2.48
cc_32 N_VDD_M1003_b N_A_27_115#_M1002_g 0.0756766f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=5.085
cc_33 N_VDD_c_28_p N_A_27_115#_M1002_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.905
+ $Y2=5.085
cc_34 N_VDD_c_29_p N_A_27_115#_M1002_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.905
+ $Y2=5.085
cc_35 N_VDD_c_35_p N_A_27_115#_M1002_g 0.00606474f $X=1.02 $Y=6.44 $X2=0.905
+ $Y2=5.085
cc_36 N_VDD_M1003_b N_A_27_115#_c_84_n 0.0187682f $X=-0.045 $Y=2.905 $X2=1.18
+ $Y2=2.935
cc_37 N_VDD_M1003_b N_A_27_115#_c_88_n 0.0580517f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.475
cc_38 N_VDD_c_27_p N_A_27_115#_c_88_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=4.475
cc_39 N_VDD_c_29_p N_A_27_115#_c_88_n 0.00476261f $X=1.02 $Y=6.49 $X2=0.26
+ $Y2=4.475
cc_40 N_VDD_M1003_b N_Y_c_135_n 0.0107503f $X=-0.045 $Y=2.905 $X2=1.12 $Y2=2.96
cc_41 N_VDD_M1003_b N_Y_c_139_n 0.051089f $X=-0.045 $Y=2.905 $X2=1.12 $Y2=2.96
cc_42 N_VDD_c_29_p N_Y_c_139_n 0.00476261f $X=1.02 $Y=6.49 $X2=1.12 $Y2=2.96
cc_43 N_VDD_c_35_p N_Y_c_139_n 0.00736239f $X=1.02 $Y=6.44 $X2=1.12 $Y2=2.96
cc_44 N_A_M1001_g N_A_27_115#_M1000_g 0.0527922f $X=0.475 $Y=0.945 $X2=0.905
+ $Y2=0.945
cc_45 A N_A_27_115#_M1002_g 0.00419145f $X=0.635 $Y=3.33 $X2=0.905 $Y2=5.085
cc_46 N_A_M1001_g N_A_27_115#_c_83_n 0.00260138f $X=0.475 $Y=0.945 $X2=1.18
+ $Y2=2.86
cc_47 N_A_M1003_g N_A_27_115#_c_83_n 0.00209773f $X=0.475 $Y=5.085 $X2=1.18
+ $Y2=2.86
cc_48 N_A_c_49_n N_A_27_115#_c_83_n 0.00361737f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_49 N_A_c_50_n N_A_27_115#_c_83_n 0.0139096f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.86
cc_50 N_A_M1003_g N_A_27_115#_c_84_n 0.0639305f $X=0.475 $Y=5.085 $X2=1.18
+ $Y2=2.935
cc_51 N_A_c_49_n N_A_27_115#_c_84_n 0.00468272f $X=0.635 $Y=2.48 $X2=1.18
+ $Y2=2.935
cc_52 N_A_M1001_g N_A_27_115#_c_85_n 0.0264643f $X=0.475 $Y=0.945 $X2=0.26
+ $Y2=0.825
cc_53 N_A_M1001_g N_A_27_115#_c_88_n 0.0668001f $X=0.475 $Y=0.945 $X2=0.26
+ $Y2=4.475
cc_54 A N_A_27_115#_c_88_n 0.0155137f $X=0.635 $Y=3.33 $X2=0.26 $Y2=4.475
cc_55 N_A_c_49_n N_A_27_115#_c_88_n 0.0696932f $X=0.635 $Y=2.48 $X2=0.26
+ $Y2=4.475
cc_56 N_A_M1001_g N_A_27_115#_c_89_n 0.0207696f $X=0.475 $Y=0.945 $X2=0.88
+ $Y2=1.935
cc_57 N_A_c_49_n N_A_27_115#_c_89_n 0.00886797f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_58 N_A_c_50_n N_A_27_115#_c_89_n 0.00273049f $X=0.635 $Y=2.48 $X2=0.88
+ $Y2=1.935
cc_59 N_A_M1001_g N_A_27_115#_c_91_n 6.59135e-19 $X=0.475 $Y=0.945 $X2=0.965
+ $Y2=1.935
cc_60 N_A_M1001_g Y 0.00310306f $X=0.475 $Y=0.945 $X2=1.07 $Y2=2.26
cc_61 N_A_c_49_n Y 0.0200396f $X=0.635 $Y=2.48 $X2=1.07 $Y2=2.26
cc_62 N_A_c_50_n Y 0.00441844f $X=0.635 $Y=2.48 $X2=1.07 $Y2=2.26
cc_63 N_A_M1001_g N_Y_c_134_n 0.00102215f $X=0.475 $Y=0.945 $X2=1.12 $Y2=1.48
cc_64 N_A_c_49_n N_Y_c_135_n 0.00609526f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_65 A N_Y_c_139_n 0.00731851f $X=0.635 $Y=3.33 $X2=1.12 $Y2=2.96
cc_66 N_A_c_49_n N_Y_c_139_n 0.0203054f $X=0.635 $Y=2.48 $X2=1.12 $Y2=2.96
cc_67 N_A_27_115#_M1000_g Y 0.00406656f $X=0.905 $Y=0.945 $X2=1.07 $Y2=2.26
cc_68 N_A_27_115#_c_83_n Y 0.0310322f $X=1.18 $Y=2.86 $X2=1.07 $Y2=2.26
cc_69 N_A_27_115#_c_89_n Y 8.73078e-19 $X=0.88 $Y=1.935 $X2=1.07 $Y2=2.26
cc_70 N_A_27_115#_c_91_n Y 0.0121742f $X=0.965 $Y=1.935 $X2=1.07 $Y2=2.26
cc_71 N_A_27_115#_c_92_n Y 0.0161039f $X=1.18 $Y=1.935 $X2=1.07 $Y2=2.26
cc_72 N_A_27_115#_M1000_g N_Y_c_134_n 0.00714414f $X=0.905 $Y=0.945 $X2=1.12
+ $Y2=1.48
cc_73 N_A_27_115#_c_91_n N_Y_c_134_n 0.00278861f $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=1.48
cc_74 N_A_27_115#_c_92_n N_Y_c_134_n 0.0014753f $X=1.18 $Y=1.935 $X2=1.12
+ $Y2=1.48
cc_75 N_A_27_115#_M1002_g N_Y_c_135_n 0.0015856f $X=0.905 $Y=5.085 $X2=1.12
+ $Y2=2.96
cc_76 N_A_27_115#_c_83_n N_Y_c_135_n 0.00226191f $X=1.18 $Y=2.86 $X2=1.12
+ $Y2=2.96
cc_77 N_A_27_115#_c_84_n N_Y_c_135_n 0.00513726f $X=1.18 $Y=2.935 $X2=1.12
+ $Y2=2.96
cc_78 N_A_27_115#_M1002_g N_Y_c_139_n 0.0402429f $X=0.905 $Y=5.085 $X2=1.12
+ $Y2=2.96
cc_79 N_A_27_115#_c_84_n N_Y_c_139_n 0.0134943f $X=1.18 $Y=2.935 $X2=1.12
+ $Y2=2.96
cc_80 N_A_27_115#_M1000_g N_Y_c_136_n 0.0152627f $X=0.905 $Y=0.945 $X2=1.12
+ $Y2=0.825
cc_81 N_A_27_115#_c_91_n N_Y_c_136_n 7.50437e-19 $X=0.965 $Y=1.935 $X2=1.12
+ $Y2=0.825
cc_82 N_A_27_115#_c_92_n N_Y_c_136_n 0.00477112f $X=1.18 $Y=1.935 $X2=1.12
+ $Y2=0.825
