* File: sky130_osu_sc_12T_ls__and2_l.pex.spice
* Created: Fri Nov 12 15:34:19 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__AND2_L%GND 1 17 19 26 35 38
r34 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r35 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r36 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r37 17 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r38 17 19 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r39 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r40 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AND2_L%VDD 1 2 17 21 23 30 36 38 41
r28 38 41 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r29 28 36 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r30 28 30 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.275
r31 26 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r32 24 35 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r33 24 26 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r34 23 36 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r35 23 26 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r36 19 35 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r37 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.275
r38 17 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r39 17 35 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r40 2 30 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=3.025 $X2=1.12 $Y2=3.275
r41 1 21 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.275
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AND2_L%A 3 7 12 15 23
c33 15 0 1.6558e-19 $X=0.27 $Y=2.48
r34 21 23 0.001703 $w=3.67e-07 $l=5e-09 $layer=MET1_cond $X=0.322 $Y=2.48
+ $X2=0.322 $Y2=2.485
r35 15 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.48
r36 15 18 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.66
r37 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.66 $X2=0.27 $Y2=2.66
r38 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.66
+ $X2=0.475 $Y2=2.66
r39 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.825
+ $X2=0.475 $Y2=2.66
r40 5 7 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.475 $Y=2.825
+ $X2=0.475 $Y2=3.445
r41 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.495
+ $X2=0.475 $Y2=2.66
r42 1 3 892.213 $w=1.5e-07 $l=1.74e-06 $layer=POLY_cond $X=0.475 $Y=2.495
+ $X2=0.475 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AND2_L%B 3 7 10 14 20
c41 10 0 1.06013e-19 $X=0.95 $Y=2.31
c42 7 0 3.10762e-20 $X=0.905 $Y=3.445
r43 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.48
+ $X2=0.95 $Y2=2.48
r44 14 17 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.95 $Y=2.31
+ $X2=0.95 $Y2=2.48
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.31 $X2=0.95 $Y2=2.31
r46 10 12 47.0643 $w=3.25e-07 $l=1.7e-07 $layer=POLY_cond $X=0.922 $Y=2.31
+ $X2=0.922 $Y2=2.48
r47 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.31
+ $X2=0.922 $Y2=2.145
r48 7 12 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=0.905 $Y=3.445
+ $X2=0.905 $Y2=2.48
r49 3 11 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=0.835 $Y=0.755
+ $X2=0.835 $Y2=2.145
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AND2_L%A_27_115# 1 3 11 15 17 19 20 25 27 28 33
+ 37 39 40 41
c71 27 0 1.6558e-19 $X=0.525 $Y=1.755
r72 40 41 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.025
+ $X2=0.65 $Y2=3.195
r73 35 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.755
+ $X2=0.61 $Y2=1.755
r74 35 37 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.755
+ $X2=1.43 $Y2=1.755
r75 33 41 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.275 $X2=0.69
+ $Y2=3.195
r76 29 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.84 $X2=0.61
+ $Y2=1.755
r77 29 40 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=0.61 $Y=1.84
+ $X2=0.61 $Y2=3.025
r78 27 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.755
+ $X2=0.61 $Y2=1.755
r79 27 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.755
+ $X2=0.345 $Y2=1.755
r80 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.67
+ $X2=0.345 $Y2=1.755
r81 23 25 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.26 $Y=1.67
+ $X2=0.26 $Y2=0.74
r82 22 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.755 $X2=1.43 $Y2=1.755
r83 19 20 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.7
+ $X2=1.352 $Y2=2.85
r84 17 22 50.6121 $w=2.83e-07 $l=2.55137e-07 $layer=POLY_cond $X=1.37 $Y=1.99
+ $X2=1.412 $Y2=1.755
r85 17 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.99
+ $X2=1.37 $Y2=2.7
r86 15 20 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.335 $Y=3.445
+ $X2=1.335 $Y2=2.85
r87 9 22 38.6899 $w=2.83e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.59
+ $X2=1.412 $Y2=1.755
r88 9 11 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=1.335 $Y=1.59
+ $X2=1.335 $Y2=0.755
r89 3 33 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.025 $X2=0.69 $Y2=3.275
r90 1 25 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__AND2_L%Y 1 3 10 16 24 27 30
c33 30 0 1.37089e-19 $X=1.55 $Y=2.48
r34 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.48
r35 22 24 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.11
r36 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.485
+ $X2=1.55 $Y2=1.37
r37 21 24 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.485
+ $X2=1.55 $Y2=2.11
r38 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.48
r39 16 19 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=3.275
r40 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.37
+ $X2=1.55 $Y2=1.37
r41 10 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.37
r42 3 19 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=3.025 $X2=1.55 $Y2=3.275
r43 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

