magic
tech sky130A
magscale 1 2
timestamp 1612373379
<< nwell >>
rect -9 529 287 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 166 243
rect 110 131 121 215
rect 155 131 166 215
rect 110 115 166 131
rect 196 215 249 243
rect 196 131 207 215
rect 241 131 249 215
rect 196 115 249 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 949 166 965
rect 110 605 121 949
rect 155 605 166 949
rect 110 565 166 605
rect 196 949 249 965
rect 196 605 207 949
rect 241 605 249 949
rect 196 565 249 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 207 131 241 215
<< pdiffc >>
rect 35 741 69 949
rect 121 605 155 949
rect 207 605 241 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 992
rect 80 540 110 565
rect 166 540 196 565
rect 80 510 196 540
rect 80 442 110 510
rect 80 426 134 442
rect 80 392 90 426
rect 124 392 134 426
rect 80 376 134 392
rect 80 318 110 376
rect 80 268 196 318
rect 80 243 110 268
rect 166 243 196 268
rect 80 89 110 115
rect 166 89 196 115
<< polycont >>
rect 90 392 124 426
<< locali >>
rect 0 1089 286 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 286 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 121 949 155 965
rect 47 426 81 597
rect 121 557 155 605
rect 207 949 241 1049
rect 207 589 241 605
rect 47 392 90 426
rect 124 392 140 426
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 227
rect 121 115 155 131
rect 207 215 241 231
rect 207 61 241 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 47 597 81 631
rect 121 523 155 557
rect 121 227 155 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 286 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 286 1089
rect 0 1049 286 1055
rect 35 631 93 637
rect 35 597 47 631
rect 81 597 127 631
rect 35 591 93 597
rect 109 557 167 563
rect 109 523 121 557
rect 155 523 167 557
rect 109 517 167 523
rect 121 267 155 517
rect 109 261 167 267
rect 109 227 121 261
rect 155 227 167 261
rect 109 221 167 227
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 152 388 152 388 1 Y
port 1 n
rlabel viali 64 613 64 613 1 A
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
