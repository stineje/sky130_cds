* File: sky130_osu_sc_18T_hs__tbufi_l.spice
* Created: Thu Oct 29 17:10:09 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_hs__tbufi_l.pex.spice"
.subckt sky130_osu_sc_18T_hs__tbufi_l  GND VDD OE A Y
* 
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_OE_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1000 A_196_115# N_OE_M1000_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.1036 PD=0.95 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_196_115# N_GND_M1002_b NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VDD_M1005_d N_OE_M1005_g N_A_27_115#_M1005_s N_VDD_M1005_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1003 A_196_817# N_A_27_115#_M1003_g N_VDD_M1005_d N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.5 A=0.3 P=4.3 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g A_196_817# N_VDD_M1005_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.21 PD=4.53 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1005_b NWDIODE A=7.296 P=11.44
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__tbufi_l.pxi.spice"
*
.ends
*
*
