* File: sky130_osu_sc_12T_hs__addh_1.pxi.spice
* Created: Fri Nov 12 15:06:27 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%GND N_GND_M1007_d N_GND_M1002_d N_GND_M1007_b
+ N_GND_c_4_p N_GND_c_5_p N_GND_c_38_p N_GND_c_8_p GND N_GND_c_6_p
+ PM_SKY130_OSU_SC_12T_HS__ADDH_1%GND
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%VDD N_VDD_M1000_d N_VDD_M1003_d N_VDD_M1013_d
+ N_VDD_M1000_b N_VDD_c_106_p N_VDD_c_107_p N_VDD_c_120_p N_VDD_c_128_p
+ N_VDD_c_110_p N_VDD_c_113_p N_VDD_c_115_p VDD N_VDD_c_108_p
+ PM_SKY130_OSU_SC_12T_HS__ADDH_1%VDD
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%CON N_CON_M1011_d N_CON_M1013_s N_CON_M1009_d
+ N_CON_M1007_g N_CON_M1000_g N_CON_c_163_n N_CON_c_164_n N_CON_c_168_n
+ N_CON_c_170_n N_CON_c_201_n N_CON_c_171_n N_CON_c_172_n N_CON_c_173_n
+ N_CON_c_175_n N_CON_c_176_n N_CON_c_177_n N_CON_c_206_n N_CON_c_179_n
+ N_CON_c_181_n N_CON_c_182_n N_CON_c_183_n N_CON_c_186_n N_CON_c_188_n
+ N_CON_c_190_n N_CON_c_192_n N_CON_c_194_n CON
+ PM_SKY130_OSU_SC_12T_HS__ADDH_1%CON
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%B N_B_M1008_g N_B_M1001_g N_B_M1004_g
+ N_B_M1006_g N_B_c_312_n N_B_c_314_n N_B_c_315_n N_B_c_316_n N_B_c_317_n
+ N_B_c_318_n B PM_SKY130_OSU_SC_12T_HS__ADDH_1%B
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%A N_A_M1010_g N_A_M1003_g N_A_M1009_g
+ N_A_M1005_g N_A_c_412_n N_A_c_413_n N_A_c_414_n N_A_c_415_n N_A_c_416_n A
+ N_A_c_418_n PM_SKY130_OSU_SC_12T_HS__ADDH_1%A
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%A_208_521# N_A_208_521#_M1010_d
+ N_A_208_521#_M1001_d N_A_208_521#_c_493_n N_A_208_521#_M1012_g
+ N_A_208_521#_c_495_n N_A_208_521#_c_496_n N_A_208_521#_c_497_n
+ N_A_208_521#_M1002_g N_A_208_521#_c_501_n N_A_208_521#_c_503_n
+ N_A_208_521#_M1011_g N_A_208_521#_M1013_g N_A_208_521#_c_507_n
+ N_A_208_521#_c_508_n N_A_208_521#_c_509_n N_A_208_521#_c_523_n
+ N_A_208_521#_c_526_n N_A_208_521#_c_529_n N_A_208_521#_c_510_n
+ N_A_208_521#_c_513_n N_A_208_521#_c_514_n
+ PM_SKY130_OSU_SC_12T_HS__ADDH_1%A_208_521#
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%S N_S_M1007_s N_S_M1000_s N_S_c_606_n
+ N_S_c_614_n S N_S_c_611_n N_S_c_620_n PM_SKY130_OSU_SC_12T_HS__ADDH_1%S
x_PM_SKY130_OSU_SC_12T_HS__ADDH_1%CO N_CO_M1002_s N_CO_M1012_d N_CO_c_640_n
+ N_CO_c_649_n N_CO_c_643_n N_CO_c_646_n N_CO_c_647_n CO
+ PM_SKY130_OSU_SC_12T_HS__ADDH_1%CO
cc_1 N_GND_M1007_b N_CON_M1000_g 0.0588644f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_2 N_GND_M1007_b N_CON_c_163_n 0.0413766f $X=-0.045 $Y=0 $X2=0.35 $Y2=1.4
cc_3 N_GND_M1007_b N_CON_c_164_n 0.0224388f $X=-0.045 $Y=0 $X2=0.382 $Y2=1.235
cc_4 N_GND_c_4_p N_CON_c_164_n 0.00606474f $X=0.665 $Y=0.152 $X2=0.382 $Y2=1.235
cc_5 N_GND_c_5_p N_CON_c_164_n 0.0061123f $X=0.75 $Y=0.755 $X2=0.382 $Y2=1.235
cc_6 N_GND_c_6_p N_CON_c_164_n 0.00468827f $X=3.74 $Y=0.19 $X2=0.382 $Y2=1.235
cc_7 N_GND_M1007_b N_CON_c_168_n 3.10614e-19 $X=-0.045 $Y=0 $X2=2.62 $Y2=1.455
cc_8 N_GND_c_8_p N_CON_c_168_n 0.00333172f $X=2.56 $Y=0.755 $X2=2.62 $Y2=1.455
cc_9 N_GND_M1007_b N_CON_c_170_n 0.0156018f $X=-0.045 $Y=0 $X2=2.62 $Y2=2.385
cc_10 N_GND_M1007_b N_CON_c_171_n 0.00849691f $X=-0.045 $Y=0 $X2=3.335 $Y2=1.37
cc_11 N_GND_M1007_b N_CON_c_172_n 0.0112921f $X=-0.045 $Y=0 $X2=3.755 $Y2=2.47
cc_12 N_GND_M1007_b N_CON_c_173_n 0.0123217f $X=-0.045 $Y=0 $X2=3.335 $Y2=0.635
cc_13 N_GND_c_6_p N_CON_c_173_n 0.00708954f $X=3.74 $Y=0.19 $X2=3.335 $Y2=0.635
cc_14 N_GND_M1007_b N_CON_c_175_n 0.00433753f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.285
cc_15 N_GND_M1007_b N_CON_c_176_n 0.00334447f $X=-0.045 $Y=0 $X2=3.42 $Y2=0.755
cc_16 N_GND_M1007_b N_CON_c_177_n 0.0122917f $X=-0.045 $Y=0 $X2=3.765 $Y2=0.635
cc_17 N_GND_c_6_p N_CON_c_177_n 0.00708954f $X=3.74 $Y=0.19 $X2=3.765 $Y2=0.635
cc_18 N_GND_M1007_b N_CON_c_179_n 0.00654377f $X=-0.045 $Y=0 $X2=0.635 $Y2=1.37
cc_19 N_GND_c_5_p N_CON_c_179_n 0.00183327f $X=0.75 $Y=0.755 $X2=0.635 $Y2=1.37
cc_20 N_GND_M1007_b N_CON_c_181_n 0.00269067f $X=-0.045 $Y=0 $X2=0.55 $Y2=1.385
cc_21 N_GND_M1007_b N_CON_c_182_n 2.79926e-19 $X=-0.045 $Y=0 $X2=2.62 $Y2=2.47
cc_22 N_GND_M1007_b N_CON_c_183_n 0.00977498f $X=-0.045 $Y=0 $X2=2.99 $Y2=0.635
cc_23 N_GND_c_8_p N_CON_c_183_n 0.00134209f $X=2.56 $Y=0.755 $X2=2.99 $Y2=0.635
cc_24 N_GND_c_6_p N_CON_c_183_n 0.00474945f $X=3.74 $Y=0.19 $X2=2.99 $Y2=0.635
cc_25 N_GND_M1007_b N_CON_c_186_n 0.0102363f $X=-0.045 $Y=0 $X2=3.42 $Y2=0.635
cc_26 N_GND_c_6_p N_CON_c_186_n 0.0048888f $X=3.74 $Y=0.19 $X2=3.42 $Y2=0.635
cc_27 N_GND_M1007_b N_CON_c_188_n 0.0104745f $X=-0.045 $Y=0 $X2=3.85 $Y2=0.635
cc_28 N_GND_c_6_p N_CON_c_188_n 0.00474945f $X=3.74 $Y=0.19 $X2=3.85 $Y2=0.635
cc_29 N_GND_M1007_b N_CON_c_190_n 0.0196895f $X=-0.045 $Y=0 $X2=2.475 $Y2=1.37
cc_30 N_GND_c_5_p N_CON_c_190_n 0.00237883f $X=0.75 $Y=0.755 $X2=2.475 $Y2=1.37
cc_31 N_GND_M1007_b N_CON_c_192_n 0.0134764f $X=-0.045 $Y=0 $X2=0.78 $Y2=1.37
cc_32 N_GND_c_5_p N_CON_c_192_n 0.00429244f $X=0.75 $Y=0.755 $X2=0.78 $Y2=1.37
cc_33 N_GND_M1007_b N_CON_c_194_n 0.00124672f $X=-0.045 $Y=0 $X2=2.62 $Y2=1.37
cc_34 N_GND_c_8_p N_CON_c_194_n 0.00508608f $X=2.56 $Y=0.755 $X2=2.62 $Y2=1.37
cc_35 N_GND_M1007_b CON 0.00374951f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.37
cc_36 N_GND_M1007_b N_B_M1008_g 0.0329711f $X=-0.045 $Y=0 $X2=0.965 $Y2=0.85
cc_37 N_GND_c_5_p N_B_M1008_g 0.00318344f $X=0.75 $Y=0.755 $X2=0.965 $Y2=0.85
cc_38 N_GND_c_38_p N_B_M1008_g 0.00606474f $X=2.475 $Y=0.152 $X2=0.965 $Y2=0.85
cc_39 N_GND_c_6_p N_B_M1008_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.965 $Y2=0.85
cc_40 N_GND_M1007_b N_B_M1001_g 0.0282323f $X=-0.045 $Y=0 $X2=0.965 $Y2=3.235
cc_41 N_GND_M1007_b N_B_M1004_g 0.0385592f $X=-0.045 $Y=0 $X2=3.205 $Y2=0.85
cc_42 N_GND_c_6_p N_B_M1004_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.205 $Y2=0.85
cc_43 N_GND_M1007_b N_B_M1006_g 0.0272084f $X=-0.045 $Y=0 $X2=3.265 $Y2=3.235
cc_44 N_GND_M1007_b N_B_c_312_n 0.0279691f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.74
cc_45 N_GND_c_5_p N_B_c_312_n 0.00173465f $X=0.75 $Y=0.755 $X2=0.905 $Y2=1.74
cc_46 N_GND_M1007_b N_B_c_314_n 0.0299556f $X=-0.045 $Y=0 $X2=3.205 $Y2=1.74
cc_47 N_GND_M1007_b N_B_c_315_n 0.00407254f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.74
cc_48 N_GND_M1007_b N_B_c_316_n 0.00365598f $X=-0.045 $Y=0 $X2=3.205 $Y2=1.74
cc_49 N_GND_M1007_b N_B_c_317_n 0.00206723f $X=-0.045 $Y=0 $X2=1.05 $Y2=1.74
cc_50 N_GND_M1007_b N_B_c_318_n 0.0175509f $X=-0.045 $Y=0 $X2=3.06 $Y2=1.74
cc_51 N_GND_M1007_b B 0.00164195f $X=-0.045 $Y=0 $X2=3.21 $Y2=1.74
cc_52 N_GND_M1007_b N_A_M1010_g 0.0542089f $X=-0.045 $Y=0 $X2=1.325 $Y2=0.85
cc_53 N_GND_c_38_p N_A_M1010_g 0.00606474f $X=2.475 $Y=0.152 $X2=1.325 $Y2=0.85
cc_54 N_GND_c_6_p N_A_M1010_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.325 $Y2=0.85
cc_55 N_GND_M1007_b N_A_M1003_g 0.00835457f $X=-0.045 $Y=0 $X2=1.395 $Y2=3.235
cc_56 N_GND_M1007_b N_A_M1009_g 0.0108664f $X=-0.045 $Y=0 $X2=3.625 $Y2=3.235
cc_57 N_GND_M1007_b N_A_M1005_g 0.0831928f $X=-0.045 $Y=0 $X2=3.635 $Y2=0.85
cc_58 N_GND_c_6_p N_A_M1005_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.635 $Y2=0.85
cc_59 N_GND_M1007_b N_A_c_412_n 0.0253796f $X=-0.045 $Y=0 $X2=1.385 $Y2=2.11
cc_60 N_GND_M1007_b N_A_c_413_n 0.034256f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.11
cc_61 N_GND_M1007_b N_A_c_414_n 9.49347e-19 $X=-0.045 $Y=0 $X2=1.385 $Y2=2.11
cc_62 N_GND_M1007_b N_A_c_415_n 0.00995238f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.11
cc_63 N_GND_M1007_b N_A_c_416_n 0.00430309f $X=-0.045 $Y=0 $X2=1.53 $Y2=2.11
cc_64 N_GND_M1007_b A 0.00380188f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.11
cc_65 N_GND_M1007_b N_A_c_418_n 0.0115394f $X=-0.045 $Y=0 $X2=3.54 $Y2=2.11
cc_66 N_GND_M1007_b N_A_208_521#_c_493_n 0.0270254f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=2.115
cc_67 N_GND_M1007_b N_A_208_521#_M1012_g 0.00928694f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=3.235
cc_68 N_GND_M1007_b N_A_208_521#_c_495_n 0.0169485f $X=-0.045 $Y=0 $X2=2.21
+ $Y2=1.32
cc_69 N_GND_M1007_b N_A_208_521#_c_496_n 0.0619559f $X=-0.045 $Y=0 $X2=2.76
+ $Y2=2.19
cc_70 N_GND_M1007_b N_A_208_521#_c_497_n 0.0222111f $X=-0.045 $Y=0 $X2=2.285
+ $Y2=1.245
cc_71 N_GND_c_38_p N_A_208_521#_c_497_n 0.00558991f $X=2.475 $Y=0.152 $X2=2.285
+ $Y2=1.245
cc_72 N_GND_c_8_p N_A_208_521#_c_497_n 0.00608877f $X=2.56 $Y=0.755 $X2=2.285
+ $Y2=1.245
cc_73 N_GND_c_6_p N_A_208_521#_c_497_n 0.00468827f $X=3.74 $Y=0.19 $X2=2.285
+ $Y2=1.245
cc_74 N_GND_M1007_b N_A_208_521#_c_501_n 0.0264701f $X=-0.045 $Y=0 $X2=2.7
+ $Y2=1.32
cc_75 N_GND_c_8_p N_A_208_521#_c_501_n 0.00351744f $X=2.56 $Y=0.755 $X2=2.7
+ $Y2=1.32
cc_76 N_GND_M1007_b N_A_208_521#_c_503_n 0.023503f $X=-0.045 $Y=0 $X2=2.775
+ $Y2=1.245
cc_77 N_GND_c_8_p N_A_208_521#_c_503_n 0.00280941f $X=2.56 $Y=0.755 $X2=2.775
+ $Y2=1.245
cc_78 N_GND_c_6_p N_A_208_521#_c_503_n 0.00468827f $X=3.74 $Y=0.19 $X2=2.775
+ $Y2=1.245
cc_79 N_GND_M1007_b N_A_208_521#_M1013_g 0.00900107f $X=-0.045 $Y=0 $X2=2.835
+ $Y2=3.235
cc_80 N_GND_M1007_b N_A_208_521#_c_507_n 0.0385573f $X=-0.045 $Y=0 $X2=1.825
+ $Y2=1.32
cc_81 N_GND_M1007_b N_A_208_521#_c_508_n 0.00492701f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=2.19
cc_82 N_GND_M1007_b N_A_208_521#_c_509_n 0.0061448f $X=-0.045 $Y=0 $X2=2.285
+ $Y2=1.32
cc_83 N_GND_M1007_b N_A_208_521#_c_510_n 0.00551537f $X=-0.045 $Y=0 $X2=1.54
+ $Y2=0.755
cc_84 N_GND_c_38_p N_A_208_521#_c_510_n 0.00741243f $X=2.475 $Y=0.152 $X2=1.54
+ $Y2=0.755
cc_85 N_GND_c_6_p N_A_208_521#_c_510_n 0.00476261f $X=3.74 $Y=0.19 $X2=1.54
+ $Y2=0.755
cc_86 N_GND_M1007_b N_A_208_521#_c_513_n 0.0137594f $X=-0.045 $Y=0 $X2=1.725
+ $Y2=2.445
cc_87 N_GND_M1007_b N_A_208_521#_c_514_n 0.00684174f $X=-0.045 $Y=0 $X2=1.725
+ $Y2=1.475
cc_88 N_GND_M1007_b N_S_c_606_n 0.001552f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.755
cc_89 N_GND_c_4_p N_S_c_606_n 0.00720145f $X=0.665 $Y=0.152 $X2=0.26 $Y2=0.755
cc_90 N_GND_c_5_p N_S_c_606_n 0.00826522f $X=0.75 $Y=0.755 $X2=0.26 $Y2=0.755
cc_91 N_GND_c_6_p N_S_c_606_n 0.00471702f $X=3.74 $Y=0.19 $X2=0.26 $Y2=0.755
cc_92 N_GND_M1007_b S 0.0627303f $X=-0.045 $Y=0 $X2=0.25 $Y2=1.905
cc_93 N_GND_M1007_b N_S_c_611_n 0.00973258f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.995
cc_94 N_GND_c_4_p N_S_c_611_n 0.00255092f $X=0.665 $Y=0.152 $X2=0.26 $Y2=0.995
cc_95 N_GND_c_5_p N_S_c_611_n 0.00132248f $X=0.75 $Y=0.755 $X2=0.26 $Y2=0.995
cc_96 N_GND_M1007_b N_CO_c_640_n 0.00153988f $X=-0.045 $Y=0 $X2=2.07 $Y2=0.755
cc_97 N_GND_c_38_p N_CO_c_640_n 0.00719884f $X=2.475 $Y=0.152 $X2=2.07 $Y2=0.755
cc_98 N_GND_c_6_p N_CO_c_640_n 0.00465624f $X=3.74 $Y=0.19 $X2=2.07 $Y2=0.755
cc_99 N_GND_c_38_p N_CO_c_643_n 0.00116296f $X=2.475 $Y=0.152 $X2=2.175
+ $Y2=0.992
cc_100 N_GND_c_8_p N_CO_c_643_n 0.00176942f $X=2.56 $Y=0.755 $X2=2.175 $Y2=0.992
cc_101 N_GND_c_6_p N_CO_c_643_n 0.0022687f $X=3.74 $Y=0.19 $X2=2.175 $Y2=0.992
cc_102 N_GND_M1007_b N_CO_c_646_n 0.00130468f $X=-0.045 $Y=0 $X2=2.175 $Y2=2.48
cc_103 N_GND_M1007_b N_CO_c_647_n 0.0155801f $X=-0.045 $Y=0 $X2=2.137 $Y2=2.395
cc_104 N_GND_M1007_b CO 0.00219851f $X=-0.045 $Y=0 $X2=2.175 $Y2=2.48
cc_105 N_VDD_M1000_b N_CON_M1000_g 0.0274231f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_106 N_VDD_c_106_p N_CON_M1000_g 0.00606474f $X=0.665 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_107 N_VDD_c_107_p N_CON_M1000_g 0.0129275f $X=0.75 $Y=2.955 $X2=0.475
+ $Y2=3.235
cc_108 N_VDD_c_108_p N_CON_M1000_g 0.00468827f $X=3.74 $Y=4.25 $X2=0.475
+ $Y2=3.235
cc_109 N_VDD_M1000_b N_CON_c_201_n 0.0024633f $X=-0.045 $Y=2.425 $X2=2.62
+ $Y2=2.955
cc_110 N_VDD_c_110_p N_CON_c_201_n 0.00751506f $X=2.965 $Y=4.287 $X2=2.62
+ $Y2=2.955
cc_111 N_VDD_c_108_p N_CON_c_201_n 0.00476261f $X=3.74 $Y=4.25 $X2=2.62
+ $Y2=2.955
cc_112 N_VDD_M1000_b N_CON_c_172_n 0.0218233f $X=-0.045 $Y=2.425 $X2=3.755
+ $Y2=2.47
cc_113 N_VDD_c_113_p N_CON_c_172_n 0.0133353f $X=3.05 $Y=2.955 $X2=3.755
+ $Y2=2.47
cc_114 N_VDD_M1000_b N_CON_c_206_n 0.00375952f $X=-0.045 $Y=2.425 $X2=3.84
+ $Y2=2.955
cc_115 N_VDD_c_115_p N_CON_c_206_n 0.00736239f $X=3.74 $Y=4.22 $X2=3.84
+ $Y2=2.955
cc_116 N_VDD_c_108_p N_CON_c_206_n 0.00476261f $X=3.74 $Y=4.25 $X2=3.84
+ $Y2=2.955
cc_117 N_VDD_M1000_b N_CON_c_182_n 0.00108117f $X=-0.045 $Y=2.425 $X2=2.62
+ $Y2=2.47
cc_118 N_VDD_M1000_b N_B_M1001_g 0.0212391f $X=-0.045 $Y=2.425 $X2=0.965
+ $Y2=3.235
cc_119 N_VDD_c_107_p N_B_M1001_g 0.00353221f $X=0.75 $Y=2.955 $X2=0.965
+ $Y2=3.235
cc_120 N_VDD_c_120_p N_B_M1001_g 0.00606474f $X=1.525 $Y=4.287 $X2=0.965
+ $Y2=3.235
cc_121 N_VDD_c_108_p N_B_M1001_g 0.00468827f $X=3.74 $Y=4.25 $X2=0.965 $Y2=3.235
cc_122 N_VDD_M1000_b N_B_M1006_g 0.0181844f $X=-0.045 $Y=2.425 $X2=3.265
+ $Y2=3.235
cc_123 N_VDD_c_113_p N_B_M1006_g 0.00337744f $X=3.05 $Y=2.955 $X2=3.265
+ $Y2=3.235
cc_124 N_VDD_c_115_p N_B_M1006_g 0.00606474f $X=3.74 $Y=4.22 $X2=3.265 $Y2=3.235
cc_125 N_VDD_c_108_p N_B_M1006_g 0.00468827f $X=3.74 $Y=4.25 $X2=3.265 $Y2=3.235
cc_126 N_VDD_M1000_b N_A_M1003_g 0.019386f $X=-0.045 $Y=2.425 $X2=1.395
+ $Y2=3.235
cc_127 N_VDD_c_120_p N_A_M1003_g 0.00606474f $X=1.525 $Y=4.287 $X2=1.395
+ $Y2=3.235
cc_128 N_VDD_c_128_p N_A_M1003_g 0.00353221f $X=1.61 $Y=3.295 $X2=1.395
+ $Y2=3.235
cc_129 N_VDD_c_108_p N_A_M1003_g 0.00468827f $X=3.74 $Y=4.25 $X2=1.395 $Y2=3.235
cc_130 N_VDD_M1000_b N_A_M1009_g 0.0239507f $X=-0.045 $Y=2.425 $X2=3.625
+ $Y2=3.235
cc_131 N_VDD_c_115_p N_A_M1009_g 0.00606474f $X=3.74 $Y=4.22 $X2=3.625 $Y2=3.235
cc_132 N_VDD_c_108_p N_A_M1009_g 0.00468827f $X=3.74 $Y=4.25 $X2=3.625 $Y2=3.235
cc_133 N_VDD_M1000_b N_A_208_521#_M1012_g 0.0243727f $X=-0.045 $Y=2.425
+ $X2=1.885 $Y2=3.235
cc_134 N_VDD_c_128_p N_A_208_521#_M1012_g 0.00995677f $X=1.61 $Y=3.295 $X2=1.885
+ $Y2=3.235
cc_135 N_VDD_c_110_p N_A_208_521#_M1012_g 0.00606474f $X=2.965 $Y=4.287
+ $X2=1.885 $Y2=3.235
cc_136 N_VDD_c_108_p N_A_208_521#_M1012_g 0.00468827f $X=3.74 $Y=4.25 $X2=1.885
+ $Y2=3.235
cc_137 N_VDD_M1000_b N_A_208_521#_M1013_g 0.0248258f $X=-0.045 $Y=2.425
+ $X2=2.835 $Y2=3.235
cc_138 N_VDD_c_110_p N_A_208_521#_M1013_g 0.00606474f $X=2.965 $Y=4.287
+ $X2=2.835 $Y2=3.235
cc_139 N_VDD_c_113_p N_A_208_521#_M1013_g 0.00337744f $X=3.05 $Y=2.955 $X2=2.835
+ $Y2=3.235
cc_140 N_VDD_c_108_p N_A_208_521#_M1013_g 0.00468827f $X=3.74 $Y=4.25 $X2=2.835
+ $Y2=3.235
cc_141 N_VDD_M1000_b N_A_208_521#_c_523_n 0.00155118f $X=-0.045 $Y=2.425
+ $X2=1.18 $Y2=3.295
cc_142 N_VDD_c_120_p N_A_208_521#_c_523_n 0.0073901f $X=1.525 $Y=4.287 $X2=1.18
+ $Y2=3.295
cc_143 N_VDD_c_108_p N_A_208_521#_c_523_n 0.00475776f $X=3.74 $Y=4.25 $X2=1.18
+ $Y2=3.295
cc_144 N_VDD_M1003_d N_A_208_521#_c_526_n 0.00559263f $X=1.47 $Y=2.605 $X2=1.64
+ $Y2=2.53
cc_145 N_VDD_M1000_b N_A_208_521#_c_526_n 0.00273697f $X=-0.045 $Y=2.425
+ $X2=1.64 $Y2=2.53
cc_146 N_VDD_c_128_p N_A_208_521#_c_526_n 0.00681335f $X=1.61 $Y=3.295 $X2=1.64
+ $Y2=2.53
cc_147 N_VDD_M1000_b N_A_208_521#_c_529_n 0.00518782f $X=-0.045 $Y=2.425
+ $X2=1.265 $Y2=2.53
cc_148 N_VDD_M1000_b N_A_208_521#_c_513_n 3.89739e-19 $X=-0.045 $Y=2.425
+ $X2=1.725 $Y2=2.445
cc_149 N_VDD_M1000_b N_S_c_614_n 0.00156053f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=2.85
cc_150 N_VDD_c_106_p N_S_c_614_n 0.00736239f $X=0.665 $Y=4.287 $X2=0.26 $Y2=2.85
cc_151 N_VDD_c_107_p N_S_c_614_n 0.0262407f $X=0.75 $Y=2.955 $X2=0.26 $Y2=2.85
cc_152 N_VDD_c_108_p N_S_c_614_n 0.00476261f $X=3.74 $Y=4.25 $X2=0.26 $Y2=2.85
cc_153 N_VDD_M1000_b S 0.00951645f $X=-0.045 $Y=2.425 $X2=0.25 $Y2=1.905
cc_154 N_VDD_c_107_p S 2.19343e-19 $X=0.75 $Y=2.955 $X2=0.25 $Y2=1.905
cc_155 N_VDD_M1000_b N_S_c_620_n 0.0102428f $X=-0.045 $Y=2.425 $X2=0.26 $Y2=2.85
cc_156 N_VDD_c_107_p N_S_c_620_n 0.00553039f $X=0.75 $Y=2.955 $X2=0.26 $Y2=2.85
cc_157 N_VDD_M1000_b N_CO_c_649_n 0.00231154f $X=-0.045 $Y=2.425 $X2=2.1
+ $Y2=2.955
cc_158 N_VDD_c_110_p N_CO_c_649_n 0.00756638f $X=2.965 $Y=4.287 $X2=2.1
+ $Y2=2.955
cc_159 N_VDD_c_108_p N_CO_c_649_n 0.00476261f $X=3.74 $Y=4.25 $X2=2.1 $Y2=2.955
cc_160 N_VDD_M1000_b N_CO_c_646_n 0.00360959f $X=-0.045 $Y=2.425 $X2=2.175
+ $Y2=2.48
cc_161 N_VDD_M1000_b CO 0.0105263f $X=-0.045 $Y=2.425 $X2=2.175 $Y2=2.48
cc_162 N_CON_c_164_n N_B_M1008_g 0.0329987f $X=0.382 $Y=1.235 $X2=0.965 $Y2=0.85
cc_163 N_CON_c_179_n N_B_M1008_g 0.00371117f $X=0.635 $Y=1.37 $X2=0.965 $Y2=0.85
cc_164 N_CON_c_190_n N_B_M1008_g 0.0103778f $X=2.475 $Y=1.37 $X2=0.965 $Y2=0.85
cc_165 N_CON_c_192_n N_B_M1008_g 9.80511e-19 $X=0.78 $Y=1.37 $X2=0.965 $Y2=0.85
cc_166 N_CON_M1000_g N_B_M1001_g 0.0512242f $X=0.475 $Y=3.235 $X2=0.965
+ $Y2=3.235
cc_167 N_CON_c_170_n N_B_M1004_g 0.00298059f $X=2.62 $Y=2.385 $X2=3.205 $Y2=0.85
cc_168 N_CON_c_171_n N_B_M1004_g 0.0111215f $X=3.335 $Y=1.37 $X2=3.205 $Y2=0.85
cc_169 N_CON_c_173_n N_B_M1004_g 0.00781392f $X=3.335 $Y=0.635 $X2=3.205
+ $Y2=0.85
cc_170 N_CON_c_176_n N_B_M1004_g 0.00441254f $X=3.42 $Y=0.755 $X2=3.205 $Y2=0.85
cc_171 N_CON_c_194_n N_B_M1004_g 4.77705e-19 $X=2.62 $Y=1.37 $X2=3.205 $Y2=0.85
cc_172 CON N_B_M1004_g 0.00323231f $X=3.42 $Y=1.37 $X2=3.205 $Y2=0.85
cc_173 N_CON_c_170_n N_B_M1006_g 0.00509671f $X=2.62 $Y=2.385 $X2=3.265
+ $Y2=3.235
cc_174 N_CON_c_172_n N_B_M1006_g 0.0160357f $X=3.755 $Y=2.47 $X2=3.265 $Y2=3.235
cc_175 N_CON_M1000_g N_B_c_312_n 0.0198105f $X=0.475 $Y=3.235 $X2=0.905 $Y2=1.74
cc_176 N_CON_c_190_n N_B_c_312_n 0.0017113f $X=2.475 $Y=1.37 $X2=0.905 $Y2=1.74
cc_177 N_CON_c_170_n N_B_c_314_n 0.00527976f $X=2.62 $Y=2.385 $X2=3.205 $Y2=1.74
cc_178 N_CON_c_171_n N_B_c_314_n 0.00297725f $X=3.335 $Y=1.37 $X2=3.205 $Y2=1.74
cc_179 N_CON_c_172_n N_B_c_314_n 0.00235541f $X=3.755 $Y=2.47 $X2=3.205 $Y2=1.74
cc_180 CON N_B_c_314_n 0.00117979f $X=3.42 $Y=1.37 $X2=3.205 $Y2=1.74
cc_181 N_CON_M1000_g N_B_c_315_n 0.00376362f $X=0.475 $Y=3.235 $X2=0.905
+ $Y2=1.74
cc_182 N_CON_c_190_n N_B_c_315_n 0.00387996f $X=2.475 $Y=1.37 $X2=0.905 $Y2=1.74
cc_183 N_CON_c_192_n N_B_c_315_n 0.00117441f $X=0.78 $Y=1.37 $X2=0.905 $Y2=1.74
cc_184 N_CON_c_170_n N_B_c_316_n 0.00612449f $X=2.62 $Y=2.385 $X2=3.205 $Y2=1.74
cc_185 N_CON_c_171_n N_B_c_316_n 0.0159093f $X=3.335 $Y=1.37 $X2=3.205 $Y2=1.74
cc_186 N_CON_c_172_n N_B_c_316_n 0.00416532f $X=3.755 $Y=2.47 $X2=3.205 $Y2=1.74
cc_187 N_CON_c_175_n N_B_c_316_n 0.00205373f $X=3.42 $Y=1.285 $X2=3.205 $Y2=1.74
cc_188 CON N_B_c_316_n 9.81883e-19 $X=3.42 $Y=1.37 $X2=3.205 $Y2=1.74
cc_189 N_CON_M1000_g N_B_c_317_n 3.21736e-19 $X=0.475 $Y=3.235 $X2=1.05 $Y2=1.74
cc_190 N_CON_c_190_n N_B_c_317_n 0.024704f $X=2.475 $Y=1.37 $X2=1.05 $Y2=1.74
cc_191 N_CON_c_192_n N_B_c_317_n 0.002062f $X=0.78 $Y=1.37 $X2=1.05 $Y2=1.74
cc_192 N_CON_c_170_n N_B_c_318_n 0.0139119f $X=2.62 $Y=2.385 $X2=3.06 $Y2=1.74
cc_193 N_CON_c_171_n N_B_c_318_n 0.0132985f $X=3.335 $Y=1.37 $X2=3.06 $Y2=1.74
cc_194 N_CON_c_190_n N_B_c_318_n 0.116608f $X=2.475 $Y=1.37 $X2=3.06 $Y2=1.74
cc_195 N_CON_c_194_n N_B_c_318_n 0.0254758f $X=2.62 $Y=1.37 $X2=3.06 $Y2=1.74
cc_196 N_CON_c_170_n B 0.00223952f $X=2.62 $Y=2.385 $X2=3.21 $Y2=1.74
cc_197 N_CON_c_171_n B 0.00321159f $X=3.335 $Y=1.37 $X2=3.21 $Y2=1.74
cc_198 CON B 0.0176994f $X=3.42 $Y=1.37 $X2=3.21 $Y2=1.74
cc_199 N_CON_c_190_n N_A_M1010_g 0.0102863f $X=2.475 $Y=1.37 $X2=1.325 $Y2=0.85
cc_200 N_CON_c_172_n N_A_M1009_g 0.015762f $X=3.755 $Y=2.47 $X2=3.625 $Y2=3.235
cc_201 N_CON_c_206_n N_A_M1009_g 0.00554073f $X=3.84 $Y=2.955 $X2=3.625
+ $Y2=3.235
cc_202 N_CON_c_175_n N_A_M1005_g 0.00402015f $X=3.42 $Y=1.285 $X2=3.635 $Y2=0.85
cc_203 N_CON_c_176_n N_A_M1005_g 0.00441254f $X=3.42 $Y=0.755 $X2=3.635 $Y2=0.85
cc_204 N_CON_c_177_n N_A_M1005_g 0.0107657f $X=3.765 $Y=0.635 $X2=3.635 $Y2=0.85
cc_205 N_CON_c_188_n N_A_M1005_g 2.14912e-19 $X=3.85 $Y=0.635 $X2=3.635 $Y2=0.85
cc_206 CON N_A_M1005_g 0.0104932f $X=3.42 $Y=1.37 $X2=3.635 $Y2=0.85
cc_207 N_CON_c_172_n N_A_c_413_n 0.00303009f $X=3.755 $Y=2.47 $X2=3.685 $Y2=2.11
cc_208 N_CON_c_172_n N_A_c_415_n 0.0189273f $X=3.755 $Y=2.47 $X2=3.685 $Y2=2.11
cc_209 CON N_A_c_415_n 3.86961e-19 $X=3.42 $Y=1.37 $X2=3.685 $Y2=2.11
cc_210 N_CON_c_172_n A 0.00711502f $X=3.755 $Y=2.47 $X2=3.685 $Y2=2.11
cc_211 CON A 0.00132366f $X=3.42 $Y=1.37 $X2=3.685 $Y2=2.11
cc_212 N_CON_c_170_n N_A_c_418_n 0.0228959f $X=2.62 $Y=2.385 $X2=3.54 $Y2=2.11
cc_213 N_CON_c_172_n N_A_c_418_n 0.0305931f $X=3.755 $Y=2.47 $X2=3.54 $Y2=2.11
cc_214 N_CON_c_175_n N_A_c_418_n 8.38986e-19 $X=3.42 $Y=1.285 $X2=3.54 $Y2=2.11
cc_215 CON N_A_c_418_n 0.0098042f $X=3.42 $Y=1.37 $X2=3.54 $Y2=2.11
cc_216 N_CON_c_190_n N_A_208_521#_c_495_n 0.00235551f $X=2.475 $Y=1.37 $X2=2.21
+ $Y2=1.32
cc_217 N_CON_c_170_n N_A_208_521#_c_496_n 0.0141734f $X=2.62 $Y=2.385 $X2=2.76
+ $Y2=2.19
cc_218 N_CON_c_171_n N_A_208_521#_c_496_n 0.00258433f $X=3.335 $Y=1.37 $X2=2.76
+ $Y2=2.19
cc_219 N_CON_c_168_n N_A_208_521#_c_501_n 0.00895457f $X=2.62 $Y=1.455 $X2=2.7
+ $Y2=1.32
cc_220 N_CON_c_171_n N_A_208_521#_c_501_n 0.00965528f $X=3.335 $Y=1.37 $X2=2.7
+ $Y2=1.32
cc_221 N_CON_c_190_n N_A_208_521#_c_501_n 0.00550578f $X=2.475 $Y=1.37 $X2=2.7
+ $Y2=1.32
cc_222 N_CON_c_194_n N_A_208_521#_c_501_n 0.00766294f $X=2.62 $Y=1.37 $X2=2.7
+ $Y2=1.32
cc_223 N_CON_c_183_n N_A_208_521#_c_503_n 2.0295e-19 $X=2.99 $Y=0.635 $X2=2.775
+ $Y2=1.245
cc_224 N_CON_c_170_n N_A_208_521#_M1013_g 0.0046186f $X=2.62 $Y=2.385 $X2=2.835
+ $Y2=3.235
cc_225 N_CON_c_201_n N_A_208_521#_M1013_g 0.00554073f $X=2.62 $Y=2.955 $X2=2.835
+ $Y2=3.235
cc_226 N_CON_c_172_n N_A_208_521#_M1013_g 0.0162813f $X=3.755 $Y=2.47 $X2=2.835
+ $Y2=3.235
cc_227 N_CON_c_190_n N_A_208_521#_c_507_n 0.0103832f $X=2.475 $Y=1.37 $X2=1.825
+ $Y2=1.32
cc_228 N_CON_c_190_n N_A_208_521#_c_509_n 0.00472068f $X=2.475 $Y=1.37 $X2=2.285
+ $Y2=1.32
cc_229 N_CON_c_190_n N_A_208_521#_c_510_n 0.0108903f $X=2.475 $Y=1.37 $X2=1.54
+ $Y2=0.755
cc_230 N_CON_c_190_n N_A_208_521#_c_514_n 0.0233954f $X=2.475 $Y=1.37 $X2=1.725
+ $Y2=1.475
cc_231 N_CON_c_163_n N_S_c_606_n 0.00232333f $X=0.35 $Y=1.4 $X2=0.26 $Y2=0.755
cc_232 N_CON_c_164_n N_S_c_606_n 0.00346767f $X=0.382 $Y=1.235 $X2=0.26
+ $Y2=0.755
cc_233 N_CON_c_181_n N_S_c_606_n 0.00772296f $X=0.55 $Y=1.385 $X2=0.26 $Y2=0.755
cc_234 N_CON_M1000_g N_S_c_614_n 0.00424545f $X=0.475 $Y=3.235 $X2=0.26 $Y2=2.85
cc_235 N_CON_M1000_g S 0.0254249f $X=0.475 $Y=3.235 $X2=0.25 $Y2=1.905
cc_236 N_CON_c_163_n S 0.00737454f $X=0.35 $Y=1.4 $X2=0.25 $Y2=1.905
cc_237 N_CON_c_164_n S 0.00289801f $X=0.382 $Y=1.235 $X2=0.25 $Y2=1.905
cc_238 N_CON_c_179_n S 3.89614e-19 $X=0.635 $Y=1.37 $X2=0.25 $Y2=1.905
cc_239 N_CON_c_181_n S 0.0146482f $X=0.55 $Y=1.385 $X2=0.25 $Y2=1.905
cc_240 N_CON_c_192_n S 0.0220159f $X=0.78 $Y=1.37 $X2=0.25 $Y2=1.905
cc_241 N_CON_c_163_n N_S_c_611_n 0.00146137f $X=0.35 $Y=1.4 $X2=0.26 $Y2=0.995
cc_242 N_CON_c_164_n N_S_c_611_n 0.00567218f $X=0.382 $Y=1.235 $X2=0.26
+ $Y2=0.995
cc_243 N_CON_c_181_n N_S_c_611_n 0.0025199f $X=0.55 $Y=1.385 $X2=0.26 $Y2=0.995
cc_244 N_CON_M1000_g N_S_c_620_n 0.00263349f $X=0.475 $Y=3.235 $X2=0.26 $Y2=2.85
cc_245 N_CON_c_201_n N_CO_c_649_n 0.0551753f $X=2.62 $Y=2.955 $X2=2.1 $Y2=2.955
cc_246 N_CON_c_190_n N_CO_c_643_n 0.00507808f $X=2.475 $Y=1.37 $X2=2.175
+ $Y2=0.992
cc_247 N_CON_c_201_n N_CO_c_646_n 3.73019e-19 $X=2.62 $Y=2.955 $X2=2.175
+ $Y2=2.48
cc_248 N_CON_c_168_n N_CO_c_647_n 0.00688689f $X=2.62 $Y=1.455 $X2=2.137
+ $Y2=2.395
cc_249 N_CON_c_170_n N_CO_c_647_n 0.0448782f $X=2.62 $Y=2.385 $X2=2.137
+ $Y2=2.395
cc_250 N_CON_c_182_n N_CO_c_647_n 0.00730853f $X=2.62 $Y=2.47 $X2=2.137
+ $Y2=2.395
cc_251 N_CON_c_190_n N_CO_c_647_n 0.0122208f $X=2.475 $Y=1.37 $X2=2.137
+ $Y2=2.395
cc_252 N_CON_c_194_n N_CO_c_647_n 0.00203433f $X=2.62 $Y=1.37 $X2=2.137
+ $Y2=2.395
cc_253 N_CON_c_170_n CO 5.70376e-19 $X=2.62 $Y=2.385 $X2=2.175 $Y2=2.48
cc_254 N_CON_c_201_n CO 0.00122973f $X=2.62 $Y=2.955 $X2=2.175 $Y2=2.48
cc_255 N_CON_c_182_n CO 0.00605606f $X=2.62 $Y=2.47 $X2=2.175 $Y2=2.48
cc_256 N_B_M1008_g N_A_M1010_g 0.0576612f $X=0.965 $Y=0.85 $X2=1.325 $Y2=0.85
cc_257 N_B_c_315_n N_A_M1010_g 0.00121678f $X=0.905 $Y=1.74 $X2=1.325 $Y2=0.85
cc_258 N_B_c_317_n N_A_M1010_g 7.94897e-19 $X=1.05 $Y=1.74 $X2=1.325 $Y2=0.85
cc_259 N_B_c_318_n N_A_M1010_g 0.00595709f $X=3.06 $Y=1.74 $X2=1.325 $Y2=0.85
cc_260 N_B_M1001_g N_A_M1003_g 0.0384449f $X=0.965 $Y=3.235 $X2=1.395 $Y2=3.235
cc_261 N_B_M1004_g N_A_M1005_g 0.0328011f $X=3.205 $Y=0.85 $X2=3.635 $Y2=0.85
cc_262 N_B_c_314_n N_A_M1005_g 0.022402f $X=3.205 $Y=1.74 $X2=3.635 $Y2=0.85
cc_263 N_B_c_316_n N_A_M1005_g 0.00376362f $X=3.205 $Y=1.74 $X2=3.635 $Y2=0.85
cc_264 B N_A_M1005_g 9.23221e-19 $X=3.21 $Y=1.74 $X2=3.635 $Y2=0.85
cc_265 N_B_c_312_n N_A_c_412_n 0.0576612f $X=0.905 $Y=1.74 $X2=1.385 $Y2=2.11
cc_266 N_B_c_318_n N_A_c_412_n 7.99243e-19 $X=3.06 $Y=1.74 $X2=1.385 $Y2=2.11
cc_267 N_B_M1006_g N_A_c_413_n 0.125484f $X=3.265 $Y=3.235 $X2=3.685 $Y2=2.11
cc_268 N_B_M1001_g N_A_c_414_n 0.00286993f $X=0.965 $Y=3.235 $X2=1.385 $Y2=2.11
cc_269 N_B_c_318_n N_A_c_414_n 0.00428104f $X=3.06 $Y=1.74 $X2=1.385 $Y2=2.11
cc_270 N_B_M1006_g N_A_c_415_n 0.00278747f $X=3.265 $Y=3.235 $X2=3.685 $Y2=2.11
cc_271 N_B_M1001_g N_A_c_416_n 0.00405562f $X=0.965 $Y=3.235 $X2=1.53 $Y2=2.11
cc_272 N_B_c_318_n N_A_c_416_n 0.0263377f $X=3.06 $Y=1.74 $X2=1.53 $Y2=2.11
cc_273 N_B_M1006_g A 7.94897e-19 $X=3.265 $Y=3.235 $X2=3.685 $Y2=2.11
cc_274 N_B_M1006_g N_A_c_418_n 0.00633265f $X=3.265 $Y=3.235 $X2=3.54 $Y2=2.11
cc_275 N_B_c_314_n N_A_c_418_n 0.00210214f $X=3.205 $Y=1.74 $X2=3.54 $Y2=2.11
cc_276 N_B_c_316_n N_A_c_418_n 0.00225835f $X=3.205 $Y=1.74 $X2=3.54 $Y2=2.11
cc_277 N_B_c_318_n N_A_c_418_n 0.128931f $X=3.06 $Y=1.74 $X2=3.54 $Y2=2.11
cc_278 B N_A_c_418_n 0.0270107f $X=3.21 $Y=1.74 $X2=3.54 $Y2=2.11
cc_279 N_B_c_318_n N_A_208_521#_c_493_n 0.00725075f $X=3.06 $Y=1.74 $X2=1.885
+ $Y2=2.115
cc_280 N_B_c_318_n N_A_208_521#_c_495_n 0.00116539f $X=3.06 $Y=1.74 $X2=2.21
+ $Y2=1.32
cc_281 N_B_M1006_g N_A_208_521#_c_496_n 0.0358659f $X=3.265 $Y=3.235 $X2=2.76
+ $Y2=2.19
cc_282 N_B_c_318_n N_A_208_521#_c_496_n 0.00178159f $X=3.06 $Y=1.74 $X2=2.76
+ $Y2=2.19
cc_283 N_B_M1004_g N_A_208_521#_c_503_n 0.0265386f $X=3.205 $Y=0.85 $X2=2.775
+ $Y2=1.245
cc_284 N_B_M1001_g N_A_208_521#_c_529_n 0.00507079f $X=0.965 $Y=3.235 $X2=1.265
+ $Y2=2.53
cc_285 N_B_c_318_n N_A_208_521#_c_529_n 0.0051538f $X=3.06 $Y=1.74 $X2=1.265
+ $Y2=2.53
cc_286 N_B_c_315_n N_A_208_521#_c_513_n 0.00316158f $X=0.905 $Y=1.74 $X2=1.725
+ $Y2=2.445
cc_287 N_B_c_317_n N_A_208_521#_c_513_n 0.00129846f $X=1.05 $Y=1.74 $X2=1.725
+ $Y2=2.445
cc_288 N_B_c_318_n N_A_208_521#_c_513_n 0.0153226f $X=3.06 $Y=1.74 $X2=1.725
+ $Y2=2.445
cc_289 N_B_c_317_n N_A_208_521#_c_514_n 5.15761e-19 $X=1.05 $Y=1.74 $X2=1.725
+ $Y2=1.475
cc_290 N_B_c_318_n N_A_208_521#_c_514_n 0.00890945f $X=3.06 $Y=1.74 $X2=1.725
+ $Y2=1.475
cc_291 N_B_M1008_g S 4.14782e-19 $X=0.965 $Y=0.85 $X2=0.25 $Y2=1.905
cc_292 N_B_c_315_n S 0.00429487f $X=0.905 $Y=1.74 $X2=0.25 $Y2=1.905
cc_293 N_B_c_317_n S 0.0134542f $X=1.05 $Y=1.74 $X2=0.25 $Y2=1.905
cc_294 N_B_M1008_g N_S_c_611_n 7.50611e-19 $X=0.965 $Y=0.85 $X2=0.26 $Y2=0.995
cc_295 N_B_c_318_n N_CO_c_647_n 0.0136552f $X=3.06 $Y=1.74 $X2=2.137 $Y2=2.395
cc_296 N_A_M1010_g N_A_208_521#_c_493_n 0.00833244f $X=1.325 $Y=0.85 $X2=1.885
+ $Y2=2.115
cc_297 N_A_c_412_n N_A_208_521#_c_493_n 0.0147848f $X=1.385 $Y=2.11 $X2=1.885
+ $Y2=2.115
cc_298 N_A_c_418_n N_A_208_521#_c_493_n 0.00210973f $X=3.54 $Y=2.11 $X2=1.885
+ $Y2=2.115
cc_299 N_A_M1003_g N_A_208_521#_M1012_g 0.0405735f $X=1.395 $Y=3.235 $X2=1.885
+ $Y2=3.235
cc_300 N_A_c_418_n N_A_208_521#_c_496_n 0.0140186f $X=3.54 $Y=2.11 $X2=2.76
+ $Y2=2.19
cc_301 N_A_M1010_g N_A_208_521#_c_507_n 0.0166986f $X=1.325 $Y=0.85 $X2=1.825
+ $Y2=1.32
cc_302 N_A_c_418_n N_A_208_521#_c_508_n 0.00700381f $X=3.54 $Y=2.11 $X2=1.885
+ $Y2=2.19
cc_303 N_A_M1003_g N_A_208_521#_c_526_n 0.0147914f $X=1.395 $Y=3.235 $X2=1.64
+ $Y2=2.53
cc_304 N_A_c_412_n N_A_208_521#_c_526_n 0.00348735f $X=1.385 $Y=2.11 $X2=1.64
+ $Y2=2.53
cc_305 N_A_c_414_n N_A_208_521#_c_526_n 0.0111584f $X=1.385 $Y=2.11 $X2=1.64
+ $Y2=2.53
cc_306 N_A_c_416_n N_A_208_521#_c_526_n 0.00509311f $X=1.53 $Y=2.11 $X2=1.64
+ $Y2=2.53
cc_307 N_A_c_418_n N_A_208_521#_c_526_n 0.00467069f $X=3.54 $Y=2.11 $X2=1.64
+ $Y2=2.53
cc_308 N_A_c_412_n N_A_208_521#_c_529_n 7.25782e-19 $X=1.385 $Y=2.11 $X2=1.265
+ $Y2=2.53
cc_309 N_A_c_416_n N_A_208_521#_c_529_n 0.00124978f $X=1.53 $Y=2.11 $X2=1.265
+ $Y2=2.53
cc_310 N_A_M1010_g N_A_208_521#_c_510_n 0.00944415f $X=1.325 $Y=0.85 $X2=1.54
+ $Y2=0.755
cc_311 N_A_M1010_g N_A_208_521#_c_513_n 0.00392362f $X=1.325 $Y=0.85 $X2=1.725
+ $Y2=2.445
cc_312 N_A_M1003_g N_A_208_521#_c_513_n 0.00360042f $X=1.395 $Y=3.235 $X2=1.725
+ $Y2=2.445
cc_313 N_A_c_412_n N_A_208_521#_c_513_n 0.00193142f $X=1.385 $Y=2.11 $X2=1.725
+ $Y2=2.445
cc_314 N_A_c_414_n N_A_208_521#_c_513_n 0.0224238f $X=1.385 $Y=2.11 $X2=1.725
+ $Y2=2.445
cc_315 N_A_c_416_n N_A_208_521#_c_513_n 0.00168305f $X=1.53 $Y=2.11 $X2=1.725
+ $Y2=2.445
cc_316 N_A_c_418_n N_A_208_521#_c_513_n 0.0185059f $X=3.54 $Y=2.11 $X2=1.725
+ $Y2=2.445
cc_317 N_A_M1010_g N_A_208_521#_c_514_n 0.00736605f $X=1.325 $Y=0.85 $X2=1.725
+ $Y2=1.475
cc_318 N_A_c_412_n N_A_208_521#_c_514_n 0.00175929f $X=1.385 $Y=2.11 $X2=1.725
+ $Y2=1.475
cc_319 N_A_c_414_n N_A_208_521#_c_514_n 2.52704e-19 $X=1.385 $Y=2.11 $X2=1.725
+ $Y2=1.475
cc_320 N_A_c_418_n N_CO_c_646_n 0.00105312f $X=3.54 $Y=2.11 $X2=2.175 $Y2=2.48
cc_321 N_A_c_418_n N_CO_c_647_n 0.0133707f $X=3.54 $Y=2.11 $X2=2.137 $Y2=2.395
cc_322 N_A_c_418_n CO 0.0346374f $X=3.54 $Y=2.11 $X2=2.175 $Y2=2.48
cc_323 N_A_208_521#_c_510_n N_CO_c_640_n 0.013807f $X=1.54 $Y=0.755 $X2=2.07
+ $Y2=0.755
cc_324 N_A_208_521#_c_495_n N_CO_c_643_n 0.00425808f $X=2.21 $Y=1.32 $X2=2.175
+ $Y2=0.992
cc_325 N_A_208_521#_c_497_n N_CO_c_643_n 0.00712614f $X=2.285 $Y=1.245 $X2=2.175
+ $Y2=0.992
cc_326 N_A_208_521#_c_503_n N_CO_c_643_n 6.90609e-19 $X=2.775 $Y=1.245 $X2=2.175
+ $Y2=0.992
cc_327 N_A_208_521#_c_510_n N_CO_c_643_n 0.00752809f $X=1.54 $Y=0.755 $X2=2.175
+ $Y2=0.992
cc_328 N_A_208_521#_M1012_g N_CO_c_646_n 0.00839391f $X=1.885 $Y=3.235 $X2=2.175
+ $Y2=2.48
cc_329 N_A_208_521#_c_496_n N_CO_c_646_n 0.00140819f $X=2.76 $Y=2.19 $X2=2.175
+ $Y2=2.48
cc_330 N_A_208_521#_c_526_n N_CO_c_646_n 0.0104146f $X=1.64 $Y=2.53 $X2=2.175
+ $Y2=2.48
cc_331 N_A_208_521#_c_513_n N_CO_c_646_n 0.00298908f $X=1.725 $Y=2.445 $X2=2.175
+ $Y2=2.48
cc_332 N_A_208_521#_M1012_g N_CO_c_647_n 0.00273706f $X=1.885 $Y=3.235 $X2=2.137
+ $Y2=2.395
cc_333 N_A_208_521#_c_495_n N_CO_c_647_n 0.00814611f $X=2.21 $Y=1.32 $X2=2.137
+ $Y2=2.395
cc_334 N_A_208_521#_c_496_n N_CO_c_647_n 0.0137597f $X=2.76 $Y=2.19 $X2=2.137
+ $Y2=2.395
cc_335 N_A_208_521#_c_497_n N_CO_c_647_n 0.00629561f $X=2.285 $Y=1.245 $X2=2.137
+ $Y2=2.395
cc_336 N_A_208_521#_c_503_n N_CO_c_647_n 8.21103e-19 $X=2.775 $Y=1.245 $X2=2.137
+ $Y2=2.395
cc_337 N_A_208_521#_M1013_g N_CO_c_647_n 8.14457e-19 $X=2.835 $Y=3.235 $X2=2.137
+ $Y2=2.395
cc_338 N_A_208_521#_c_507_n N_CO_c_647_n 0.011021f $X=1.825 $Y=1.32 $X2=2.137
+ $Y2=2.395
cc_339 N_A_208_521#_c_509_n N_CO_c_647_n 0.00392207f $X=2.285 $Y=1.32 $X2=2.137
+ $Y2=2.395
cc_340 N_A_208_521#_c_510_n N_CO_c_647_n 0.00791989f $X=1.54 $Y=0.755 $X2=2.137
+ $Y2=2.395
cc_341 N_A_208_521#_c_513_n N_CO_c_647_n 0.0354244f $X=1.725 $Y=2.445 $X2=2.137
+ $Y2=2.395
cc_342 N_A_208_521#_c_514_n N_CO_c_647_n 0.0222722f $X=1.725 $Y=1.475 $X2=2.137
+ $Y2=2.395
cc_343 N_A_208_521#_M1012_g CO 7.58429e-19 $X=1.885 $Y=3.235 $X2=2.175 $Y2=2.48
cc_344 N_A_208_521#_c_496_n CO 0.0027071f $X=2.76 $Y=2.19 $X2=2.175 $Y2=2.48
cc_345 N_A_208_521#_c_526_n CO 0.00111652f $X=1.64 $Y=2.53 $X2=2.175 $Y2=2.48
cc_346 N_A_208_521#_c_513_n CO 0.0012063f $X=1.725 $Y=2.445 $X2=2.175 $Y2=2.48
