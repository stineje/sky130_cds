* File: sky130_osu_sc_18T_hs__or2_l.pxi.spice
* Created: Fri Nov 12 13:52:56 2021
* 
x_PM_SKY130_OSU_SC_18T_HS__OR2_L%GND N_GND_M1002_s N_GND_M1000_d N_GND_M1002_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_HS__OR2_L%GND
x_PM_SKY130_OSU_SC_18T_HS__OR2_L%VDD N_VDD_M1003_d N_VDD_M1005_b N_VDD_c_37_p
+ N_VDD_c_43_p N_VDD_c_49_p VDD N_VDD_c_38_p PM_SKY130_OSU_SC_18T_HS__OR2_L%VDD
x_PM_SKY130_OSU_SC_18T_HS__OR2_L%B N_B_M1002_g N_B_M1005_g N_B_c_66_n N_B_c_67_n
+ B PM_SKY130_OSU_SC_18T_HS__OR2_L%B
x_PM_SKY130_OSU_SC_18T_HS__OR2_L%A N_A_M1000_g N_A_M1003_g N_A_c_95_n N_A_c_96_n
+ A PM_SKY130_OSU_SC_18T_HS__OR2_L%A
x_PM_SKY130_OSU_SC_18T_HS__OR2_L%A_27_817# N_A_27_817#_M1002_d
+ N_A_27_817#_M1005_s N_A_27_817#_M1001_g N_A_27_817#_M1004_g
+ N_A_27_817#_c_136_n N_A_27_817#_c_137_n N_A_27_817#_c_138_n
+ N_A_27_817#_c_150_n N_A_27_817#_c_153_n N_A_27_817#_c_154_n
+ N_A_27_817#_c_139_n N_A_27_817#_c_140_n N_A_27_817#_c_143_n
+ N_A_27_817#_c_144_n PM_SKY130_OSU_SC_18T_HS__OR2_L%A_27_817#
x_PM_SKY130_OSU_SC_18T_HS__OR2_L%Y N_Y_M1001_d N_Y_M1004_d N_Y_c_203_n
+ N_Y_c_206_n Y N_Y_c_208_n N_Y_c_209_n PM_SKY130_OSU_SC_18T_HS__OR2_L%Y
cc_1 N_GND_M1002_b N_B_M1002_g 0.105092f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_B_M1002_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_B_M1002_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.945
cc_4 N_GND_c_4_p N_B_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.945
cc_5 N_GND_M1002_b N_B_M1005_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=5.085
cc_6 N_GND_M1002_b N_B_c_66_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.675
cc_7 N_GND_M1002_b N_B_c_67_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.675
cc_8 N_GND_M1002_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.96
cc_9 N_GND_M1002_b N_A_M1000_g 0.0580646f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.945
cc_10 N_GND_c_3_p N_A_M1000_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.945
cc_11 N_GND_c_11_p N_A_M1000_g 0.00354579f $X=1.12 $Y=0.825 $X2=0.905 $Y2=0.945
cc_12 N_GND_c_4_p N_A_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=0.945
cc_13 N_GND_M1002_b N_A_M1003_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=5.085
cc_14 N_GND_M1002_b N_A_c_95_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.385
cc_15 N_GND_M1002_b N_A_c_96_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.385
cc_16 N_GND_M1002_b N_A_27_817#_M1001_g 0.0449913f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.945
cc_17 N_GND_c_11_p N_A_27_817#_M1001_g 0.00354579f $X=1.12 $Y=0.825 $X2=1.335
+ $Y2=0.945
cc_18 N_GND_c_18_p N_A_27_817#_M1001_g 0.00606474f $X=1.12 $Y=0.152 $X2=1.335
+ $Y2=0.945
cc_19 N_GND_c_4_p N_A_27_817#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=0.945
cc_20 N_GND_M1002_b N_A_27_817#_c_136_n 0.0364586f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.1
cc_21 N_GND_M1002_b N_A_27_817#_c_137_n 0.0466273f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.81
cc_22 N_GND_M1002_b N_A_27_817#_c_138_n 0.0076653f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.96
cc_23 N_GND_M1002_b N_A_27_817#_c_139_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.545
cc_24 N_GND_M1002_b N_A_27_817#_c_140_n 0.0134398f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.825
cc_25 N_GND_c_3_p N_A_27_817#_c_140_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.825
cc_26 N_GND_c_4_p N_A_27_817#_c_140_n 0.00475776f $X=1.02 $Y=0.19 $X2=0.69
+ $Y2=0.825
cc_27 N_GND_M1002_b N_A_27_817#_c_143_n 0.0235867f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_28 N_GND_M1002_b N_A_27_817#_c_144_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.935
cc_29 N_GND_M1002_b N_Y_c_203_n 0.0115904f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_30 N_GND_c_18_p N_Y_c_203_n 0.00757793f $X=1.12 $Y=0.152 $X2=1.55 $Y2=0.825
cc_31 N_GND_c_4_p N_Y_c_203_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.825
cc_32 N_GND_M1002_b N_Y_c_206_n 0.016457f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_33 N_GND_M1002_b Y 0.039938f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_34 N_GND_M1002_b N_Y_c_208_n 0.0157042f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.48
cc_35 N_GND_M1002_b N_Y_c_209_n 0.0141689f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_36 N_VDD_M1005_b N_B_M1005_g 0.0918303f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_37 N_VDD_c_37_p N_B_M1005_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=5.085
cc_38 N_VDD_c_38_p N_B_M1005_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=5.085
cc_39 N_VDD_M1005_b N_B_c_67_n 0.00375034f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.675
cc_40 N_VDD_M1005_b B 0.0108395f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.96
cc_41 N_VDD_M1005_b N_A_M1003_g 0.0703255f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=5.085
cc_42 N_VDD_c_37_p N_A_M1003_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=5.085
cc_43 N_VDD_c_43_p N_A_M1003_g 0.00354579f $X=1.12 $Y=4.815 $X2=0.905 $Y2=5.085
cc_44 N_VDD_c_38_p N_A_M1003_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.905 $Y2=5.085
cc_45 N_VDD_M1005_b N_A_c_96_n 0.00479112f $X=-0.045 $Y=2.905 $X2=0.95 $Y2=2.385
cc_46 N_VDD_M1005_b A 0.0200864f $X=-0.045 $Y=2.905 $X2=0.95 $Y2=3.33
cc_47 N_VDD_M1005_b N_A_27_817#_M1004_g 0.0777475f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=5.085
cc_48 N_VDD_c_43_p N_A_27_817#_M1004_g 0.00354579f $X=1.12 $Y=4.815 $X2=1.335
+ $Y2=5.085
cc_49 N_VDD_c_49_p N_A_27_817#_M1004_g 0.00606474f $X=1.12 $Y=6.507 $X2=1.335
+ $Y2=5.085
cc_50 N_VDD_c_38_p N_A_27_817#_M1004_g 0.00468827f $X=1.02 $Y=6.47 $X2=1.335
+ $Y2=5.085
cc_51 N_VDD_M1005_b N_A_27_817#_c_138_n 0.00525234f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.96
cc_52 N_VDD_M1005_b N_A_27_817#_c_150_n 0.0190556f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.815
cc_53 N_VDD_c_37_p N_A_27_817#_c_150_n 0.00736239f $X=1.035 $Y=6.507 $X2=0.26
+ $Y2=4.815
cc_54 N_VDD_c_38_p N_A_27_817#_c_150_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26
+ $Y2=4.815
cc_55 N_VDD_M1005_b N_A_27_817#_c_153_n 0.0103569f $X=-0.045 $Y=2.905 $X2=0.525
+ $Y2=3.63
cc_56 N_VDD_M1005_b N_A_27_817#_c_154_n 0.00927559f $X=-0.045 $Y=2.905 $X2=0.345
+ $Y2=3.63
cc_57 N_VDD_M1005_b N_A_27_817#_c_139_n 0.00377157f $X=-0.045 $Y=2.905 $X2=0.61
+ $Y2=3.545
cc_58 N_VDD_M1005_b N_Y_c_206_n 0.0591925f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.59
cc_59 N_VDD_c_49_p N_Y_c_206_n 0.00757793f $X=1.12 $Y=6.507 $X2=1.55 $Y2=2.59
cc_60 N_VDD_c_38_p N_Y_c_206_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.55 $Y2=2.59
cc_61 N_B_M1002_g N_A_M1000_g 0.052095f $X=0.475 $Y=0.945 $X2=0.905 $Y2=0.945
cc_62 N_B_c_66_n N_A_M1003_g 0.15786f $X=0.475 $Y=2.675 $X2=0.905 $Y2=5.085
cc_63 N_B_M1002_g N_A_c_95_n 0.0148656f $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.385
cc_64 N_B_M1002_g N_A_c_96_n 0.00121111f $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.385
cc_65 N_B_M1005_g N_A_27_817#_c_150_n 0.0256225f $X=0.475 $Y=5.085 $X2=0.26
+ $Y2=4.815
cc_66 N_B_M1005_g N_A_27_817#_c_153_n 0.0162328f $X=0.475 $Y=5.085 $X2=0.525
+ $Y2=3.63
cc_67 B N_A_27_817#_c_153_n 0.00520961f $X=0.27 $Y=2.96 $X2=0.525 $Y2=3.63
cc_68 N_B_c_67_n N_A_27_817#_c_154_n 0.00389696f $X=0.27 $Y=2.675 $X2=0.345
+ $Y2=3.63
cc_69 B N_A_27_817#_c_154_n 0.00433184f $X=0.27 $Y=2.96 $X2=0.345 $Y2=3.63
cc_70 N_B_M1002_g N_A_27_817#_c_139_n 0.0231435f $X=0.475 $Y=0.945 $X2=0.61
+ $Y2=3.545
cc_71 N_B_M1005_g N_A_27_817#_c_139_n 0.026563f $X=0.475 $Y=5.085 $X2=0.61
+ $Y2=3.545
cc_72 N_B_c_66_n N_A_27_817#_c_139_n 0.00764878f $X=0.475 $Y=2.675 $X2=0.61
+ $Y2=3.545
cc_73 N_B_c_67_n N_A_27_817#_c_139_n 0.0350086f $X=0.27 $Y=2.675 $X2=0.61
+ $Y2=3.545
cc_74 B N_A_27_817#_c_139_n 0.00758489f $X=0.27 $Y=2.96 $X2=0.61 $Y2=3.545
cc_75 N_B_M1002_g N_A_27_817#_c_140_n 0.0142017f $X=0.475 $Y=0.945 $X2=0.69
+ $Y2=0.825
cc_76 N_B_M1002_g N_A_27_817#_c_144_n 0.0113001f $X=0.475 $Y=0.945 $X2=0.65
+ $Y2=1.935
cc_77 N_A_M1000_g N_A_27_817#_M1001_g 0.044975f $X=0.905 $Y=0.945 $X2=1.335
+ $Y2=0.945
cc_78 A N_A_27_817#_M1004_g 0.00374181f $X=0.95 $Y=3.33 $X2=1.335 $Y2=5.085
cc_79 N_A_M1000_g N_A_27_817#_c_136_n 0.0119161f $X=0.905 $Y=0.945 $X2=1.37
+ $Y2=2.1
cc_80 N_A_M1003_g N_A_27_817#_c_137_n 0.00914307f $X=0.905 $Y=5.085 $X2=1.352
+ $Y2=2.81
cc_81 N_A_c_95_n N_A_27_817#_c_137_n 0.0204279f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.81
cc_82 N_A_c_96_n N_A_27_817#_c_137_n 0.00375034f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.81
cc_83 N_A_M1003_g N_A_27_817#_c_138_n 0.0855856f $X=0.905 $Y=5.085 $X2=1.352
+ $Y2=2.96
cc_84 N_A_c_96_n N_A_27_817#_c_138_n 0.00434324f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.96
cc_85 N_A_M1003_g N_A_27_817#_c_153_n 0.00457566f $X=0.905 $Y=5.085 $X2=0.525
+ $Y2=3.63
cc_86 N_A_M1000_g N_A_27_817#_c_139_n 0.00429604f $X=0.905 $Y=0.945 $X2=0.61
+ $Y2=3.545
cc_87 N_A_M1003_g N_A_27_817#_c_139_n 0.00776428f $X=0.905 $Y=5.085 $X2=0.61
+ $Y2=3.545
cc_88 N_A_c_95_n N_A_27_817#_c_139_n 0.0021255f $X=0.95 $Y=2.385 $X2=0.61
+ $Y2=3.545
cc_89 N_A_c_96_n N_A_27_817#_c_139_n 0.0825894f $X=0.95 $Y=2.385 $X2=0.61
+ $Y2=3.545
cc_90 A N_A_27_817#_c_139_n 0.00866797f $X=0.95 $Y=3.33 $X2=0.61 $Y2=3.545
cc_91 N_A_M1000_g N_A_27_817#_c_140_n 0.0142017f $X=0.905 $Y=0.945 $X2=0.69
+ $Y2=0.825
cc_92 N_A_M1000_g N_A_27_817#_c_143_n 0.0163305f $X=0.905 $Y=0.945 $X2=1.43
+ $Y2=1.935
cc_93 N_A_c_95_n N_A_27_817#_c_143_n 0.00276813f $X=0.95 $Y=2.385 $X2=1.43
+ $Y2=1.935
cc_94 N_A_c_96_n N_A_27_817#_c_143_n 0.0114342f $X=0.95 $Y=2.385 $X2=1.43
+ $Y2=1.935
cc_95 N_A_c_96_n N_Y_c_206_n 0.0300473f $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_96 A N_Y_c_206_n 0.00659455f $X=0.95 $Y=3.33 $X2=1.55 $Y2=2.59
cc_97 N_A_M1000_g Y 6.73508e-19 $X=0.905 $Y=0.945 $X2=1.555 $Y2=2.22
cc_98 N_A_c_96_n Y 0.00825539f $X=0.95 $Y=2.385 $X2=1.555 $Y2=2.22
cc_99 N_A_M1000_g N_Y_c_208_n 0.00102215f $X=0.905 $Y=0.945 $X2=1.55 $Y2=1.48
cc_100 N_A_c_95_n N_Y_c_209_n 3.65268e-19 $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_101 N_A_c_96_n N_Y_c_209_n 0.00535705f $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_102 N_A_27_817#_M1001_g N_Y_c_203_n 0.0152627f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=0.825
cc_103 N_A_27_817#_c_136_n N_Y_c_203_n 0.00168f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=0.825
cc_104 N_A_27_817#_c_143_n N_Y_c_203_n 0.00530006f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_105 N_A_27_817#_M1004_g N_Y_c_206_n 0.0488265f $X=1.335 $Y=5.085 $X2=1.55
+ $Y2=2.59
cc_106 N_A_27_817#_c_136_n N_Y_c_206_n 0.00125776f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_107 N_A_27_817#_c_137_n N_Y_c_206_n 0.0115869f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_108 N_A_27_817#_c_143_n N_Y_c_206_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_109 N_A_27_817#_M1001_g Y 0.00406656f $X=1.335 $Y=0.945 $X2=1.555 $Y2=2.22
cc_110 N_A_27_817#_c_136_n Y 0.00704613f $X=1.37 $Y=2.1 $X2=1.555 $Y2=2.22
cc_111 N_A_27_817#_c_137_n Y 0.00892438f $X=1.352 $Y=2.81 $X2=1.555 $Y2=2.22
cc_112 N_A_27_817#_c_143_n Y 0.0151477f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_113 N_A_27_817#_M1001_g N_Y_c_208_n 0.00715333f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=1.48
cc_114 N_A_27_817#_c_136_n N_Y_c_208_n 0.00154864f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=1.48
cc_115 N_A_27_817#_c_143_n N_Y_c_208_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.48
cc_116 N_A_27_817#_c_136_n N_Y_c_209_n 4.58687e-19 $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_117 N_A_27_817#_c_137_n N_Y_c_209_n 0.00721849f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_118 N_A_27_817#_c_143_n N_Y_c_209_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
