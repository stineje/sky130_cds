* File: sky130_osu_sc_12T_hs__inv_3.pxi.spice
* Created: Fri Nov 12 15:10:53 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__INV_3%GND N_GND_M1001_d N_GND_M1002_d N_GND_M1001_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p N_GND_c_17_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_HS__INV_3%GND
x_PM_SKY130_OSU_SC_12T_HS__INV_3%VDD N_VDD_M1000_s N_VDD_M1004_s N_VDD_M1000_b
+ N_VDD_c_50_p N_VDD_c_51_p N_VDD_c_56_p N_VDD_c_62_p VDD N_VDD_c_52_p
+ PM_SKY130_OSU_SC_12T_HS__INV_3%VDD
x_PM_SKY130_OSU_SC_12T_HS__INV_3%A N_A_c_82_n N_A_M1001_g N_A_c_86_n N_A_c_109_n
+ N_A_M1000_g N_A_c_87_n N_A_c_88_n N_A_c_89_n N_A_M1002_g N_A_c_114_n
+ N_A_M1004_g N_A_c_93_n N_A_c_95_n N_A_c_96_n N_A_M1003_g N_A_c_120_n
+ N_A_M1005_g N_A_c_100_n N_A_c_101_n N_A_c_102_n N_A_c_103_n N_A_c_104_n
+ N_A_c_105_n N_A_c_106_n N_A_c_107_n N_A_c_108_n A
+ PM_SKY130_OSU_SC_12T_HS__INV_3%A
x_PM_SKY130_OSU_SC_12T_HS__INV_3%Y N_Y_M1001_s N_Y_M1003_s N_Y_M1000_d
+ N_Y_M1005_d N_Y_c_178_n N_Y_c_199_n N_Y_c_182_n N_Y_c_186_n N_Y_c_187_n
+ N_Y_c_205_n Y N_Y_c_191_n N_Y_c_206_n N_Y_c_195_n N_Y_c_198_n
+ PM_SKY130_OSU_SC_12T_HS__INV_3%Y
cc_1 N_GND_M1001_b N_A_c_82_n 0.018528f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.22
cc_2 N_GND_c_2_p N_A_c_82_n 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=1.22
cc_3 N_GND_c_3_p N_A_c_82_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.22
cc_4 N_GND_c_4_p N_A_c_82_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.22
cc_5 N_GND_M1001_b N_A_c_86_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.33
cc_6 N_GND_M1001_b N_A_c_87_n 0.0162043f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.295
cc_7 N_GND_M1001_b N_A_c_88_n 0.0114349f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.405
cc_8 N_GND_M1001_b N_A_c_89_n 0.0152079f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.22
cc_9 N_GND_c_3_p N_A_c_89_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.22
cc_10 N_GND_c_10_p N_A_c_89_n 0.00311745f $X=1.12 $Y=0.755 $X2=0.905 $Y2=1.22
cc_11 N_GND_c_4_p N_A_c_89_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=1.22
cc_12 N_GND_M1001_b N_A_c_93_n 0.037872f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.295
cc_13 N_GND_c_10_p N_A_c_93_n 0.00283047f $X=1.12 $Y=0.755 $X2=1.26 $Y2=1.295
cc_14 N_GND_M1001_b N_A_c_95_n 0.0305509f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.405
cc_15 N_GND_M1001_b N_A_c_96_n 0.0205268f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.22
cc_16 N_GND_c_10_p N_A_c_96_n 0.00311745f $X=1.12 $Y=0.755 $X2=1.335 $Y2=1.22
cc_17 N_GND_c_17_p N_A_c_96_n 0.00606474f $X=1.12 $Y=0.152 $X2=1.335 $Y2=1.22
cc_18 N_GND_c_4_p N_A_c_96_n 0.00468827f $X=1.02 $Y=0.19 $X2=1.335 $Y2=1.22
cc_19 N_GND_M1001_b N_A_c_100_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.295
cc_20 N_GND_M1001_b N_A_c_101_n 0.0348407f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_21 N_GND_M1001_b N_A_c_102_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.66
cc_22 N_GND_M1001_b N_A_c_103_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.405
cc_23 N_GND_M1001_b N_A_c_104_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.295
cc_24 N_GND_M1001_b N_A_c_105_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.405
cc_25 N_GND_M1001_b N_A_c_106_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.85
cc_26 N_GND_M1001_b N_A_c_107_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.825
cc_27 N_GND_M1001_b N_A_c_108_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_28 N_GND_M1001_b N_Y_c_178_n 0.00154299f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.755
cc_29 N_GND_c_3_p N_Y_c_178_n 0.00740081f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.755
cc_30 N_GND_c_10_p N_Y_c_178_n 8.14297e-19 $X=1.12 $Y=0.755 $X2=0.69 $Y2=0.755
cc_31 N_GND_c_4_p N_Y_c_178_n 0.0047139f $X=1.02 $Y=0.19 $X2=0.69 $Y2=0.755
cc_32 N_GND_M1001_b N_Y_c_182_n 0.00155228f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_33 N_GND_c_10_p N_Y_c_182_n 8.14297e-19 $X=1.12 $Y=0.755 $X2=1.55 $Y2=0.755
cc_34 N_GND_c_17_p N_Y_c_182_n 0.0074222f $X=1.12 $Y=0.152 $X2=1.55 $Y2=0.755
cc_35 N_GND_c_4_p N_Y_c_182_n 0.00471849f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.755
cc_36 N_GND_M1001_b N_Y_c_186_n 0.00312976f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.48
cc_37 N_GND_c_2_p N_Y_c_187_n 0.00134236f $X=0.26 $Y=0.755 $X2=0.69 $Y2=1.115
cc_38 N_GND_c_3_p N_Y_c_187_n 0.00245319f $X=1.035 $Y=0.152 $X2=0.69 $Y2=1.115
cc_39 N_GND_c_10_p N_Y_c_187_n 7.53951e-19 $X=1.12 $Y=0.755 $X2=0.69 $Y2=1.115
cc_40 N_GND_M1001_b Y 0.0453816f $X=-0.045 $Y=0 $X2=0.76 $Y2=1.72
cc_41 N_GND_M1002_d N_Y_c_191_n 0.0100144f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1
cc_42 N_GND_c_3_p N_Y_c_191_n 0.0028844f $X=1.035 $Y=0.152 $X2=1.405 $Y2=1
cc_43 N_GND_c_10_p N_Y_c_191_n 0.0142303f $X=1.12 $Y=0.755 $X2=1.405 $Y2=1
cc_44 N_GND_c_17_p N_Y_c_191_n 0.0028844f $X=1.12 $Y=0.152 $X2=1.405 $Y2=1
cc_45 N_GND_M1001_b N_Y_c_195_n 0.0101598f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.115
cc_46 N_GND_c_10_p N_Y_c_195_n 7.53951e-19 $X=1.12 $Y=0.755 $X2=1.55 $Y2=1.115
cc_47 N_GND_c_17_p N_Y_c_195_n 0.00253787f $X=1.12 $Y=0.152 $X2=1.55 $Y2=1.115
cc_48 N_GND_M1001_b N_Y_c_198_n 0.0945652f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.365
cc_49 N_VDD_M1000_b N_A_c_109_n 0.0181616f $X=-0.045 $Y=2.425 $X2=0.475 $Y2=2.48
cc_50 N_VDD_c_50_p N_A_c_109_n 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=2.48
cc_51 N_VDD_c_51_p N_A_c_109_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=2.48
cc_52 N_VDD_c_52_p N_A_c_109_n 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=2.48
cc_53 N_VDD_M1000_b N_A_c_88_n 0.00448664f $X=-0.045 $Y=2.425 $X2=0.83 $Y2=2.405
cc_54 N_VDD_M1000_b N_A_c_114_n 0.0159283f $X=-0.045 $Y=2.425 $X2=0.905 $Y2=2.48
cc_55 N_VDD_c_51_p N_A_c_114_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=2.48
cc_56 N_VDD_c_56_p N_A_c_114_n 0.00337744f $X=1.12 $Y=2.955 $X2=0.905 $Y2=2.48
cc_57 N_VDD_c_52_p N_A_c_114_n 0.00468827f $X=1.02 $Y=4.25 $X2=0.905 $Y2=2.48
cc_58 N_VDD_M1000_b N_A_c_95_n 0.00774816f $X=-0.045 $Y=2.425 $X2=1.26 $Y2=2.405
cc_59 N_VDD_c_56_p N_A_c_95_n 0.00341318f $X=1.12 $Y=2.955 $X2=1.26 $Y2=2.405
cc_60 N_VDD_M1000_b N_A_c_120_n 0.0221472f $X=-0.045 $Y=2.425 $X2=1.335 $Y2=2.48
cc_61 N_VDD_c_56_p N_A_c_120_n 0.00337744f $X=1.12 $Y=2.955 $X2=1.335 $Y2=2.48
cc_62 N_VDD_c_62_p N_A_c_120_n 0.00606474f $X=1.12 $Y=4.287 $X2=1.335 $Y2=2.48
cc_63 N_VDD_c_52_p N_A_c_120_n 0.00468827f $X=1.02 $Y=4.25 $X2=1.335 $Y2=2.48
cc_64 N_VDD_M1000_b N_A_c_103_n 0.00244521f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.405
cc_65 N_VDD_M1000_b N_A_c_105_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.405
cc_66 N_VDD_M1000_s N_A_c_106_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.85
cc_67 N_VDD_M1000_b N_A_c_106_n 0.00618364f $X=-0.045 $Y=2.425 $X2=0.32 $Y2=2.85
cc_68 N_VDD_c_50_p N_A_c_106_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_69 N_VDD_M1000_s A 0.0162774f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.845
cc_70 N_VDD_c_50_p A 0.00522047f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.845
cc_71 N_VDD_c_56_p A 9.09141e-19 $X=1.12 $Y=2.955 $X2=0.32 $Y2=2.845
cc_72 N_VDD_M1000_b N_Y_c_199_n 0.00361433f $X=-0.045 $Y=2.425 $X2=0.69 $Y2=2.48
cc_73 N_VDD_c_51_p N_Y_c_199_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69 $Y2=2.48
cc_74 N_VDD_c_52_p N_Y_c_199_n 0.00475776f $X=1.02 $Y=4.25 $X2=0.69 $Y2=2.48
cc_75 N_VDD_M1000_b N_Y_c_186_n 0.00745764f $X=-0.045 $Y=2.425 $X2=1.55 $Y2=2.48
cc_76 N_VDD_c_62_p N_Y_c_186_n 0.00757793f $X=1.12 $Y=4.287 $X2=1.55 $Y2=2.48
cc_77 N_VDD_c_52_p N_Y_c_186_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.55 $Y2=2.48
cc_78 N_VDD_M1000_b N_Y_c_205_n 0.00248543f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=2.365
cc_79 N_VDD_M1000_b N_Y_c_206_n 0.00520877f $X=-0.045 $Y=2.425 $X2=1.405
+ $Y2=2.48
cc_80 N_VDD_c_56_p N_Y_c_206_n 0.0090257f $X=1.12 $Y=2.955 $X2=1.405 $Y2=2.48
cc_81 N_VDD_M1000_b N_Y_c_198_n 0.0111011f $X=-0.045 $Y=2.425 $X2=1.55 $Y2=2.365
cc_82 A N_Y_M1000_d 0.00250716f $X=0.32 $Y=2.845 $X2=0.55 $Y2=2.605
cc_83 N_A_c_82_n N_Y_c_178_n 0.00182852f $X=0.475 $Y=1.22 $X2=0.69 $Y2=0.755
cc_84 N_A_c_87_n N_Y_c_178_n 0.00251439f $X=0.83 $Y=1.295 $X2=0.69 $Y2=0.755
cc_85 N_A_c_89_n N_Y_c_178_n 0.00182852f $X=0.905 $Y=1.22 $X2=0.69 $Y2=0.755
cc_86 N_A_c_108_n N_Y_c_178_n 0.00109947f $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.755
cc_87 N_A_c_109_n N_Y_c_199_n 0.00183112f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.48
cc_88 N_A_c_88_n N_Y_c_199_n 0.00864247f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.48
cc_89 N_A_c_114_n N_Y_c_199_n 0.00335296f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.48
cc_90 N_A_c_101_n N_Y_c_199_n 2.38128e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_91 N_A_c_106_n N_Y_c_199_n 0.0226156f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_92 N_A_c_108_n N_Y_c_199_n 0.00165526f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_93 A N_Y_c_199_n 0.00938699f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.48
cc_94 N_A_c_96_n N_Y_c_182_n 0.00356431f $X=1.335 $Y=1.22 $X2=1.55 $Y2=0.755
cc_95 N_A_c_95_n N_Y_c_186_n 0.0109268f $X=1.26 $Y=2.405 $X2=1.55 $Y2=2.48
cc_96 N_A_c_82_n N_Y_c_187_n 0.00880716f $X=0.475 $Y=1.22 $X2=0.69 $Y2=1.115
cc_97 N_A_c_89_n N_Y_c_187_n 0.00198464f $X=0.905 $Y=1.22 $X2=0.69 $Y2=1.115
cc_98 N_A_c_101_n N_Y_c_187_n 6.32153e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=1.115
cc_99 N_A_c_109_n N_Y_c_205_n 0.00169643f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.365
cc_100 N_A_c_88_n N_Y_c_205_n 0.00259868f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.365
cc_101 N_A_c_114_n N_Y_c_205_n 0.00144225f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.365
cc_102 N_A_c_101_n N_Y_c_205_n 2.98633e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.365
cc_103 N_A_c_103_n N_Y_c_205_n 0.00102602f $X=0.475 $Y=2.405 $X2=0.69 $Y2=2.365
cc_104 N_A_c_105_n N_Y_c_205_n 0.00150284f $X=0.905 $Y=2.405 $X2=0.69 $Y2=2.365
cc_105 N_A_c_106_n N_Y_c_205_n 0.0071561f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.365
cc_106 N_A_c_108_n N_Y_c_205_n 0.00173027f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.365
cc_107 A N_Y_c_205_n 0.00805971f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.365
cc_108 N_A_c_82_n Y 0.00150089f $X=0.475 $Y=1.22 $X2=0.76 $Y2=1.72
cc_109 N_A_c_86_n Y 0.00792324f $X=0.475 $Y=2.33 $X2=0.76 $Y2=1.72
cc_110 N_A_c_87_n Y 0.0163225f $X=0.83 $Y=1.295 $X2=0.76 $Y2=1.72
cc_111 N_A_c_88_n Y 0.0038871f $X=0.83 $Y=2.405 $X2=0.76 $Y2=1.72
cc_112 N_A_c_89_n Y 0.00150089f $X=0.905 $Y=1.22 $X2=0.76 $Y2=1.72
cc_113 N_A_c_101_n Y 0.00610708f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_114 N_A_c_102_n Y 0.00675469f $X=0.535 $Y=1.66 $X2=0.76 $Y2=1.72
cc_115 N_A_c_106_n Y 0.0182346f $X=0.32 $Y=2.85 $X2=0.76 $Y2=1.72
cc_116 N_A_c_108_n Y 0.0178517f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_117 N_A_c_89_n N_Y_c_191_n 0.00871678f $X=0.905 $Y=1.22 $X2=1.405 $Y2=1
cc_118 N_A_c_93_n N_Y_c_191_n 0.0022289f $X=1.26 $Y=1.295 $X2=1.405 $Y2=1
cc_119 N_A_c_96_n N_Y_c_191_n 0.00869047f $X=1.335 $Y=1.22 $X2=1.405 $Y2=1
cc_120 N_A_c_114_n N_Y_c_206_n 0.0069535f $X=0.905 $Y=2.48 $X2=1.405 $Y2=2.48
cc_121 N_A_c_95_n N_Y_c_206_n 0.0176406f $X=1.26 $Y=2.405 $X2=1.405 $Y2=2.48
cc_122 N_A_c_120_n N_Y_c_206_n 0.00693713f $X=1.335 $Y=2.48 $X2=1.405 $Y2=2.48
cc_123 N_A_c_105_n N_Y_c_206_n 0.00560085f $X=0.905 $Y=2.405 $X2=1.405 $Y2=2.48
cc_124 N_A_c_96_n N_Y_c_195_n 0.00300301f $X=1.335 $Y=1.22 $X2=1.55 $Y2=1.115
cc_125 N_A_c_95_n N_Y_c_198_n 0.00397242f $X=1.26 $Y=2.405 $X2=1.55 $Y2=2.365
cc_126 N_A_c_96_n N_Y_c_198_n 0.00700756f $X=1.335 $Y=1.22 $X2=1.55 $Y2=2.365
cc_127 N_A_c_120_n N_Y_c_198_n 0.00214586f $X=1.335 $Y=2.48 $X2=1.55 $Y2=2.365
