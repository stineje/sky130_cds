* File: sky130_osu_sc_15T_hs__or2_1.spice
* Created: Fri Nov 12 14:32:31 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__or2_1.pex.spice"
.subckt sky130_osu_sc_15T_hs__or2_1  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1004 N_A_27_565#_M1004_d N_B_M1004_g N_GND_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_GND_M1000_d N_A_M1000_g N_A_27_565#_M1004_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_Y_M1001_d N_A_27_565#_M1001_g N_GND_M1000_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 A_110_565# N_B_M1005_g N_A_27_565#_M1005_s N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=8.3528 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1002 N_VDD_M1002_d N_A_M1002_g A_110_565# N_VDD_M1005_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=8.3528 M=1 R=13.3333 SA=75000.6
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1003 N_Y_M1003_d N_A_27_565#_M1003_g N_VDD_M1002_d N_VDD_M1005_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1005_b NWDIODE A=5.64925 P=9.73
pX7_noxref noxref_8 B B PROBETYPE=1
pX8_noxref noxref_9 A A PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__or2_1.pxi.spice"
*
.ends
*
*
