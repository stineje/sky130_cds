* File: sky130_osu_sc_12T_ls__oai22_l.pex.spice
* Created: Fri Nov 12 15:39:20 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%GND 1 23 25 33 48 50
r44 48 50 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r45 35 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r46 31 44 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r47 31 33 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r48 25 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r49 23 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r50 23 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r51 23 35 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r52 23 25 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r53 1 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%VDD 1 2 21 25 27 36 45 49
r22 45 49 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.7 $Y2=4.287
r23 41 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r24 34 43 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.91 $Y=4.135
+ $X2=1.91 $Y2=4.287
r25 34 36 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.91 $Y=4.135
+ $X2=1.91 $Y2=3.35
r26 32 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=4.25 $X2=1.7
+ $Y2=4.25
r27 30 32 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r28 28 41 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r29 28 30 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r30 27 43 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=4.287
+ $X2=1.91 $Y2=4.287
r31 27 32 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=4.287
+ $X2=1.7 $Y2=4.287
r32 23 41 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r33 23 25 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.35
r34 21 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r35 21 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r36 21 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r37 2 36 300 $w=1.7e-07 $l=8.11988e-07 $layer=licon1_PDIFF $count=2 $X=1.77
+ $Y=2.605 $X2=1.91 $Y2=3.35
r38 1 25 300 $w=1.7e-07 $l=8.05078e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.35
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%A0 2 5 7 9 13 18 24
r28 18 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.345 $Y=2.11
+ $X2=0.345 $Y2=2.11
r29 18 21 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.345 $Y=2.11
+ $X2=0.345 $Y2=2.275
r30 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.345
+ $Y=2.275 $X2=0.345 $Y2=2.275
r31 11 13 62.1936 $w=1.55e-07 $l=1.3e-07 $layer=POLY_cond $X=0.345 $Y=1.307
+ $X2=0.475 $Y2=1.307
r32 7 16 39.3623 $w=2.99e-07 $l=2.1225e-07 $layer=POLY_cond $X=0.475 $Y=2.445
+ $X2=0.38 $Y2=2.275
r33 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=2.445
+ $X2=0.475 $Y2=3.235
r34 3 13 3.61756 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=0.475 $Y=1.23
+ $X2=0.475 $Y2=1.307
r35 3 5 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=1.23
+ $X2=0.475 $Y2=0.835
r36 2 16 39.5263 $w=2.99e-07 $l=2.06761e-07 $layer=POLY_cond $X=0.345 $Y=2.085
+ $X2=0.38 $Y2=2.275
r37 1 11 0.573156 $w=1.7e-07 $l=7.8e-08 $layer=POLY_cond $X=0.345 $Y=1.385
+ $X2=0.345 $Y2=1.307
r38 1 2 295.965 $w=1.7e-07 $l=7e-07 $layer=POLY_cond $X=0.345 $Y=1.385 $X2=0.345
+ $Y2=2.085
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%A1 3 7 10 14 19
c43 19 0 5.77118e-21 $X=0.815 $Y=1.74
c44 10 0 3.09989e-20 $X=0.815 $Y=1.74
c45 7 0 1.78354e-19 $X=0.905 $Y=0.835
r46 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.815 $Y=1.74
+ $X2=0.815 $Y2=1.74
r47 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=1.74 $X2=0.815 $Y2=1.74
r48 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.815 $Y=1.74
+ $X2=0.815 $Y2=1.875
r49 10 11 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.815 $Y=1.74
+ $X2=0.815 $Y2=1.605
r50 7 11 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.905 $Y=0.835
+ $X2=0.905 $Y2=1.605
r51 3 12 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.835 $Y=3.235
+ $X2=0.835 $Y2=1.875
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%B0 3 7 10 15 20 23
c55 10 0 5.77118e-21 $X=1.325 $Y=1.85
r56 17 20 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.85
+ $X2=1.325 $Y2=1.85
r57 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.48 $X2=1.2
+ $Y2=2.48
r58 13 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=2.015 $X2=1.2
+ $Y2=1.85
r59 13 15 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.2 $Y=2.015
+ $X2=1.2 $Y2=2.48
r60 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.85 $X2=1.325 $Y2=1.85
r61 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.85
+ $X2=1.325 $Y2=2.015
r62 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.85
+ $X2=1.325 $Y2=1.685
r63 7 12 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.335 $Y=3.235
+ $X2=1.335 $Y2=2.015
r64 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.335 $Y=0.835
+ $X2=1.335 $Y2=1.685
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%B1 1 3 6 11 16
r24 11 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.005 $Y=2.115
+ $X2=2.005 $Y2=2.115
r25 9 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=2.115 $X2=2.005 $Y2=2.115
r26 4 9 38.7288 $w=3.45e-07 $l=2.16852e-07 $layer=POLY_cond $X=1.765 $Y=1.95
+ $X2=1.885 $Y2=2.115
r27 4 6 571.734 $w=1.5e-07 $l=1.115e-06 $layer=POLY_cond $X=1.765 $Y=1.95
+ $X2=1.765 $Y2=0.835
r28 1 9 72.2592 $w=3.45e-07 $l=4.90892e-07 $layer=POLY_cond $X=1.695 $Y=2.52
+ $X2=1.885 $Y2=2.115
r29 1 3 229.753 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.695 $Y=2.52
+ $X2=1.695 $Y2=3.235
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%Y 1 3 11 15 16 17 20 24
c41 24 0 3.09989e-20 $X=1.665 $Y=1.74
c42 17 0 1.78354e-19 $X=1.665 $Y=1.235
r43 20 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.665 $Y=1.74
+ $X2=1.665 $Y2=1.74
r44 18 20 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=1.665 $Y=2.745
+ $X2=1.665 $Y2=1.74
r45 17 22 12.496 $w=3.47e-07 $l=3.10153e-07 $layer=LI1_cond $X=1.665 $Y=1.235
+ $X2=1.567 $Y2=0.97
r46 17 20 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.665 $Y=1.235
+ $X2=1.665 $Y2=1.74
r47 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=2.83
+ $X2=1.665 $Y2=2.745
r48 15 16 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.58 $Y=2.83
+ $X2=1.17 $Y2=2.83
r49 11 13 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.085 $Y=3.01
+ $X2=1.085 $Y2=3.69
r50 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.085 $Y=2.915
+ $X2=1.17 $Y2=2.83
r51 9 11 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.085 $Y=2.915
+ $X2=1.085 $Y2=3.01
r52 3 13 400 $w=1.7e-07 $l=1.16923e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.605 $X2=1.085 $Y2=3.69
r53 3 11 400 $w=1.7e-07 $l=4.84665e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.605 $X2=1.085 $Y2=3.01
r54 1 22 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.97
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OAI22_L%A_27_115# 1 2 3 15 17 18 23 24 25
r32 25 28 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.98 $Y=0.63
+ $X2=1.98 $Y2=0.74
r33 23 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.63
+ $X2=1.98 $Y2=0.63
r34 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=0.63
+ $X2=1.205 $Y2=0.63
r35 20 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.12 $Y=1.075
+ $X2=1.12 $Y2=0.825
r36 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.715
+ $X2=1.205 $Y2=0.63
r37 19 22 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.12 $Y=0.715
+ $X2=1.12 $Y2=0.825
r38 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=1.12 $Y2=1.075
r39 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.345 $Y2=1.16
r40 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.345 $Y2=1.16
r41 13 15 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.26 $Y2=0.825
r42 3 28 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.74
r43 2 22 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r44 1 15 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

