* File: sky130_osu_sc_12T_hs__nand2_l.pex.spice
* Created: Fri Nov 12 15:11:52 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__NAND2_L%GND 1 17 19 26 33 36
r24 33 36 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r25 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r26 17 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r27 17 24 4.26217 $w=1.7e-07 $l=2.14243e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=1.05 $Y2=0.305
r28 17 19 3.29607 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=0.965 $Y2=0.152
r29 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r30 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__NAND2_L%VDD 1 2 17 21 23 30 35 38
r20 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r21 28 30 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.615
r22 26 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r23 24 33 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r24 24 26 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r25 23 28 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.135
r26 23 26 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r27 19 33 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r28 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.615
r29 17 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r30 17 33 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r31 2 30 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=3.025 $X2=1.12 $Y2=3.615
r32 1 21 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.615
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__NAND2_L%A 3 7 10 14 20
r32 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r33 14 17 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.32 $Y=2.575
+ $X2=0.32 $Y2=2.85
r34 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.575 $X2=0.32 $Y2=2.575
r35 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.575
+ $X2=0.367 $Y2=2.74
r36 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.575
+ $X2=0.367 $Y2=2.41
r37 7 12 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=3.445
+ $X2=0.475 $Y2=2.74
r38 3 11 833.245 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.475 $Y=0.785
+ $X2=0.475 $Y2=2.41
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__NAND2_L%B 3 7 10 14 19 22
c37 10 0 1.91696e-19 $X=0.915 $Y=1.825
c38 3 0 1.57512e-19 $X=0.835 $Y=0.785
r39 17 19 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.915 $Y=1.825
+ $X2=1.06 $Y2=1.825
r40 14 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.06 $Y=2.85
+ $X2=1.06 $Y2=2.85
r41 12 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.91
+ $X2=1.06 $Y2=1.825
r42 12 14 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.06 $Y=1.91
+ $X2=1.06 $Y2=2.85
r43 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=1.825 $X2=0.915 $Y2=1.825
r44 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.825
+ $X2=0.905 $Y2=1.66
r45 5 10 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.99
+ $X2=0.905 $Y2=1.825
r46 5 7 746.074 $w=1.5e-07 $l=1.455e-06 $layer=POLY_cond $X=0.905 $Y=1.99
+ $X2=0.905 $Y2=3.445
r47 3 11 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.835 $Y=0.785
+ $X2=0.835 $Y2=1.66
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__NAND2_L%Y 1 3 10 16 21 22 26 32
c37 22 0 1.57512e-19 $X=0.405 $Y=1.37
c38 16 0 1.91696e-19 $X=0.69 $Y=2.48
r39 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.48
r40 24 26 0.12036 $w=1.7e-07 $l=1.25e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.24
r41 23 26 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=0.69 $Y=1.455
+ $X2=0.69 $Y2=2.24
r42 22 29 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=1.37
+ $X2=0.26 $Y2=1.37
r43 21 23 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=1.37
+ $X2=0.69 $Y2=1.455
r44 21 22 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=1.37
+ $X2=0.405 $Y2=1.37
r45 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r46 16 19 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=3.615
r47 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=1.37
r48 10 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.26 $Y=0.74
+ $X2=0.26 $Y2=1.37
r49 3 19 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.025 $X2=0.69 $Y2=3.615
r50 1 10 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

