magic
tech sky130A
magscale 1 2
timestamp 1604007753
<< checkpaint >>
rect -1269 2461 1615 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1615 -1129
<< nwell >>
rect -9 529 355 1119
<< locali >>
rect 0 1049 352 1110
rect 0 0 352 61
<< metal1 >>
rect 0 1049 352 1110
rect 0 0 352 61
<< labels >>
rlabel metal1 196 30 196 30 1 gnd
rlabel metal1 199 1078 199 1078 1 vdd
<< end >>
