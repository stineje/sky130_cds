* File: sky130_osu_sc_15T_ms__dffsr_1.pxi.spice
* Created: Fri Nov 12 14:43:05 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%GND N_GND_M1017_s N_GND_M1033_s N_GND_M1000_d
+ N_GND_M1002_s N_GND_M1022_d N_GND_M1003_d N_GND_M1009_s N_GND_M1024_d
+ N_GND_M1004_d N_GND_M1017_b N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_14_p
+ N_GND_c_48_p N_GND_c_49_p N_GND_c_89_p N_GND_c_50_p N_GND_c_108_p N_GND_c_51_p
+ N_GND_c_113_p N_GND_c_52_p N_GND_c_17_p N_GND_c_18_p N_GND_c_193_p
+ N_GND_c_194_p GND N_GND_c_5_p PM_SKY130_OSU_SC_15T_MS__DFFSR_1%GND
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%VDD N_VDD_M1026_s N_VDD_M1010_d N_VDD_M1014_s
+ N_VDD_M1030_d N_VDD_M1015_d N_VDD_M1021_d N_VDD_M1016_d N_VDD_M1026_b
+ N_VDD_c_251_p N_VDD_c_252_p N_VDD_c_270_p N_VDD_c_285_p N_VDD_c_286_p
+ N_VDD_c_294_p N_VDD_c_279_p N_VDD_c_304_p N_VDD_c_280_p N_VDD_c_309_p
+ N_VDD_c_273_p N_VDD_c_263_p N_VDD_c_347_p N_VDD_c_363_p VDD N_VDD_c_253_p
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%VDD
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%RN N_RN_M1017_g N_RN_c_400_n N_RN_M1026_g
+ N_RN_c_402_n N_RN_c_403_n RN PM_SKY130_OSU_SC_15T_MS__DFFSR_1%RN
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_110_115# N_A_110_115#_M1017_d
+ N_A_110_115#_M1026_d N_A_110_115#_c_435_n N_A_110_115#_M1025_g
+ N_A_110_115#_c_437_n N_A_110_115#_M1033_g N_A_110_115#_c_441_n
+ N_A_110_115#_M1024_g N_A_110_115#_M1013_g N_A_110_115#_c_446_n
+ N_A_110_115#_c_447_n N_A_110_115#_c_448_n N_A_110_115#_c_450_n
+ N_A_110_115#_c_452_n N_A_110_115#_c_453_n N_A_110_115#_c_457_n
+ N_A_110_115#_c_458_n N_A_110_115#_c_459_n N_A_110_115#_c_461_n
+ N_A_110_115#_c_462_n N_A_110_115#_c_463_n N_A_110_115#_c_465_n
+ N_A_110_115#_c_467_n N_A_110_115#_c_479_n N_A_110_115#_c_481_n
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_110_115#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%SN N_SN_c_644_n N_SN_c_645_n N_SN_M1010_g
+ N_SN_M1011_g N_SN_M1001_g N_SN_M1007_g N_SN_c_654_n N_SN_c_655_n N_SN_c_656_n
+ N_SN_c_657_n N_SN_c_658_n N_SN_c_659_n N_SN_c_660_n N_SN_c_661_n SN
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%SN
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_432_468# N_A_432_468#_M1034_d
+ N_A_432_468#_M1005_d N_A_432_468#_M1000_g N_A_432_468#_M1012_g
+ N_A_432_468#_c_821_n N_A_432_468#_c_822_n N_A_432_468#_c_823_n
+ N_A_432_468#_c_826_n N_A_432_468#_c_838_n N_A_432_468#_c_868_n
+ N_A_432_468#_c_827_n N_A_432_468#_c_828_n N_A_432_468#_c_841_n
+ N_A_432_468#_c_849_n PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_432_468#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%D N_D_M1002_g N_D_M1014_g N_D_c_912_n
+ N_D_c_913_n D PM_SKY130_OSU_SC_15T_MS__DFFSR_1%D
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%CK N_CK_M1005_g N_CK_M1029_g N_CK_M1023_g
+ N_CK_M1027_g N_CK_M1008_g N_CK_c_946_n N_CK_M1020_g N_CK_c_947_n N_CK_c_948_n
+ N_CK_c_949_n N_CK_c_950_n N_CK_c_953_n N_CK_c_954_n N_CK_c_957_n N_CK_c_958_n
+ N_CK_c_963_n N_CK_c_964_n N_CK_c_965_n N_CK_c_966_n N_CK_c_967_n N_CK_c_968_n
+ N_CK_c_969_n N_CK_c_970_n N_CK_c_971_n N_CK_c_972_n N_CK_c_973_n N_CK_c_974_n
+ N_CK_c_975_n CK PM_SKY130_OSU_SC_15T_MS__DFFSR_1%CK
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_217_565# N_A_217_565#_M1033_d
+ N_A_217_565#_M1025_s N_A_217_565#_M1022_g N_A_217_565#_M1030_g
+ N_A_217_565#_c_1183_n N_A_217_565#_c_1185_n N_A_217_565#_c_1186_n
+ N_A_217_565#_c_1187_n N_A_217_565#_M1028_g N_A_217_565#_M1032_g
+ N_A_217_565#_c_1192_n N_A_217_565#_c_1193_n N_A_217_565#_c_1194_n
+ N_A_217_565#_c_1195_n N_A_217_565#_c_1198_n N_A_217_565#_c_1199_n
+ N_A_217_565#_c_1201_n N_A_217_565#_c_1202_n N_A_217_565#_c_1252_n
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_217_565#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_704_89# N_A_704_89#_M1008_d
+ N_A_704_89#_M1020_d N_A_704_89#_c_1344_n N_A_704_89#_M1034_g
+ N_A_704_89#_c_1347_n N_A_704_89#_c_1348_n N_A_704_89#_c_1349_n
+ N_A_704_89#_M1035_g N_A_704_89#_c_1351_n N_A_704_89#_M1031_g
+ N_A_704_89#_c_1353_n N_A_704_89#_c_1354_n N_A_704_89#_M1018_g
+ N_A_704_89#_c_1355_n N_A_704_89#_c_1356_n N_A_704_89#_c_1357_n
+ N_A_704_89#_c_1358_n N_A_704_89#_c_1359_n N_A_704_89#_c_1362_n
+ N_A_704_89#_c_1364_n N_A_704_89#_c_1369_n N_A_704_89#_c_1379_n
+ N_A_704_89#_c_1370_n N_A_704_89#_c_1371_n N_A_704_89#_c_1372_n
+ N_A_704_89#_c_1383_n PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_704_89#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_1246_89# N_A_1246_89#_M1001_d
+ N_A_1246_89#_M1013_d N_A_1246_89#_M1003_g N_A_1246_89#_M1015_g
+ N_A_1246_89#_M1004_g N_A_1246_89#_M1016_g N_A_1246_89#_c_1540_n
+ N_A_1246_89#_c_1541_n N_A_1246_89#_c_1542_n N_A_1246_89#_c_1543_n
+ N_A_1246_89#_c_1548_n N_A_1246_89#_c_1549_n N_A_1246_89#_c_1550_n
+ N_A_1246_89#_c_1551_n N_A_1246_89#_c_1552_n N_A_1246_89#_c_1555_n
+ N_A_1246_89#_c_1556_n N_A_1246_89#_c_1557_n N_A_1246_89#_c_1558_n
+ N_A_1246_89#_c_1559_n N_A_1246_89#_c_1560_n
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_1246_89#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_1084_115# N_A_1084_115#_M1023_d
+ N_A_1084_115#_M1031_d N_A_1084_115#_c_1707_n N_A_1084_115#_c_1708_n
+ N_A_1084_115#_M1009_g N_A_1084_115#_M1021_g N_A_1084_115#_c_1712_n
+ N_A_1084_115#_c_1714_n N_A_1084_115#_c_1715_n N_A_1084_115#_c_1740_n
+ N_A_1084_115#_c_1741_n N_A_1084_115#_c_1759_n N_A_1084_115#_c_1807_n
+ N_A_1084_115#_c_1716_n N_A_1084_115#_c_1732_n N_A_1084_115#_c_1719_n
+ N_A_1084_115#_c_1721_n N_A_1084_115#_c_1724_n N_A_1084_115#_c_1725_n
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_1084_115#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%QN N_QN_M1004_s N_QN_M1016_s N_QN_M1006_g
+ N_QN_M1019_g N_QN_c_1868_n N_QN_c_1869_n N_QN_c_1873_n N_QN_c_1874_n
+ N_QN_c_1876_n N_QN_c_1877_n N_QN_c_1878_n N_QN_c_1879_n QN
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%QN
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_300_565# N_A_300_565#_M1025_d
+ N_A_300_565#_M1012_d N_A_300_565#_c_1946_n N_A_300_565#_c_1949_n
+ N_A_300_565#_c_1960_n N_A_300_565#_c_1952_n
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_300_565#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_1469_565# N_A_1469_565#_M1021_s
+ N_A_1469_565#_M1007_d N_A_1469_565#_c_1970_n N_A_1469_565#_c_1973_n
+ N_A_1469_565#_c_1982_n N_A_1469_565#_c_1975_n
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%A_1469_565#
x_PM_SKY130_OSU_SC_15T_MS__DFFSR_1%Q N_Q_M1006_d N_Q_M1019_d N_Q_c_1989_n
+ N_Q_c_1993_n N_Q_c_1991_n N_Q_c_1992_n N_Q_c_1997_n Q
+ PM_SKY130_OSU_SC_15T_MS__DFFSR_1%Q
cc_1 N_GND_M1017_b N_RN_M1017_g 0.0635803f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_RN_M1017_g 0.00866533f $X=0.26 $Y=0.865 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_RN_M1017_g 0.00606474f $X=1.135 $Y=0.152 $X2=0.475 $Y2=0.945
cc_4 N_GND_c_4_p N_RN_M1017_g 0.0035726f $X=1.22 $Y=0.74 $X2=0.475 $Y2=0.945
cc_5 N_GND_c_5_p N_RN_M1017_g 0.00468827f $X=9.855 $Y=0.19 $X2=0.475 $Y2=0.945
cc_6 N_GND_M1017_b N_RN_c_400_n 0.0367521f $X=-0.05 $Y=0 $X2=0.475 $Y2=2.21
cc_7 N_GND_M1017_b N_RN_M1026_g 0.0318003f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.825
cc_8 N_GND_M1017_b N_RN_c_402_n 0.0149094f $X=-0.05 $Y=0 $X2=0.32 $Y2=3.07
cc_9 N_GND_M1017_b N_RN_c_403_n 0.0203125f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.045
cc_10 N_GND_M1017_b N_A_110_115#_c_435_n 0.0563099f $X=-0.05 $Y=0 $X2=1.29
+ $Y2=2.485
cc_11 N_GND_M1017_b N_A_110_115#_M1025_g 5.04534e-19 $X=-0.05 $Y=0 $X2=1.425
+ $Y2=3.825
cc_12 N_GND_M1017_b N_A_110_115#_c_437_n 0.0188039f $X=-0.05 $Y=0 $X2=1.435
+ $Y2=1.205
cc_13 N_GND_c_4_p N_A_110_115#_c_437_n 0.00502587f $X=1.22 $Y=0.74 $X2=1.435
+ $Y2=1.205
cc_14 N_GND_c_14_p N_A_110_115#_c_437_n 0.00606474f $X=2.415 $Y=0.152 $X2=1.435
+ $Y2=1.205
cc_15 N_GND_c_5_p N_A_110_115#_c_437_n 0.00468827f $X=9.855 $Y=0.19 $X2=1.435
+ $Y2=1.205
cc_16 N_GND_M1017_b N_A_110_115#_c_441_n 0.0186872f $X=-0.05 $Y=0 $X2=8.535
+ $Y2=1.205
cc_17 N_GND_c_17_p N_A_110_115#_c_441_n 0.00606474f $X=8.665 $Y=0.152 $X2=8.535
+ $Y2=1.205
cc_18 N_GND_c_18_p N_A_110_115#_c_441_n 0.00502587f $X=8.75 $Y=0.74 $X2=8.535
+ $Y2=1.205
cc_19 N_GND_c_5_p N_A_110_115#_c_441_n 0.00468827f $X=9.855 $Y=0.19 $X2=8.535
+ $Y2=1.205
cc_20 N_GND_M1017_b N_A_110_115#_M1013_g 5.06723e-19 $X=-0.05 $Y=0 $X2=8.545
+ $Y2=3.825
cc_21 N_GND_M1017_b N_A_110_115#_c_446_n 0.0508801f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=2.345
cc_22 N_GND_M1017_b N_A_110_115#_c_447_n 0.0211399f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=2.56
cc_23 N_GND_M1017_b N_A_110_115#_c_448_n 0.0418952f $X=-0.05 $Y=0 $X2=1.29
+ $Y2=1.37
cc_24 N_GND_c_4_p N_A_110_115#_c_448_n 0.00117914f $X=1.22 $Y=0.74 $X2=1.29
+ $Y2=1.37
cc_25 N_GND_M1017_b N_A_110_115#_c_450_n 0.0502942f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=1.37
cc_26 N_GND_c_18_p N_A_110_115#_c_450_n 0.00264977f $X=8.75 $Y=0.74 $X2=8.8
+ $Y2=1.37
cc_27 N_GND_M1017_b N_A_110_115#_c_452_n 0.0393083f $X=-0.05 $Y=0 $X2=8.545
+ $Y2=2.49
cc_28 N_GND_M1017_b N_A_110_115#_c_453_n 0.00156177f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=0.865
cc_29 N_GND_c_3_p N_A_110_115#_c_453_n 0.00760188f $X=1.135 $Y=0.152 $X2=0.69
+ $Y2=0.865
cc_30 N_GND_c_4_p N_A_110_115#_c_453_n 0.013807f $X=1.22 $Y=0.74 $X2=0.69
+ $Y2=0.865
cc_31 N_GND_c_5_p N_A_110_115#_c_453_n 0.00476945f $X=9.855 $Y=0.19 $X2=0.69
+ $Y2=0.865
cc_32 N_GND_M1017_b N_A_110_115#_c_457_n 0.00214428f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=3.205
cc_33 N_GND_M1017_b N_A_110_115#_c_458_n 0.0206181f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.395
cc_34 N_GND_M1017_b N_A_110_115#_c_459_n 0.0093348f $X=-0.05 $Y=0 $X2=1.145
+ $Y2=1.37
cc_35 N_GND_c_4_p N_A_110_115#_c_459_n 2.18563e-19 $X=1.22 $Y=0.74 $X2=1.145
+ $Y2=1.37
cc_36 N_GND_M1017_b N_A_110_115#_c_461_n 0.0133271f $X=-0.05 $Y=0 $X2=0.955
+ $Y2=1.37
cc_37 N_GND_M1017_b N_A_110_115#_c_462_n 0.0161505f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.48
cc_38 N_GND_M1017_b N_A_110_115#_c_463_n 0.00277795f $X=-0.05 $Y=0 $X2=1.23
+ $Y2=1.37
cc_39 N_GND_c_4_p N_A_110_115#_c_463_n 0.00841029f $X=1.22 $Y=0.74 $X2=1.23
+ $Y2=1.37
cc_40 N_GND_M1017_b N_A_110_115#_c_465_n 0.00613204f $X=-0.05 $Y=0 $X2=8.86
+ $Y2=1.22
cc_41 N_GND_c_18_p N_A_110_115#_c_465_n 0.00520267f $X=8.75 $Y=0.74 $X2=8.86
+ $Y2=1.22
cc_42 N_GND_M1000_d N_A_110_115#_c_467_n 0.00506015f $X=2.36 $Y=0.575 $X2=8.715
+ $Y2=1.22
cc_43 N_GND_M1002_s N_A_110_115#_c_467_n 0.00506021f $X=2.895 $Y=0.575 $X2=8.715
+ $Y2=1.22
cc_44 N_GND_M1022_d N_A_110_115#_c_467_n 0.0107322f $X=4.63 $Y=0.575 $X2=8.715
+ $Y2=1.22
cc_45 N_GND_M1003_d N_A_110_115#_c_467_n 0.00557645f $X=6.38 $Y=0.575 $X2=8.715
+ $Y2=1.22
cc_46 N_GND_M1009_s N_A_110_115#_c_467_n 0.00564702f $X=7.345 $Y=0.575 $X2=8.715
+ $Y2=1.22
cc_47 N_GND_M1017_b N_A_110_115#_c_467_n 0.0324342f $X=-0.05 $Y=0 $X2=8.715
+ $Y2=1.22
cc_48 N_GND_c_48_p N_A_110_115#_c_467_n 0.0118179f $X=2.5 $Y=0.865 $X2=8.715
+ $Y2=1.22
cc_49 N_GND_c_49_p N_A_110_115#_c_467_n 0.0118117f $X=3.02 $Y=0.865 $X2=8.715
+ $Y2=1.22
cc_50 N_GND_c_50_p N_A_110_115#_c_467_n 0.00602612f $X=4.77 $Y=0.74 $X2=8.715
+ $Y2=1.22
cc_51 N_GND_c_51_p N_A_110_115#_c_467_n 0.0119903f $X=6.52 $Y=0.865 $X2=8.715
+ $Y2=1.22
cc_52 N_GND_c_52_p N_A_110_115#_c_467_n 0.0139059f $X=7.47 $Y=0.865 $X2=8.715
+ $Y2=1.22
cc_53 N_GND_c_18_p N_A_110_115#_c_467_n 0.00198961f $X=8.75 $Y=0.74 $X2=8.715
+ $Y2=1.22
cc_54 N_GND_M1017_b N_A_110_115#_c_479_n 0.00688624f $X=-0.05 $Y=0 $X2=1.375
+ $Y2=1.22
cc_55 N_GND_c_4_p N_A_110_115#_c_479_n 0.00482641f $X=1.22 $Y=0.74 $X2=1.375
+ $Y2=1.22
cc_56 N_GND_M1017_b N_A_110_115#_c_481_n 0.00895912f $X=-0.05 $Y=0 $X2=8.86
+ $Y2=1.22
cc_57 N_GND_c_18_p N_A_110_115#_c_481_n 0.00356558f $X=8.75 $Y=0.74 $X2=8.86
+ $Y2=1.22
cc_58 N_GND_M1017_b N_SN_c_644_n 0.00804573f $X=-0.05 $Y=0 $X2=1.89 $Y2=1.625
cc_59 N_GND_M1017_b N_SN_c_645_n 0.0186775f $X=-0.05 $Y=0 $X2=1.89 $Y2=1.945
cc_60 N_GND_M1017_b N_SN_M1010_g 0.0180465f $X=-0.05 $Y=0 $X2=1.855 $Y2=3.825
cc_61 N_GND_M1017_b N_SN_M1011_g 0.0218297f $X=-0.05 $Y=0 $X2=1.925 $Y2=0.945
cc_62 N_GND_c_14_p N_SN_M1011_g 0.00606474f $X=2.415 $Y=0.152 $X2=1.925
+ $Y2=0.945
cc_63 N_GND_c_5_p N_SN_M1011_g 0.00468827f $X=9.855 $Y=0.19 $X2=1.925 $Y2=0.945
cc_64 N_GND_M1017_b N_SN_M1001_g 0.0429403f $X=-0.05 $Y=0 $X2=8.045 $Y2=0.945
cc_65 N_GND_c_17_p N_SN_M1001_g 0.00606474f $X=8.665 $Y=0.152 $X2=8.045
+ $Y2=0.945
cc_66 N_GND_c_5_p N_SN_M1001_g 0.00468827f $X=9.855 $Y=0.19 $X2=8.045 $Y2=0.945
cc_67 N_GND_M1017_b N_SN_M1007_g 0.0290585f $X=-0.05 $Y=0 $X2=8.115 $Y2=3.825
cc_68 N_GND_M1017_b N_SN_c_654_n 0.0380769f $X=-0.05 $Y=0 $X2=1.855 $Y2=2.11
cc_69 N_GND_M1017_b N_SN_c_655_n 0.0336181f $X=-0.05 $Y=0 $X2=8.025 $Y2=1.995
cc_70 N_GND_M1017_b N_SN_c_656_n 0.00274437f $X=-0.05 $Y=0 $X2=1.71 $Y2=2.7
cc_71 N_GND_M1017_b N_SN_c_657_n 0.00920532f $X=-0.05 $Y=0 $X2=7.935 $Y2=2.7
cc_72 N_GND_M1017_b N_SN_c_658_n 0.00222947f $X=-0.05 $Y=0 $X2=1.71 $Y2=2.11
cc_73 N_GND_M1017_b N_SN_c_659_n 0.00365816f $X=-0.05 $Y=0 $X2=8.025 $Y2=1.995
cc_74 N_GND_M1017_b N_SN_c_660_n 0.0528874f $X=-0.05 $Y=0 $X2=7.79 $Y2=2.7
cc_75 N_GND_M1017_b N_SN_c_661_n 0.00107924f $X=-0.05 $Y=0 $X2=1.855 $Y2=2.7
cc_76 N_GND_M1017_b SN 0.00268604f $X=-0.05 $Y=0 $X2=7.935 $Y2=2.7
cc_77 N_GND_M1017_b N_A_432_468#_M1000_g 0.0741657f $X=-0.05 $Y=0 $X2=2.285
+ $Y2=0.945
cc_78 N_GND_c_14_p N_A_432_468#_M1000_g 0.00606474f $X=2.415 $Y=0.152 $X2=2.285
+ $Y2=0.945
cc_79 N_GND_c_48_p N_A_432_468#_M1000_g 0.00868259f $X=2.5 $Y=0.865 $X2=2.285
+ $Y2=0.945
cc_80 N_GND_c_5_p N_A_432_468#_M1000_g 0.00468827f $X=9.855 $Y=0.19 $X2=2.285
+ $Y2=0.945
cc_81 N_GND_M1017_b N_A_432_468#_c_821_n 0.0343446f $X=-0.05 $Y=0 $X2=2.295
+ $Y2=2.505
cc_82 N_GND_M1017_b N_A_432_468#_c_822_n 0.0239207f $X=-0.05 $Y=0 $X2=2.295
+ $Y2=2.505
cc_83 N_GND_M1017_b N_A_432_468#_c_823_n 0.0278215f $X=-0.05 $Y=0 $X2=3.71
+ $Y2=1.505
cc_84 N_GND_c_48_p N_A_432_468#_c_823_n 0.00673409f $X=2.5 $Y=0.865 $X2=3.71
+ $Y2=1.505
cc_85 N_GND_c_49_p N_A_432_468#_c_823_n 0.00673409f $X=3.02 $Y=0.865 $X2=3.71
+ $Y2=1.505
cc_86 N_GND_M1017_b N_A_432_468#_c_826_n 0.00154034f $X=-0.05 $Y=0 $X2=2.38
+ $Y2=1.505
cc_87 N_GND_M1017_b N_A_432_468#_c_827_n 0.00198494f $X=-0.05 $Y=0 $X2=3.795
+ $Y2=1.42
cc_88 N_GND_M1017_b N_A_432_468#_c_828_n 0.00313474f $X=-0.05 $Y=0 $X2=3.895
+ $Y2=0.865
cc_89 N_GND_c_89_p N_A_432_468#_c_828_n 0.0148765f $X=4.685 $Y=0.152 $X2=3.895
+ $Y2=0.865
cc_90 N_GND_c_5_p N_A_432_468#_c_828_n 0.00955491f $X=9.855 $Y=0.19 $X2=3.895
+ $Y2=0.865
cc_91 N_GND_M1017_b N_D_M1002_g 0.0440753f $X=-0.05 $Y=0 $X2=3.235 $Y2=0.945
cc_92 N_GND_c_49_p N_D_M1002_g 0.0086813f $X=3.02 $Y=0.865 $X2=3.235 $Y2=0.945
cc_93 N_GND_c_89_p N_D_M1002_g 0.00606474f $X=4.685 $Y=0.152 $X2=3.235 $Y2=0.945
cc_94 N_GND_c_5_p N_D_M1002_g 0.00468827f $X=9.855 $Y=0.19 $X2=3.235 $Y2=0.945
cc_95 N_GND_M1017_b N_D_M1014_g 0.0445147f $X=-0.05 $Y=0 $X2=3.235 $Y2=3.825
cc_96 N_GND_M1017_b N_D_c_912_n 0.0337053f $X=-0.05 $Y=0 $X2=3.295 $Y2=1.96
cc_97 N_GND_M1017_b N_D_c_913_n 0.00170741f $X=-0.05 $Y=0 $X2=3.295 $Y2=1.96
cc_98 N_GND_M1017_b D 0.0155354f $X=-0.05 $Y=0 $X2=3.295 $Y2=1.96
cc_99 N_GND_M1017_b N_CK_c_946_n 0.0294225f $X=-0.05 $Y=0 $X2=6.735 $Y2=2.67
cc_100 N_GND_M1017_b N_CK_c_947_n 0.0432725f $X=-0.05 $Y=0 $X2=6.79 $Y2=2.34
cc_101 N_GND_M1017_b N_CK_c_948_n 0.0240652f $X=-0.05 $Y=0 $X2=3.655 $Y2=2.505
cc_102 N_GND_M1017_b N_CK_c_949_n 0.0254608f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.59
cc_103 N_GND_M1017_b N_CK_c_950_n 0.0173906f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.425
cc_104 N_GND_c_89_p N_CK_c_950_n 0.00606474f $X=4.685 $Y=0.152 $X2=4.135
+ $Y2=1.425
cc_105 N_GND_c_5_p N_CK_c_950_n 0.00468827f $X=9.855 $Y=0.19 $X2=4.135 $Y2=1.425
cc_106 N_GND_M1017_b N_CK_c_953_n 0.0252285f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.59
cc_107 N_GND_M1017_b N_CK_c_954_n 0.0175305f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.425
cc_108 N_GND_c_108_p N_CK_c_954_n 0.00606474f $X=6.435 $Y=0.152 $X2=5.405
+ $Y2=1.425
cc_109 N_GND_c_5_p N_CK_c_954_n 0.00468827f $X=9.855 $Y=0.19 $X2=5.405 $Y2=1.425
cc_110 N_GND_M1017_b N_CK_c_957_n 0.0230394f $X=-0.05 $Y=0 $X2=5.885 $Y2=2.505
cc_111 N_GND_M1017_b N_CK_c_958_n 0.0183851f $X=-0.05 $Y=0 $X2=6.762 $Y2=1.425
cc_112 N_GND_c_51_p N_CK_c_958_n 0.00390533f $X=6.52 $Y=0.865 $X2=6.762
+ $Y2=1.425
cc_113 N_GND_c_113_p N_CK_c_958_n 0.00606474f $X=7.385 $Y=0.152 $X2=6.762
+ $Y2=1.425
cc_114 N_GND_c_52_p N_CK_c_958_n 0.00409021f $X=7.47 $Y=0.865 $X2=6.762
+ $Y2=1.425
cc_115 N_GND_c_5_p N_CK_c_958_n 0.00468827f $X=9.855 $Y=0.19 $X2=6.762 $Y2=1.425
cc_116 N_GND_M1017_b N_CK_c_963_n 0.0130903f $X=-0.05 $Y=0 $X2=6.762 $Y2=1.575
cc_117 N_GND_M1017_b N_CK_c_964_n 0.00600607f $X=-0.05 $Y=0 $X2=4.05 $Y2=2.33
cc_118 N_GND_M1017_b N_CK_c_965_n 0.00921066f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.59
cc_119 N_GND_M1017_b N_CK_c_966_n 0.00838835f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.59
cc_120 N_GND_M1017_b N_CK_c_967_n 0.00543853f $X=-0.05 $Y=0 $X2=5.8 $Y2=2.33
cc_121 N_GND_M1017_b N_CK_c_968_n 5.00459e-19 $X=-0.05 $Y=0 $X2=5.49 $Y2=2.33
cc_122 N_GND_M1017_b N_CK_c_969_n 7.61111e-19 $X=-0.05 $Y=0 $X2=6.88 $Y2=2.33
cc_123 N_GND_M1017_b N_CK_c_970_n 0.00276905f $X=-0.05 $Y=0 $X2=3.655 $Y2=2.33
cc_124 N_GND_M1017_b N_CK_c_971_n 0.00265612f $X=-0.05 $Y=0 $X2=5.885 $Y2=2.33
cc_125 N_GND_M1017_b N_CK_c_972_n 0.0238264f $X=-0.05 $Y=0 $X2=5.74 $Y2=2.33
cc_126 N_GND_M1017_b N_CK_c_973_n 0.00704113f $X=-0.05 $Y=0 $X2=3.8 $Y2=2.33
cc_127 N_GND_M1017_b N_CK_c_974_n 0.00818551f $X=-0.05 $Y=0 $X2=6.735 $Y2=2.33
cc_128 N_GND_M1017_b N_CK_c_975_n 0.0038305f $X=-0.05 $Y=0 $X2=6.03 $Y2=2.33
cc_129 N_GND_M1017_b CK 0.00234237f $X=-0.05 $Y=0 $X2=6.88 $Y2=2.33
cc_130 N_GND_M1017_b N_A_217_565#_M1022_g 0.0171814f $X=-0.05 $Y=0 $X2=4.555
+ $Y2=0.945
cc_131 N_GND_c_89_p N_A_217_565#_M1022_g 0.00606474f $X=4.685 $Y=0.152 $X2=4.555
+ $Y2=0.945
cc_132 N_GND_c_50_p N_A_217_565#_M1022_g 0.00308284f $X=4.77 $Y=0.74 $X2=4.555
+ $Y2=0.945
cc_133 N_GND_c_5_p N_A_217_565#_M1022_g 0.00468827f $X=9.855 $Y=0.19 $X2=4.555
+ $Y2=0.945
cc_134 N_GND_M1017_b N_A_217_565#_c_1183_n 0.024077f $X=-0.05 $Y=0 $X2=4.91
+ $Y2=1.59
cc_135 N_GND_c_50_p N_A_217_565#_c_1183_n 8.60298e-19 $X=4.77 $Y=0.74 $X2=4.91
+ $Y2=1.59
cc_136 N_GND_M1017_b N_A_217_565#_c_1185_n 0.0105855f $X=-0.05 $Y=0 $X2=4.63
+ $Y2=1.59
cc_137 N_GND_M1017_b N_A_217_565#_c_1186_n 0.023252f $X=-0.05 $Y=0 $X2=4.91
+ $Y2=2.505
cc_138 N_GND_M1017_b N_A_217_565#_c_1187_n 0.0103717f $X=-0.05 $Y=0 $X2=4.63
+ $Y2=2.505
cc_139 N_GND_M1017_b N_A_217_565#_M1028_g 0.0163216f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=0.945
cc_140 N_GND_c_50_p N_A_217_565#_M1028_g 0.00308284f $X=4.77 $Y=0.74 $X2=4.985
+ $Y2=0.945
cc_141 N_GND_c_108_p N_A_217_565#_M1028_g 0.00606474f $X=6.435 $Y=0.152
+ $X2=4.985 $Y2=0.945
cc_142 N_GND_c_5_p N_A_217_565#_M1028_g 0.00468827f $X=9.855 $Y=0.19 $X2=4.985
+ $Y2=0.945
cc_143 N_GND_M1017_b N_A_217_565#_c_1192_n 0.00601555f $X=-0.05 $Y=0 $X2=1.21
+ $Y2=3.545
cc_144 N_GND_M1017_b N_A_217_565#_c_1193_n 0.00757526f $X=-0.05 $Y=0 $X2=1.625
+ $Y2=1.76
cc_145 N_GND_M1017_b N_A_217_565#_c_1194_n 0.00180429f $X=-0.05 $Y=0 $X2=1.295
+ $Y2=1.76
cc_146 N_GND_M1017_b N_A_217_565#_c_1195_n 0.00633193f $X=-0.05 $Y=0 $X2=1.71
+ $Y2=0.865
cc_147 N_GND_c_14_p N_A_217_565#_c_1195_n 0.00736239f $X=2.415 $Y=0.152 $X2=1.71
+ $Y2=0.865
cc_148 N_GND_c_5_p N_A_217_565#_c_1195_n 0.00476261f $X=9.855 $Y=0.19 $X2=1.71
+ $Y2=0.865
cc_149 N_GND_M1017_b N_A_217_565#_c_1198_n 0.0087185f $X=-0.05 $Y=0 $X2=4.725
+ $Y2=2.505
cc_150 N_GND_M1017_b N_A_217_565#_c_1199_n 0.00236783f $X=-0.05 $Y=0 $X2=4.725
+ $Y2=1.59
cc_151 N_GND_c_50_p N_A_217_565#_c_1199_n 0.00215957f $X=4.77 $Y=0.74 $X2=4.725
+ $Y2=1.59
cc_152 N_GND_M1017_b N_A_217_565#_c_1201_n 0.047915f $X=-0.05 $Y=0 $X2=4.49
+ $Y2=1.59
cc_153 N_GND_M1017_b N_A_217_565#_c_1202_n 0.00355505f $X=-0.05 $Y=0 $X2=1.855
+ $Y2=1.59
cc_154 N_GND_M1017_b N_A_704_89#_c_1344_n 0.0173059f $X=-0.05 $Y=0 $X2=3.595
+ $Y2=1.425
cc_155 N_GND_c_89_p N_A_704_89#_c_1344_n 0.00606474f $X=4.685 $Y=0.152 $X2=3.595
+ $Y2=1.425
cc_156 N_GND_c_5_p N_A_704_89#_c_1344_n 0.00468827f $X=9.855 $Y=0.19 $X2=3.595
+ $Y2=1.425
cc_157 N_GND_M1017_b N_A_704_89#_c_1347_n 0.0203057f $X=-0.05 $Y=0 $X2=3.715
+ $Y2=1.965
cc_158 N_GND_M1017_b N_A_704_89#_c_1348_n 0.0187566f $X=-0.05 $Y=0 $X2=4.12
+ $Y2=2.04
cc_159 N_GND_M1017_b N_A_704_89#_c_1349_n 0.00755029f $X=-0.05 $Y=0 $X2=3.79
+ $Y2=2.04
cc_160 N_GND_M1017_b N_A_704_89#_M1035_g 0.0321382f $X=-0.05 $Y=0 $X2=4.195
+ $Y2=3.825
cc_161 N_GND_M1017_b N_A_704_89#_c_1351_n 0.0559794f $X=-0.05 $Y=0 $X2=5.27
+ $Y2=2.04
cc_162 N_GND_M1017_b N_A_704_89#_M1031_g 0.0316517f $X=-0.05 $Y=0 $X2=5.345
+ $Y2=3.825
cc_163 N_GND_M1017_b N_A_704_89#_c_1353_n 0.0270462f $X=-0.05 $Y=0 $X2=5.75
+ $Y2=2.04
cc_164 N_GND_M1017_b N_A_704_89#_c_1354_n 0.0125754f $X=-0.05 $Y=0 $X2=5.825
+ $Y2=1.965
cc_165 N_GND_M1017_b N_A_704_89#_c_1355_n 0.0141451f $X=-0.05 $Y=0 $X2=3.715
+ $Y2=1.5
cc_166 N_GND_M1017_b N_A_704_89#_c_1356_n 0.00426512f $X=-0.05 $Y=0 $X2=4.195
+ $Y2=2.04
cc_167 N_GND_M1017_b N_A_704_89#_c_1357_n 0.00426512f $X=-0.05 $Y=0 $X2=5.345
+ $Y2=2.04
cc_168 N_GND_M1017_b N_A_704_89#_c_1358_n 0.0256431f $X=-0.05 $Y=0 $X2=5.885
+ $Y2=1.59
cc_169 N_GND_M1017_b N_A_704_89#_c_1359_n 0.01755f $X=-0.05 $Y=0 $X2=5.885
+ $Y2=1.425
cc_170 N_GND_c_108_p N_A_704_89#_c_1359_n 0.00606474f $X=6.435 $Y=0.152
+ $X2=5.885 $Y2=1.425
cc_171 N_GND_c_5_p N_A_704_89#_c_1359_n 0.00468827f $X=9.855 $Y=0.19 $X2=5.885
+ $Y2=1.425
cc_172 N_GND_M1017_b N_A_704_89#_c_1362_n 0.0116005f $X=-0.05 $Y=0 $X2=6.865
+ $Y2=1.59
cc_173 N_GND_c_51_p N_A_704_89#_c_1362_n 0.00564434f $X=6.52 $Y=0.865 $X2=6.865
+ $Y2=1.59
cc_174 N_GND_M1017_b N_A_704_89#_c_1364_n 0.00557295f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=0.865
cc_175 N_GND_c_51_p N_A_704_89#_c_1364_n 4.65312e-19 $X=6.52 $Y=0.865 $X2=6.95
+ $Y2=0.865
cc_176 N_GND_c_113_p N_A_704_89#_c_1364_n 0.0074445f $X=7.385 $Y=0.152 $X2=6.95
+ $Y2=0.865
cc_177 N_GND_c_52_p N_A_704_89#_c_1364_n 0.0245588f $X=7.47 $Y=0.865 $X2=6.95
+ $Y2=0.865
cc_178 N_GND_c_5_p N_A_704_89#_c_1364_n 0.00476261f $X=9.855 $Y=0.19 $X2=6.95
+ $Y2=0.865
cc_179 N_GND_M1017_b N_A_704_89#_c_1369_n 0.00299027f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=1.845
cc_180 N_GND_M1017_b N_A_704_89#_c_1370_n 0.011861f $X=-0.05 $Y=0 $X2=7.22
+ $Y2=2.84
cc_181 N_GND_M1017_b N_A_704_89#_c_1371_n 0.001308f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=1.59
cc_182 N_GND_M1017_b N_A_704_89#_c_1372_n 0.00945336f $X=-0.05 $Y=0 $X2=7.22
+ $Y2=1.93
cc_183 N_GND_M1017_b N_A_1246_89#_M1003_g 0.0319752f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=0.945
cc_184 N_GND_c_108_p N_A_1246_89#_M1003_g 0.00606474f $X=6.435 $Y=0.152
+ $X2=6.305 $Y2=0.945
cc_185 N_GND_c_51_p N_A_1246_89#_M1003_g 0.00394143f $X=6.52 $Y=0.865 $X2=6.305
+ $Y2=0.945
cc_186 N_GND_c_5_p N_A_1246_89#_M1003_g 0.00468827f $X=9.855 $Y=0.19 $X2=6.305
+ $Y2=0.945
cc_187 N_GND_M1017_b N_A_1246_89#_M1015_g 0.0327124f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=3.825
cc_188 N_GND_M1017_b N_A_1246_89#_c_1540_n 0.0263478f $X=-0.05 $Y=0 $X2=6.365
+ $Y2=1.93
cc_189 N_GND_M1017_b N_A_1246_89#_c_1541_n 0.0270403f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=1.93
cc_190 N_GND_M1017_b N_A_1246_89#_c_1542_n 0.0124759f $X=-0.05 $Y=0 $X2=9.382
+ $Y2=1.765
cc_191 N_GND_M1017_b N_A_1246_89#_c_1543_n 0.0165756f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=1.39
cc_192 N_GND_c_18_p N_A_1246_89#_c_1543_n 0.0035726f $X=8.75 $Y=0.74 $X2=9.47
+ $Y2=1.39
cc_193 N_GND_c_193_p N_A_1246_89#_c_1543_n 0.00606474f $X=9.625 $Y=0.152
+ $X2=9.47 $Y2=1.39
cc_194 N_GND_c_194_p N_A_1246_89#_c_1543_n 0.00388248f $X=9.71 $Y=0.865 $X2=9.47
+ $Y2=1.39
cc_195 N_GND_c_5_p N_A_1246_89#_c_1543_n 0.00468827f $X=9.855 $Y=0.19 $X2=9.47
+ $Y2=1.39
cc_196 N_GND_M1017_b N_A_1246_89#_c_1548_n 0.0132017f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=1.54
cc_197 N_GND_M1017_b N_A_1246_89#_c_1549_n 0.0284927f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=2.595
cc_198 N_GND_M1017_b N_A_1246_89#_c_1550_n 0.00455162f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=2.745
cc_199 N_GND_M1017_b N_A_1246_89#_c_1551_n 0.0039674f $X=-0.05 $Y=0 $X2=6.365
+ $Y2=1.93
cc_200 N_GND_M1017_b N_A_1246_89#_c_1552_n 0.00750073f $X=-0.05 $Y=0 $X2=8.26
+ $Y2=0.865
cc_201 N_GND_c_17_p N_A_1246_89#_c_1552_n 0.00750865f $X=8.665 $Y=0.152 $X2=8.26
+ $Y2=0.865
cc_202 N_GND_c_5_p N_A_1246_89#_c_1552_n 0.00476261f $X=9.855 $Y=0.19 $X2=8.26
+ $Y2=0.865
cc_203 N_GND_M1017_b N_A_1246_89#_c_1555_n 0.00494477f $X=-0.05 $Y=0 $X2=8.76
+ $Y2=3.545
cc_204 N_GND_M1017_b N_A_1246_89#_c_1556_n 0.020747f $X=-0.05 $Y=0 $X2=8.845
+ $Y2=1.93
cc_205 N_GND_M1017_b N_A_1246_89#_c_1557_n 0.0094386f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=1.93
cc_206 N_GND_M1017_b N_A_1246_89#_c_1558_n 0.056726f $X=-0.05 $Y=0 $X2=9.235
+ $Y2=1.93
cc_207 N_GND_M1017_b N_A_1246_89#_c_1559_n 0.00189525f $X=-0.05 $Y=0 $X2=6.51
+ $Y2=1.93
cc_208 N_GND_M1017_b N_A_1246_89#_c_1560_n 0.0014645f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=1.93
cc_209 N_GND_M1017_b N_A_1084_115#_c_1707_n 0.0450481f $X=-0.05 $Y=0 $X2=7.505
+ $Y2=2.37
cc_210 N_GND_M1017_b N_A_1084_115#_c_1708_n 0.0178887f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.43
cc_211 N_GND_c_52_p N_A_1084_115#_c_1708_n 0.00868259f $X=7.47 $Y=0.865
+ $X2=7.685 $Y2=1.43
cc_212 N_GND_c_17_p N_A_1084_115#_c_1708_n 0.00606474f $X=8.665 $Y=0.152
+ $X2=7.685 $Y2=1.43
cc_213 N_GND_c_5_p N_A_1084_115#_c_1708_n 0.00468827f $X=9.855 $Y=0.19 $X2=7.685
+ $Y2=1.43
cc_214 N_GND_M1017_b N_A_1084_115#_c_1712_n 0.0235095f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.51
cc_215 N_GND_c_52_p N_A_1084_115#_c_1712_n 0.00391038f $X=7.47 $Y=0.865
+ $X2=7.685 $Y2=1.51
cc_216 N_GND_M1017_b N_A_1084_115#_c_1714_n 0.0324837f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=2.505
cc_217 N_GND_M1017_b N_A_1084_115#_c_1715_n 0.011286f $X=-0.05 $Y=0 $X2=5.065
+ $Y2=1.59
cc_218 N_GND_M1017_b N_A_1084_115#_c_1716_n 0.00313975f $X=-0.05 $Y=0 $X2=5.645
+ $Y2=0.865
cc_219 N_GND_c_108_p N_A_1084_115#_c_1716_n 0.0149333f $X=6.435 $Y=0.152
+ $X2=5.645 $Y2=0.865
cc_220 N_GND_c_5_p N_A_1084_115#_c_1716_n 0.00958198f $X=9.855 $Y=0.19 $X2=5.645
+ $Y2=0.865
cc_221 N_GND_M1017_b N_A_1084_115#_c_1719_n 0.00582616f $X=-0.05 $Y=0 $X2=7.595
+ $Y2=1.59
cc_222 N_GND_c_52_p N_A_1084_115#_c_1719_n 0.00131024f $X=7.47 $Y=0.865
+ $X2=7.595 $Y2=1.59
cc_223 N_GND_M1017_b N_A_1084_115#_c_1721_n 0.022645f $X=-0.05 $Y=0 $X2=7.45
+ $Y2=1.59
cc_224 N_GND_c_51_p N_A_1084_115#_c_1721_n 5.03331e-19 $X=6.52 $Y=0.865 $X2=7.45
+ $Y2=1.59
cc_225 N_GND_c_52_p N_A_1084_115#_c_1721_n 3.1624e-19 $X=7.47 $Y=0.865 $X2=7.45
+ $Y2=1.59
cc_226 N_GND_M1017_b N_A_1084_115#_c_1724_n 0.00120467f $X=-0.05 $Y=0 $X2=5.21
+ $Y2=1.59
cc_227 N_GND_M1017_b N_A_1084_115#_c_1725_n 0.00169121f $X=-0.05 $Y=0 $X2=7.595
+ $Y2=1.59
cc_228 N_GND_c_52_p N_A_1084_115#_c_1725_n 4.00959e-19 $X=7.47 $Y=0.865
+ $X2=7.595 $Y2=1.59
cc_229 N_GND_M1017_b N_QN_M1006_g 0.0561552f $X=-0.05 $Y=0 $X2=9.925 $Y2=0.945
cc_230 N_GND_c_194_p N_QN_M1006_g 0.00388248f $X=9.71 $Y=0.865 $X2=9.925
+ $Y2=0.945
cc_231 N_GND_c_5_p N_QN_M1006_g 0.00468827f $X=9.855 $Y=0.19 $X2=9.925 $Y2=0.945
cc_232 N_GND_M1017_b N_QN_M1019_g 0.0186095f $X=-0.05 $Y=0 $X2=9.925 $Y2=3.825
cc_233 N_GND_M1017_b N_QN_c_1868_n 0.0291912f $X=-0.05 $Y=0 $X2=9.865 $Y2=2.135
cc_234 N_GND_M1017_b N_QN_c_1869_n 0.00463899f $X=-0.05 $Y=0 $X2=9.28 $Y2=0.865
cc_235 N_GND_c_18_p N_QN_c_1869_n 0.013807f $X=8.75 $Y=0.74 $X2=9.28 $Y2=0.865
cc_236 N_GND_c_193_p N_QN_c_1869_n 0.00736239f $X=9.625 $Y=0.152 $X2=9.28
+ $Y2=0.865
cc_237 N_GND_c_5_p N_QN_c_1869_n 0.00476261f $X=9.855 $Y=0.19 $X2=9.28 $Y2=0.865
cc_238 N_GND_M1017_b N_QN_c_1873_n 0.00102655f $X=-0.05 $Y=0 $X2=9.28 $Y2=2.7
cc_239 N_GND_M1017_b N_QN_c_1874_n 0.0133445f $X=-0.05 $Y=0 $X2=9.78 $Y2=1.59
cc_240 N_GND_c_194_p N_QN_c_1874_n 0.00827206f $X=9.71 $Y=0.865 $X2=9.78
+ $Y2=1.59
cc_241 N_GND_M1017_b N_QN_c_1876_n 0.00291105f $X=-0.05 $Y=0 $X2=9.365 $Y2=1.59
cc_242 N_GND_M1017_b N_QN_c_1877_n 0.0138424f $X=-0.05 $Y=0 $X2=9.78 $Y2=2.505
cc_243 N_GND_M1017_b N_QN_c_1878_n 0.00301984f $X=-0.05 $Y=0 $X2=9.365 $Y2=2.505
cc_244 N_GND_M1017_b N_QN_c_1879_n 0.0034889f $X=-0.05 $Y=0 $X2=9.865 $Y2=2.135
cc_245 N_GND_M1017_b QN 0.00258296f $X=-0.05 $Y=0 $X2=9.285 $Y2=2.7
cc_246 N_GND_M1017_b N_Q_c_1989_n 0.00905638f $X=-0.05 $Y=0 $X2=10.14 $Y2=0.865
cc_247 N_GND_c_5_p N_Q_c_1989_n 0.00474182f $X=9.855 $Y=0.19 $X2=10.14 $Y2=0.865
cc_248 N_GND_M1017_b N_Q_c_1991_n 0.0625704f $X=-0.05 $Y=0 $X2=10.255 $Y2=2.745
cc_249 N_GND_M1017_b N_Q_c_1992_n 0.0140324f $X=-0.05 $Y=0 $X2=10.255 $Y2=1.255
cc_250 N_VDD_M1026_b N_RN_M1026_g 0.0270317f $X=-0.05 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_251 N_VDD_c_251_p N_RN_M1026_g 0.00751602f $X=0.26 $Y=3.885 $X2=0.475
+ $Y2=3.825
cc_252 N_VDD_c_252_p N_RN_M1026_g 0.00496961f $X=1.985 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_253 N_VDD_c_253_p N_RN_M1026_g 0.00429146f $X=9.855 $Y=5.36 $X2=0.475
+ $Y2=3.825
cc_254 N_VDD_M1026_s N_RN_c_402_n 0.00953431f $X=0.135 $Y=2.825 $X2=0.32
+ $Y2=3.07
cc_255 N_VDD_M1026_b N_RN_c_402_n 0.00618364f $X=-0.05 $Y=2.645 $X2=0.32
+ $Y2=3.07
cc_256 N_VDD_c_251_p N_RN_c_402_n 0.00252874f $X=0.26 $Y=3.885 $X2=0.32 $Y2=3.07
cc_257 N_VDD_M1026_s RN 0.0162774f $X=0.135 $Y=2.825 $X2=0.325 $Y2=3.07
cc_258 N_VDD_c_251_p RN 0.00522047f $X=0.26 $Y=3.885 $X2=0.325 $Y2=3.07
cc_259 N_VDD_M1026_b N_A_110_115#_M1025_g 0.0250337f $X=-0.05 $Y=2.645 $X2=1.425
+ $Y2=3.825
cc_260 N_VDD_c_252_p N_A_110_115#_M1025_g 0.00496961f $X=1.985 $Y=5.397
+ $X2=1.425 $Y2=3.825
cc_261 N_VDD_c_253_p N_A_110_115#_M1025_g 0.00429146f $X=9.855 $Y=5.36 $X2=1.425
+ $Y2=3.825
cc_262 N_VDD_M1026_b N_A_110_115#_M1013_g 0.0250679f $X=-0.05 $Y=2.645 $X2=8.545
+ $Y2=3.825
cc_263 N_VDD_c_263_p N_A_110_115#_M1013_g 0.00496961f $X=9.625 $Y=5.397
+ $X2=8.545 $Y2=3.825
cc_264 N_VDD_c_253_p N_A_110_115#_M1013_g 0.00429146f $X=9.855 $Y=5.36 $X2=8.545
+ $Y2=3.825
cc_265 N_VDD_M1026_b N_A_110_115#_c_457_n 0.00593582f $X=-0.05 $Y=2.645 $X2=0.69
+ $Y2=3.205
cc_266 N_VDD_c_252_p N_A_110_115#_c_457_n 0.00477009f $X=1.985 $Y=5.397 $X2=0.69
+ $Y2=3.205
cc_267 N_VDD_c_253_p N_A_110_115#_c_457_n 0.00435496f $X=9.855 $Y=5.36 $X2=0.69
+ $Y2=3.205
cc_268 N_VDD_M1026_b N_SN_M1010_g 0.0192489f $X=-0.05 $Y=2.645 $X2=1.855
+ $Y2=3.825
cc_269 N_VDD_c_252_p N_SN_M1010_g 0.00496961f $X=1.985 $Y=5.397 $X2=1.855
+ $Y2=3.825
cc_270 N_VDD_c_270_p N_SN_M1010_g 0.00362996f $X=2.07 $Y=3.885 $X2=1.855
+ $Y2=3.825
cc_271 N_VDD_c_253_p N_SN_M1010_g 0.00429146f $X=9.855 $Y=5.36 $X2=1.855
+ $Y2=3.825
cc_272 N_VDD_M1026_b N_SN_M1007_g 0.0201131f $X=-0.05 $Y=2.645 $X2=8.115
+ $Y2=3.825
cc_273 N_VDD_c_273_p N_SN_M1007_g 0.00362996f $X=7.9 $Y=3.885 $X2=8.115
+ $Y2=3.825
cc_274 N_VDD_c_263_p N_SN_M1007_g 0.00496961f $X=9.625 $Y=5.397 $X2=8.115
+ $Y2=3.825
cc_275 N_VDD_c_253_p N_SN_M1007_g 0.00429146f $X=9.855 $Y=5.36 $X2=8.115
+ $Y2=3.825
cc_276 N_VDD_M1026_b N_SN_c_656_n 0.00205457f $X=-0.05 $Y=2.645 $X2=1.71 $Y2=2.7
cc_277 N_VDD_M1026_b N_SN_c_657_n 0.00449283f $X=-0.05 $Y=2.645 $X2=7.935
+ $Y2=2.7
cc_278 N_VDD_M1026_b N_SN_c_660_n 0.0566252f $X=-0.05 $Y=2.645 $X2=7.79 $Y2=2.7
cc_279 N_VDD_c_279_p N_SN_c_660_n 0.00464215f $X=4.77 $Y=3.545 $X2=7.79 $Y2=2.7
cc_280 N_VDD_c_280_p N_SN_c_660_n 0.0090257f $X=6.52 $Y=3.205 $X2=7.79 $Y2=2.7
cc_281 N_VDD_M1026_b N_SN_c_661_n 0.00372061f $X=-0.05 $Y=2.645 $X2=1.855
+ $Y2=2.7
cc_282 N_VDD_M1026_b SN 0.00292685f $X=-0.05 $Y=2.645 $X2=7.935 $Y2=2.7
cc_283 N_VDD_M1026_b N_A_432_468#_M1012_g 0.0217743f $X=-0.05 $Y=2.645 $X2=2.285
+ $Y2=3.825
cc_284 N_VDD_c_270_p N_A_432_468#_M1012_g 0.00362996f $X=2.07 $Y=3.885 $X2=2.285
+ $Y2=3.825
cc_285 N_VDD_c_285_p N_A_432_468#_M1012_g 0.00496961f $X=2.935 $Y=5.397
+ $X2=2.285 $Y2=3.825
cc_286 N_VDD_c_286_p N_A_432_468#_M1012_g 0.00620001f $X=3.02 $Y=3.545 $X2=2.285
+ $Y2=3.825
cc_287 N_VDD_c_253_p N_A_432_468#_M1012_g 0.00429146f $X=9.855 $Y=5.36 $X2=2.285
+ $Y2=3.825
cc_288 N_VDD_M1026_b N_A_432_468#_c_821_n 0.0057899f $X=-0.05 $Y=2.645 $X2=2.295
+ $Y2=2.505
cc_289 N_VDD_M1026_b N_A_432_468#_c_822_n 0.00281226f $X=-0.05 $Y=2.645
+ $X2=2.295 $Y2=2.505
cc_290 N_VDD_M1014_s N_A_432_468#_c_838_n 0.00705065f $X=2.895 $Y=2.825
+ $X2=3.725 $Y2=2.925
cc_291 N_VDD_M1026_b N_A_432_468#_c_838_n 0.013691f $X=-0.05 $Y=2.645 $X2=3.725
+ $Y2=2.925
cc_292 N_VDD_c_286_p N_A_432_468#_c_838_n 0.00850976f $X=3.02 $Y=3.545 $X2=3.725
+ $Y2=2.925
cc_293 N_VDD_M1026_b N_A_432_468#_c_841_n 0.00402069f $X=-0.05 $Y=2.645
+ $X2=3.895 $Y2=3.205
cc_294 N_VDD_c_294_p N_A_432_468#_c_841_n 0.00928728f $X=4.685 $Y=5.397
+ $X2=3.895 $Y2=3.205
cc_295 N_VDD_c_253_p N_A_432_468#_c_841_n 0.00876183f $X=9.855 $Y=5.36 $X2=3.895
+ $Y2=3.205
cc_296 N_VDD_M1026_b N_D_M1014_g 0.0228684f $X=-0.05 $Y=2.645 $X2=3.235
+ $Y2=3.825
cc_297 N_VDD_c_286_p N_D_M1014_g 0.00751602f $X=3.02 $Y=3.545 $X2=3.235
+ $Y2=3.825
cc_298 N_VDD_c_294_p N_D_M1014_g 0.00496961f $X=4.685 $Y=5.397 $X2=3.235
+ $Y2=3.825
cc_299 N_VDD_c_253_p N_D_M1014_g 0.00429146f $X=9.855 $Y=5.36 $X2=3.235
+ $Y2=3.825
cc_300 N_VDD_M1026_b N_CK_M1005_g 0.0192734f $X=-0.05 $Y=2.645 $X2=3.595
+ $Y2=3.825
cc_301 N_VDD_c_294_p N_CK_M1005_g 0.00496961f $X=4.685 $Y=5.397 $X2=3.595
+ $Y2=3.825
cc_302 N_VDD_c_253_p N_CK_M1005_g 0.00429146f $X=9.855 $Y=5.36 $X2=3.595
+ $Y2=3.825
cc_303 N_VDD_M1026_b N_CK_M1027_g 0.0192734f $X=-0.05 $Y=2.645 $X2=5.945
+ $Y2=3.825
cc_304 N_VDD_c_304_p N_CK_M1027_g 0.00496961f $X=6.435 $Y=5.397 $X2=5.945
+ $Y2=3.825
cc_305 N_VDD_c_253_p N_CK_M1027_g 0.00429146f $X=9.855 $Y=5.36 $X2=5.945
+ $Y2=3.825
cc_306 N_VDD_M1026_b N_CK_c_946_n 0.007968f $X=-0.05 $Y=2.645 $X2=6.735 $Y2=2.67
cc_307 N_VDD_M1026_b N_CK_M1020_g 0.0245312f $X=-0.05 $Y=2.645 $X2=6.735
+ $Y2=3.825
cc_308 N_VDD_c_280_p N_CK_M1020_g 0.00362996f $X=6.52 $Y=3.205 $X2=6.735
+ $Y2=3.825
cc_309 N_VDD_c_309_p N_CK_M1020_g 0.00496961f $X=7.815 $Y=5.397 $X2=6.735
+ $Y2=3.825
cc_310 N_VDD_c_253_p N_CK_M1020_g 0.00429146f $X=9.855 $Y=5.36 $X2=6.735
+ $Y2=3.825
cc_311 N_VDD_M1026_b N_CK_c_948_n 0.00508175f $X=-0.05 $Y=2.645 $X2=3.655
+ $Y2=2.505
cc_312 N_VDD_M1026_b N_CK_c_957_n 0.00508175f $X=-0.05 $Y=2.645 $X2=5.885
+ $Y2=2.505
cc_313 N_VDD_M1026_b N_CK_c_969_n 0.0010436f $X=-0.05 $Y=2.645 $X2=6.88 $Y2=2.33
cc_314 N_VDD_M1026_b N_CK_c_970_n 2.35021e-19 $X=-0.05 $Y=2.645 $X2=3.655
+ $Y2=2.33
cc_315 N_VDD_M1026_b N_CK_c_971_n 7.56914e-19 $X=-0.05 $Y=2.645 $X2=5.885
+ $Y2=2.33
cc_316 N_VDD_M1026_b N_A_217_565#_M1030_g 0.0182924f $X=-0.05 $Y=2.645 $X2=4.555
+ $Y2=3.825
cc_317 N_VDD_c_294_p N_A_217_565#_M1030_g 0.00496961f $X=4.685 $Y=5.397
+ $X2=4.555 $Y2=3.825
cc_318 N_VDD_c_279_p N_A_217_565#_M1030_g 0.00362996f $X=4.77 $Y=3.545 $X2=4.555
+ $Y2=3.825
cc_319 N_VDD_c_253_p N_A_217_565#_M1030_g 0.00429146f $X=9.855 $Y=5.36 $X2=4.555
+ $Y2=3.825
cc_320 N_VDD_c_279_p N_A_217_565#_c_1186_n 7.6376e-19 $X=4.77 $Y=3.545 $X2=4.91
+ $Y2=2.505
cc_321 N_VDD_M1026_b N_A_217_565#_M1032_g 0.0179418f $X=-0.05 $Y=2.645 $X2=4.985
+ $Y2=3.825
cc_322 N_VDD_c_279_p N_A_217_565#_M1032_g 0.00362996f $X=4.77 $Y=3.545 $X2=4.985
+ $Y2=3.825
cc_323 N_VDD_c_304_p N_A_217_565#_M1032_g 0.00496961f $X=6.435 $Y=5.397
+ $X2=4.985 $Y2=3.825
cc_324 N_VDD_c_253_p N_A_217_565#_M1032_g 0.00429146f $X=9.855 $Y=5.36 $X2=4.985
+ $Y2=3.825
cc_325 N_VDD_M1026_b N_A_217_565#_c_1192_n 0.00480682f $X=-0.05 $Y=2.645
+ $X2=1.21 $Y2=3.545
cc_326 N_VDD_c_252_p N_A_217_565#_c_1192_n 0.00463398f $X=1.985 $Y=5.397
+ $X2=1.21 $Y2=3.545
cc_327 N_VDD_c_253_p N_A_217_565#_c_1192_n 0.00435496f $X=9.855 $Y=5.36 $X2=1.21
+ $Y2=3.545
cc_328 N_VDD_M1026_b N_A_217_565#_c_1198_n 0.00208967f $X=-0.05 $Y=2.645
+ $X2=4.725 $Y2=2.505
cc_329 N_VDD_c_279_p N_A_217_565#_c_1198_n 0.00215846f $X=4.77 $Y=3.545
+ $X2=4.725 $Y2=2.505
cc_330 N_VDD_M1026_b N_A_704_89#_M1035_g 0.0203819f $X=-0.05 $Y=2.645 $X2=4.195
+ $Y2=3.825
cc_331 N_VDD_c_294_p N_A_704_89#_M1035_g 0.00496961f $X=4.685 $Y=5.397 $X2=4.195
+ $Y2=3.825
cc_332 N_VDD_c_253_p N_A_704_89#_M1035_g 0.00429146f $X=9.855 $Y=5.36 $X2=4.195
+ $Y2=3.825
cc_333 N_VDD_M1026_b N_A_704_89#_M1031_g 0.0203747f $X=-0.05 $Y=2.645 $X2=5.345
+ $Y2=3.825
cc_334 N_VDD_c_304_p N_A_704_89#_M1031_g 0.00496961f $X=6.435 $Y=5.397 $X2=5.345
+ $Y2=3.825
cc_335 N_VDD_c_253_p N_A_704_89#_M1031_g 0.00429146f $X=9.855 $Y=5.36 $X2=5.345
+ $Y2=3.825
cc_336 N_VDD_M1026_b N_A_704_89#_c_1379_n 0.00199838f $X=-0.05 $Y=2.645 $X2=6.95
+ $Y2=3.205
cc_337 N_VDD_c_309_p N_A_704_89#_c_1379_n 0.00461951f $X=7.815 $Y=5.397 $X2=6.95
+ $Y2=3.205
cc_338 N_VDD_c_253_p N_A_704_89#_c_1379_n 0.00435496f $X=9.855 $Y=5.36 $X2=6.95
+ $Y2=3.205
cc_339 N_VDD_M1026_b N_A_704_89#_c_1370_n 0.00526199f $X=-0.05 $Y=2.645 $X2=7.22
+ $Y2=2.84
cc_340 N_VDD_M1026_b N_A_704_89#_c_1383_n 0.012303f $X=-0.05 $Y=2.645 $X2=7.22
+ $Y2=2.925
cc_341 N_VDD_M1026_b N_A_1246_89#_M1015_g 0.0186387f $X=-0.05 $Y=2.645 $X2=6.305
+ $Y2=3.825
cc_342 N_VDD_c_304_p N_A_1246_89#_M1015_g 0.00496961f $X=6.435 $Y=5.397
+ $X2=6.305 $Y2=3.825
cc_343 N_VDD_c_280_p N_A_1246_89#_M1015_g 0.00362996f $X=6.52 $Y=3.205 $X2=6.305
+ $Y2=3.825
cc_344 N_VDD_c_253_p N_A_1246_89#_M1015_g 0.00429146f $X=9.855 $Y=5.36 $X2=6.305
+ $Y2=3.825
cc_345 N_VDD_M1026_b N_A_1246_89#_c_1550_n 0.0293418f $X=-0.05 $Y=2.645 $X2=9.47
+ $Y2=2.745
cc_346 N_VDD_c_263_p N_A_1246_89#_c_1550_n 0.00496961f $X=9.625 $Y=5.397
+ $X2=9.47 $Y2=2.745
cc_347 N_VDD_c_347_p N_A_1246_89#_c_1550_n 0.00362996f $X=9.71 $Y=3.205 $X2=9.47
+ $Y2=2.745
cc_348 N_VDD_c_253_p N_A_1246_89#_c_1550_n 0.00429146f $X=9.855 $Y=5.36 $X2=9.47
+ $Y2=2.745
cc_349 N_VDD_M1026_b N_A_1246_89#_c_1555_n 0.00484331f $X=-0.05 $Y=2.645
+ $X2=8.76 $Y2=3.545
cc_350 N_VDD_c_263_p N_A_1246_89#_c_1555_n 0.00473534f $X=9.625 $Y=5.397
+ $X2=8.76 $Y2=3.545
cc_351 N_VDD_c_253_p N_A_1246_89#_c_1555_n 0.00435496f $X=9.855 $Y=5.36 $X2=8.76
+ $Y2=3.545
cc_352 N_VDD_M1026_b N_A_1084_115#_M1021_g 0.0258774f $X=-0.05 $Y=2.645
+ $X2=7.685 $Y2=3.825
cc_353 N_VDD_c_309_p N_A_1084_115#_M1021_g 0.00496961f $X=7.815 $Y=5.397
+ $X2=7.685 $Y2=3.825
cc_354 N_VDD_c_273_p N_A_1084_115#_M1021_g 0.00362996f $X=7.9 $Y=3.885 $X2=7.685
+ $Y2=3.825
cc_355 N_VDD_c_253_p N_A_1084_115#_M1021_g 0.00429146f $X=9.855 $Y=5.36
+ $X2=7.685 $Y2=3.825
cc_356 N_VDD_M1026_b N_A_1084_115#_c_1715_n 0.00207418f $X=-0.05 $Y=2.645
+ $X2=5.065 $Y2=1.59
cc_357 N_VDD_M1026_b N_A_1084_115#_c_1732_n 0.00402069f $X=-0.05 $Y=2.645
+ $X2=5.645 $Y2=3.545
cc_358 N_VDD_c_304_p N_A_1084_115#_c_1732_n 0.00924384f $X=6.435 $Y=5.397
+ $X2=5.645 $Y2=3.545
cc_359 N_VDD_c_253_p N_A_1084_115#_c_1732_n 0.00876183f $X=9.855 $Y=5.36
+ $X2=5.645 $Y2=3.545
cc_360 N_VDD_M1026_b N_A_1084_115#_c_1719_n 9.87966e-19 $X=-0.05 $Y=2.645
+ $X2=7.595 $Y2=1.59
cc_361 N_VDD_M1026_b N_QN_M1019_g 0.0251095f $X=-0.05 $Y=2.645 $X2=9.925
+ $Y2=3.825
cc_362 N_VDD_c_347_p N_QN_M1019_g 0.00362996f $X=9.71 $Y=3.205 $X2=9.925
+ $Y2=3.825
cc_363 N_VDD_c_363_p N_QN_M1019_g 0.00496961f $X=9.855 $Y=5.33 $X2=9.925
+ $Y2=3.825
cc_364 N_VDD_c_253_p N_QN_M1019_g 0.00429146f $X=9.855 $Y=5.36 $X2=9.925
+ $Y2=3.825
cc_365 N_VDD_M1026_b N_QN_c_1873_n 0.0057559f $X=-0.05 $Y=2.645 $X2=9.28 $Y2=2.7
cc_366 N_VDD_c_263_p N_QN_c_1873_n 0.00452684f $X=9.625 $Y=5.397 $X2=9.28
+ $Y2=2.7
cc_367 N_VDD_c_253_p N_QN_c_1873_n 0.00435496f $X=9.855 $Y=5.36 $X2=9.28 $Y2=2.7
cc_368 N_VDD_c_347_p N_QN_c_1877_n 0.00818856f $X=9.71 $Y=3.205 $X2=9.78
+ $Y2=2.505
cc_369 N_VDD_M1026_b QN 0.0101088f $X=-0.05 $Y=2.645 $X2=9.285 $Y2=2.7
cc_370 N_VDD_M1026_b N_A_300_565#_c_1946_n 0.00198641f $X=-0.05 $Y=2.645
+ $X2=1.64 $Y2=3.545
cc_371 N_VDD_c_252_p N_A_300_565#_c_1946_n 0.0045126f $X=1.985 $Y=5.397 $X2=1.64
+ $Y2=3.545
cc_372 N_VDD_c_253_p N_A_300_565#_c_1946_n 0.00434939f $X=9.855 $Y=5.36 $X2=1.64
+ $Y2=3.545
cc_373 N_VDD_M1010_d N_A_300_565#_c_1949_n 0.00482635f $X=1.93 $Y=2.825
+ $X2=2.415 $Y2=3.37
cc_374 N_VDD_c_270_p N_A_300_565#_c_1949_n 0.0135055f $X=2.07 $Y=3.885 $X2=2.415
+ $Y2=3.37
cc_375 N_VDD_c_286_p N_A_300_565#_c_1949_n 0.00811594f $X=3.02 $Y=3.545
+ $X2=2.415 $Y2=3.37
cc_376 N_VDD_M1026_b N_A_300_565#_c_1952_n 0.00199838f $X=-0.05 $Y=2.645 $X2=2.5
+ $Y2=3.545
cc_377 N_VDD_c_285_p N_A_300_565#_c_1952_n 0.00453263f $X=2.935 $Y=5.397 $X2=2.5
+ $Y2=3.545
cc_378 N_VDD_c_286_p N_A_300_565#_c_1952_n 0.0585029f $X=3.02 $Y=3.545 $X2=2.5
+ $Y2=3.545
cc_379 N_VDD_c_253_p N_A_300_565#_c_1952_n 0.00435496f $X=9.855 $Y=5.36 $X2=2.5
+ $Y2=3.545
cc_380 N_VDD_M1026_b N_A_1469_565#_c_1970_n 0.00199838f $X=-0.05 $Y=2.645
+ $X2=7.47 $Y2=3.545
cc_381 N_VDD_c_309_p N_A_1469_565#_c_1970_n 0.00477009f $X=7.815 $Y=5.397
+ $X2=7.47 $Y2=3.545
cc_382 N_VDD_c_253_p N_A_1469_565#_c_1970_n 0.00435496f $X=9.855 $Y=5.36
+ $X2=7.47 $Y2=3.545
cc_383 N_VDD_M1021_d N_A_1469_565#_c_1973_n 0.00462014f $X=7.76 $Y=2.825
+ $X2=8.245 $Y2=3.37
cc_384 N_VDD_c_273_p N_A_1469_565#_c_1973_n 0.0135055f $X=7.9 $Y=3.885 $X2=8.245
+ $Y2=3.37
cc_385 N_VDD_M1026_b N_A_1469_565#_c_1975_n 0.00198641f $X=-0.05 $Y=2.645
+ $X2=8.33 $Y2=3.545
cc_386 N_VDD_c_263_p N_A_1469_565#_c_1975_n 0.00457631f $X=9.625 $Y=5.397
+ $X2=8.33 $Y2=3.545
cc_387 N_VDD_c_253_p N_A_1469_565#_c_1975_n 0.00434939f $X=9.855 $Y=5.36
+ $X2=8.33 $Y2=3.545
cc_388 N_VDD_M1026_b N_Q_c_1993_n 0.00199838f $X=-0.05 $Y=2.645 $X2=10.14
+ $Y2=3.07
cc_389 N_VDD_c_363_p N_Q_c_1993_n 0.00476429f $X=9.855 $Y=5.33 $X2=10.14
+ $Y2=3.07
cc_390 N_VDD_c_253_p N_Q_c_1993_n 0.00435496f $X=9.855 $Y=5.36 $X2=10.14
+ $Y2=3.07
cc_391 N_VDD_M1026_b N_Q_c_1991_n 0.00544948f $X=-0.05 $Y=2.645 $X2=10.255
+ $Y2=2.745
cc_392 N_VDD_M1026_b N_Q_c_1997_n 0.0144447f $X=-0.05 $Y=2.645 $X2=10.255
+ $Y2=2.83
cc_393 N_VDD_M1026_b Q 0.00983408f $X=-0.05 $Y=2.645 $X2=10.14 $Y2=3.07
cc_394 N_VDD_c_347_p Q 0.00673193f $X=9.71 $Y=3.205 $X2=10.14 $Y2=3.07
cc_395 RN N_A_110_115#_M1026_d 0.00414531f $X=0.325 $Y=3.07 $X2=0.55 $Y2=2.825
cc_396 N_RN_M1017_g N_A_110_115#_c_435_n 0.00347101f $X=0.475 $Y=0.945 $X2=1.29
+ $Y2=2.485
cc_397 N_RN_c_400_n N_A_110_115#_c_435_n 0.00491728f $X=0.475 $Y=2.21 $X2=1.29
+ $Y2=2.485
cc_398 N_RN_M1026_g N_A_110_115#_c_435_n 0.00426455f $X=0.475 $Y=3.825 $X2=1.29
+ $Y2=2.485
cc_399 N_RN_M1017_g N_A_110_115#_c_448_n 0.0050047f $X=0.475 $Y=0.945 $X2=1.29
+ $Y2=1.37
cc_400 N_RN_M1026_g N_A_110_115#_c_457_n 0.0100254f $X=0.475 $Y=3.825 $X2=0.69
+ $Y2=3.205
cc_401 N_RN_c_402_n N_A_110_115#_c_457_n 0.0282684f $X=0.32 $Y=3.07 $X2=0.69
+ $Y2=3.205
cc_402 RN N_A_110_115#_c_457_n 0.00974028f $X=0.325 $Y=3.07 $X2=0.69 $Y2=3.205
cc_403 N_RN_M1017_g N_A_110_115#_c_458_n 0.00939617f $X=0.475 $Y=0.945 $X2=0.87
+ $Y2=2.395
cc_404 N_RN_c_400_n N_A_110_115#_c_458_n 0.00325637f $X=0.475 $Y=2.21 $X2=0.87
+ $Y2=2.395
cc_405 N_RN_M1026_g N_A_110_115#_c_458_n 0.00186244f $X=0.475 $Y=3.825 $X2=0.87
+ $Y2=2.395
cc_406 N_RN_c_402_n N_A_110_115#_c_458_n 0.0072511f $X=0.32 $Y=3.07 $X2=0.87
+ $Y2=2.395
cc_407 N_RN_c_403_n N_A_110_115#_c_458_n 0.0248372f $X=0.32 $Y=2.045 $X2=0.87
+ $Y2=2.395
cc_408 N_RN_M1017_g N_A_110_115#_c_461_n 0.00501976f $X=0.475 $Y=0.945 $X2=0.955
+ $Y2=1.37
cc_409 N_RN_c_400_n N_A_110_115#_c_461_n 0.00149212f $X=0.475 $Y=2.21 $X2=0.955
+ $Y2=1.37
cc_410 N_RN_c_403_n N_A_110_115#_c_461_n 3.79578e-19 $X=0.32 $Y=2.045 $X2=0.955
+ $Y2=1.37
cc_411 N_RN_c_400_n N_A_110_115#_c_462_n 0.00191737f $X=0.475 $Y=2.21 $X2=0.87
+ $Y2=2.48
cc_412 N_RN_M1026_g N_A_110_115#_c_462_n 0.00207383f $X=0.475 $Y=3.825 $X2=0.87
+ $Y2=2.48
cc_413 N_RN_c_402_n N_A_110_115#_c_462_n 0.0113366f $X=0.32 $Y=3.07 $X2=0.87
+ $Y2=2.48
cc_414 N_RN_c_403_n N_A_110_115#_c_462_n 7.08415e-19 $X=0.32 $Y=2.045 $X2=0.87
+ $Y2=2.48
cc_415 N_RN_M1026_g N_A_217_565#_c_1192_n 0.00502509f $X=0.475 $Y=3.825 $X2=1.21
+ $Y2=3.545
cc_416 RN N_A_217_565#_c_1192_n 9.10636e-19 $X=0.325 $Y=3.07 $X2=1.21 $Y2=3.545
cc_417 N_A_110_115#_c_448_n N_SN_c_644_n 0.00566608f $X=1.29 $Y=1.37 $X2=1.89
+ $Y2=1.625
cc_418 N_A_110_115#_c_467_n N_SN_c_644_n 2.91248e-19 $X=8.715 $Y=1.22 $X2=1.89
+ $Y2=1.625
cc_419 N_A_110_115#_c_435_n N_SN_c_645_n 0.00566608f $X=1.29 $Y=2.485 $X2=1.89
+ $Y2=1.945
cc_420 N_A_110_115#_c_435_n N_SN_M1010_g 0.00495566f $X=1.29 $Y=2.485 $X2=1.855
+ $Y2=3.825
cc_421 N_A_110_115#_c_447_n N_SN_M1010_g 0.0464682f $X=1.425 $Y=2.56 $X2=1.855
+ $Y2=3.825
cc_422 N_A_110_115#_c_437_n N_SN_M1011_g 0.0230282f $X=1.435 $Y=1.205 $X2=1.925
+ $Y2=0.945
cc_423 N_A_110_115#_c_448_n N_SN_M1011_g 0.00298272f $X=1.29 $Y=1.37 $X2=1.925
+ $Y2=0.945
cc_424 N_A_110_115#_c_467_n N_SN_M1011_g 0.0106787f $X=8.715 $Y=1.22 $X2=1.925
+ $Y2=0.945
cc_425 N_A_110_115#_c_441_n N_SN_M1001_g 0.023075f $X=8.535 $Y=1.205 $X2=8.045
+ $Y2=0.945
cc_426 N_A_110_115#_c_450_n N_SN_M1001_g 0.00540313f $X=8.8 $Y=1.37 $X2=8.045
+ $Y2=0.945
cc_427 N_A_110_115#_c_467_n N_SN_M1001_g 0.0110943f $X=8.715 $Y=1.22 $X2=8.045
+ $Y2=0.945
cc_428 N_A_110_115#_c_452_n N_SN_M1007_g 0.0505287f $X=8.545 $Y=2.49 $X2=8.115
+ $Y2=3.825
cc_429 N_A_110_115#_c_435_n N_SN_c_654_n 0.0200438f $X=1.29 $Y=2.485 $X2=1.855
+ $Y2=2.11
cc_430 N_A_110_115#_c_446_n N_SN_c_655_n 0.00890342f $X=8.8 $Y=2.345 $X2=8.025
+ $Y2=1.995
cc_431 N_A_110_115#_c_467_n N_SN_c_655_n 0.00212668f $X=8.715 $Y=1.22 $X2=8.025
+ $Y2=1.995
cc_432 N_A_110_115#_c_435_n N_SN_c_656_n 0.00177359f $X=1.29 $Y=2.485 $X2=1.71
+ $Y2=2.7
cc_433 N_A_110_115#_c_447_n N_SN_c_656_n 0.00231894f $X=1.425 $Y=2.56 $X2=1.71
+ $Y2=2.7
cc_434 N_A_110_115#_c_435_n N_SN_c_658_n 0.00103414f $X=1.29 $Y=2.485 $X2=1.71
+ $Y2=2.11
cc_435 N_A_110_115#_c_446_n N_SN_c_659_n 2.72295e-19 $X=8.8 $Y=2.345 $X2=8.025
+ $Y2=1.995
cc_436 N_A_110_115#_c_467_n N_SN_c_659_n 0.00342638f $X=8.715 $Y=1.22 $X2=8.025
+ $Y2=1.995
cc_437 N_A_110_115#_c_447_n N_SN_c_661_n 0.00457686f $X=1.425 $Y=2.56 $X2=1.855
+ $Y2=2.7
cc_438 N_A_110_115#_c_452_n SN 0.00110631f $X=8.545 $Y=2.49 $X2=7.935 $Y2=2.7
cc_439 N_A_110_115#_c_467_n N_A_432_468#_M1034_d 0.00558831f $X=8.715 $Y=1.22
+ $X2=3.67 $Y2=0.575
cc_440 N_A_110_115#_c_467_n N_A_432_468#_M1000_g 0.0116352f $X=8.715 $Y=1.22
+ $X2=2.285 $Y2=0.945
cc_441 N_A_110_115#_c_467_n N_A_432_468#_c_823_n 0.0295499f $X=8.715 $Y=1.22
+ $X2=3.71 $Y2=1.505
cc_442 N_A_110_115#_c_467_n N_A_432_468#_c_826_n 0.00540043f $X=8.715 $Y=1.22
+ $X2=2.38 $Y2=1.505
cc_443 N_A_110_115#_c_467_n N_A_432_468#_c_827_n 0.0151351f $X=8.715 $Y=1.22
+ $X2=3.795 $Y2=1.42
cc_444 N_A_110_115#_c_467_n N_A_432_468#_c_849_n 0.0253593f $X=8.715 $Y=1.22
+ $X2=3.887 $Y2=1.155
cc_445 N_A_110_115#_c_467_n N_D_M1002_g 0.0116357f $X=8.715 $Y=1.22 $X2=3.235
+ $Y2=0.945
cc_446 N_A_110_115#_c_467_n N_CK_c_949_n 8.06574e-19 $X=8.715 $Y=1.22 $X2=4.135
+ $Y2=1.59
cc_447 N_A_110_115#_c_467_n N_CK_c_950_n 0.0106495f $X=8.715 $Y=1.22 $X2=4.135
+ $Y2=1.425
cc_448 N_A_110_115#_c_467_n N_CK_c_953_n 8.06574e-19 $X=8.715 $Y=1.22 $X2=5.405
+ $Y2=1.59
cc_449 N_A_110_115#_c_467_n N_CK_c_954_n 0.00177838f $X=8.715 $Y=1.22 $X2=5.405
+ $Y2=1.425
cc_450 N_A_110_115#_c_467_n N_CK_c_958_n 0.01159f $X=8.715 $Y=1.22 $X2=6.762
+ $Y2=1.425
cc_451 N_A_110_115#_c_467_n N_CK_c_963_n 0.00107886f $X=8.715 $Y=1.22 $X2=6.762
+ $Y2=1.575
cc_452 N_A_110_115#_c_467_n N_CK_c_965_n 0.00496158f $X=8.715 $Y=1.22 $X2=4.135
+ $Y2=1.59
cc_453 N_A_110_115#_c_467_n N_CK_c_966_n 0.00118606f $X=8.715 $Y=1.22 $X2=5.405
+ $Y2=1.59
cc_454 N_A_110_115#_c_467_n N_A_217_565#_M1033_d 0.00428739f $X=8.715 $Y=1.22
+ $X2=1.51 $Y2=0.575
cc_455 N_A_110_115#_c_467_n N_A_217_565#_M1022_g 0.0104272f $X=8.715 $Y=1.22
+ $X2=4.555 $Y2=0.945
cc_456 N_A_110_115#_c_467_n N_A_217_565#_c_1183_n 2.42482e-19 $X=8.715 $Y=1.22
+ $X2=4.91 $Y2=1.59
cc_457 N_A_110_115#_c_467_n N_A_217_565#_M1028_g 0.00491871f $X=8.715 $Y=1.22
+ $X2=4.985 $Y2=0.945
cc_458 N_A_110_115#_c_435_n N_A_217_565#_c_1192_n 0.0189043f $X=1.29 $Y=2.485
+ $X2=1.21 $Y2=3.545
cc_459 N_A_110_115#_M1025_g N_A_217_565#_c_1192_n 0.0164398f $X=1.425 $Y=3.825
+ $X2=1.21 $Y2=3.545
cc_460 N_A_110_115#_c_447_n N_A_217_565#_c_1192_n 0.00689282f $X=1.425 $Y=2.56
+ $X2=1.21 $Y2=3.545
cc_461 N_A_110_115#_c_457_n N_A_217_565#_c_1192_n 0.0963044f $X=0.69 $Y=3.205
+ $X2=1.21 $Y2=3.545
cc_462 N_A_110_115#_c_458_n N_A_217_565#_c_1192_n 0.041373f $X=0.87 $Y=2.395
+ $X2=1.21 $Y2=3.545
cc_463 N_A_110_115#_c_462_n N_A_217_565#_c_1192_n 0.0134429f $X=0.87 $Y=2.48
+ $X2=1.21 $Y2=3.545
cc_464 N_A_110_115#_c_435_n N_A_217_565#_c_1193_n 0.00783536f $X=1.29 $Y=2.485
+ $X2=1.625 $Y2=1.76
cc_465 N_A_110_115#_c_447_n N_A_217_565#_c_1193_n 0.00344703f $X=1.425 $Y=2.56
+ $X2=1.625 $Y2=1.76
cc_466 N_A_110_115#_c_448_n N_A_217_565#_c_1193_n 0.00422528f $X=1.29 $Y=1.37
+ $X2=1.625 $Y2=1.76
cc_467 N_A_110_115#_c_463_n N_A_217_565#_c_1193_n 0.00525465f $X=1.23 $Y=1.37
+ $X2=1.625 $Y2=1.76
cc_468 N_A_110_115#_c_467_n N_A_217_565#_c_1193_n 0.00645017f $X=8.715 $Y=1.22
+ $X2=1.625 $Y2=1.76
cc_469 N_A_110_115#_c_479_n N_A_217_565#_c_1193_n 4.15231e-19 $X=1.375 $Y=1.22
+ $X2=1.625 $Y2=1.76
cc_470 N_A_110_115#_c_435_n N_A_217_565#_c_1194_n 0.00463903f $X=1.29 $Y=2.485
+ $X2=1.295 $Y2=1.76
cc_471 N_A_110_115#_c_448_n N_A_217_565#_c_1194_n 0.00225048f $X=1.29 $Y=1.37
+ $X2=1.295 $Y2=1.76
cc_472 N_A_110_115#_c_458_n N_A_217_565#_c_1194_n 0.0142869f $X=0.87 $Y=2.395
+ $X2=1.295 $Y2=1.76
cc_473 N_A_110_115#_c_459_n N_A_217_565#_c_1194_n 0.0011521f $X=1.145 $Y=1.37
+ $X2=1.295 $Y2=1.76
cc_474 N_A_110_115#_c_463_n N_A_217_565#_c_1194_n 0.00901695f $X=1.23 $Y=1.37
+ $X2=1.295 $Y2=1.76
cc_475 N_A_110_115#_c_479_n N_A_217_565#_c_1194_n 0.00105745f $X=1.375 $Y=1.22
+ $X2=1.295 $Y2=1.76
cc_476 N_A_110_115#_c_437_n N_A_217_565#_c_1195_n 0.00980314f $X=1.435 $Y=1.205
+ $X2=1.71 $Y2=0.865
cc_477 N_A_110_115#_c_448_n N_A_217_565#_c_1195_n 0.00232106f $X=1.29 $Y=1.37
+ $X2=1.71 $Y2=0.865
cc_478 N_A_110_115#_c_458_n N_A_217_565#_c_1195_n 0.00354634f $X=0.87 $Y=2.395
+ $X2=1.71 $Y2=0.865
cc_479 N_A_110_115#_c_463_n N_A_217_565#_c_1195_n 0.0161718f $X=1.23 $Y=1.37
+ $X2=1.71 $Y2=0.865
cc_480 N_A_110_115#_c_467_n N_A_217_565#_c_1195_n 0.0229218f $X=8.715 $Y=1.22
+ $X2=1.71 $Y2=0.865
cc_481 N_A_110_115#_c_479_n N_A_217_565#_c_1195_n 0.00144419f $X=1.375 $Y=1.22
+ $X2=1.71 $Y2=0.865
cc_482 N_A_110_115#_c_467_n N_A_217_565#_c_1199_n 0.00527975f $X=8.715 $Y=1.22
+ $X2=4.725 $Y2=1.59
cc_483 N_A_110_115#_c_467_n N_A_217_565#_c_1201_n 0.212985f $X=8.715 $Y=1.22
+ $X2=4.49 $Y2=1.59
cc_484 N_A_110_115#_c_448_n N_A_217_565#_c_1202_n 0.00392729f $X=1.29 $Y=1.37
+ $X2=1.855 $Y2=1.59
cc_485 N_A_110_115#_c_458_n N_A_217_565#_c_1202_n 0.0049761f $X=0.87 $Y=2.395
+ $X2=1.855 $Y2=1.59
cc_486 N_A_110_115#_c_467_n N_A_217_565#_c_1202_n 0.0252928f $X=8.715 $Y=1.22
+ $X2=1.855 $Y2=1.59
cc_487 N_A_110_115#_c_467_n N_A_217_565#_c_1252_n 0.0259207f $X=8.715 $Y=1.22
+ $X2=4.635 $Y2=1.59
cc_488 N_A_110_115#_c_467_n N_A_704_89#_M1008_d 0.00421798f $X=8.715 $Y=1.22
+ $X2=6.81 $Y2=0.575
cc_489 N_A_110_115#_c_467_n N_A_704_89#_c_1344_n 0.0102209f $X=8.715 $Y=1.22
+ $X2=3.595 $Y2=1.425
cc_490 N_A_110_115#_c_467_n N_A_704_89#_c_1358_n 0.00232964f $X=8.715 $Y=1.22
+ $X2=5.885 $Y2=1.59
cc_491 N_A_110_115#_c_467_n N_A_704_89#_c_1359_n 0.0103799f $X=8.715 $Y=1.22
+ $X2=5.885 $Y2=1.425
cc_492 N_A_110_115#_c_467_n N_A_704_89#_c_1362_n 0.0115848f $X=8.715 $Y=1.22
+ $X2=6.865 $Y2=1.59
cc_493 N_A_110_115#_c_467_n N_A_704_89#_c_1364_n 0.0252668f $X=8.715 $Y=1.22
+ $X2=6.95 $Y2=0.865
cc_494 N_A_110_115#_c_467_n N_A_704_89#_c_1372_n 4.8388e-19 $X=8.715 $Y=1.22
+ $X2=7.22 $Y2=1.93
cc_495 N_A_110_115#_c_467_n N_A_1246_89#_M1001_d 0.00453588f $X=8.715 $Y=1.22
+ $X2=8.12 $Y2=0.575
cc_496 N_A_110_115#_c_467_n N_A_1246_89#_M1003_g 0.0100216f $X=8.715 $Y=1.22
+ $X2=6.305 $Y2=0.945
cc_497 N_A_110_115#_c_446_n N_A_1246_89#_c_1541_n 0.0112463f $X=8.8 $Y=2.345
+ $X2=9.38 $Y2=1.93
cc_498 N_A_110_115#_c_450_n N_A_1246_89#_c_1543_n 0.00434527f $X=8.8 $Y=1.37
+ $X2=9.47 $Y2=1.39
cc_499 N_A_110_115#_c_446_n N_A_1246_89#_c_1548_n 0.00524146f $X=8.8 $Y=2.345
+ $X2=9.47 $Y2=1.54
cc_500 N_A_110_115#_c_450_n N_A_1246_89#_c_1548_n 0.00385786f $X=8.8 $Y=1.37
+ $X2=9.47 $Y2=1.54
cc_501 N_A_110_115#_c_446_n N_A_1246_89#_c_1549_n 0.00978182f $X=8.8 $Y=2.345
+ $X2=9.47 $Y2=2.595
cc_502 N_A_110_115#_c_452_n N_A_1246_89#_c_1549_n 0.00180274f $X=8.545 $Y=2.49
+ $X2=9.47 $Y2=2.595
cc_503 N_A_110_115#_c_441_n N_A_1246_89#_c_1552_n 0.0100938f $X=8.535 $Y=1.205
+ $X2=8.26 $Y2=0.865
cc_504 N_A_110_115#_c_450_n N_A_1246_89#_c_1552_n 0.0024217f $X=8.8 $Y=1.37
+ $X2=8.26 $Y2=0.865
cc_505 N_A_110_115#_c_465_n N_A_1246_89#_c_1552_n 0.0109701f $X=8.86 $Y=1.22
+ $X2=8.26 $Y2=0.865
cc_506 N_A_110_115#_c_467_n N_A_1246_89#_c_1552_n 0.0256238f $X=8.715 $Y=1.22
+ $X2=8.26 $Y2=0.865
cc_507 N_A_110_115#_c_481_n N_A_1246_89#_c_1552_n 0.0014036f $X=8.86 $Y=1.22
+ $X2=8.26 $Y2=0.865
cc_508 N_A_110_115#_M1013_g N_A_1246_89#_c_1555_n 0.0169896f $X=8.545 $Y=3.825
+ $X2=8.76 $Y2=3.545
cc_509 N_A_110_115#_c_446_n N_A_1246_89#_c_1555_n 0.0115916f $X=8.8 $Y=2.345
+ $X2=8.76 $Y2=3.545
cc_510 N_A_110_115#_c_452_n N_A_1246_89#_c_1555_n 0.0174648f $X=8.545 $Y=2.49
+ $X2=8.76 $Y2=3.545
cc_511 N_A_110_115#_c_446_n N_A_1246_89#_c_1556_n 0.0121067f $X=8.8 $Y=2.345
+ $X2=8.845 $Y2=1.93
cc_512 N_A_110_115#_c_450_n N_A_1246_89#_c_1556_n 0.00693473f $X=8.8 $Y=1.37
+ $X2=8.845 $Y2=1.93
cc_513 N_A_110_115#_c_452_n N_A_1246_89#_c_1556_n 0.0054736f $X=8.545 $Y=2.49
+ $X2=8.845 $Y2=1.93
cc_514 N_A_110_115#_c_465_n N_A_1246_89#_c_1556_n 0.00372046f $X=8.86 $Y=1.22
+ $X2=8.845 $Y2=1.93
cc_515 N_A_110_115#_c_467_n N_A_1246_89#_c_1556_n 0.00679066f $X=8.715 $Y=1.22
+ $X2=8.845 $Y2=1.93
cc_516 N_A_110_115#_c_481_n N_A_1246_89#_c_1556_n 3.23811e-19 $X=8.86 $Y=1.22
+ $X2=8.845 $Y2=1.93
cc_517 N_A_110_115#_c_446_n N_A_1246_89#_c_1557_n 0.0039999f $X=8.8 $Y=2.345
+ $X2=9.38 $Y2=1.93
cc_518 N_A_110_115#_c_450_n N_A_1246_89#_c_1557_n 0.0023935f $X=8.8 $Y=1.37
+ $X2=9.38 $Y2=1.93
cc_519 N_A_110_115#_c_465_n N_A_1246_89#_c_1557_n 0.00479193f $X=8.86 $Y=1.22
+ $X2=9.38 $Y2=1.93
cc_520 N_A_110_115#_c_446_n N_A_1246_89#_c_1558_n 0.00275467f $X=8.8 $Y=2.345
+ $X2=9.235 $Y2=1.93
cc_521 N_A_110_115#_c_450_n N_A_1246_89#_c_1558_n 0.00187493f $X=8.8 $Y=1.37
+ $X2=9.235 $Y2=1.93
cc_522 N_A_110_115#_c_465_n N_A_1246_89#_c_1558_n 0.00255174f $X=8.86 $Y=1.22
+ $X2=9.235 $Y2=1.93
cc_523 N_A_110_115#_c_467_n N_A_1246_89#_c_1558_n 0.044242f $X=8.715 $Y=1.22
+ $X2=9.235 $Y2=1.93
cc_524 N_A_110_115#_c_481_n N_A_1246_89#_c_1558_n 0.0129068f $X=8.86 $Y=1.22
+ $X2=9.235 $Y2=1.93
cc_525 N_A_110_115#_c_446_n N_A_1246_89#_c_1560_n 8.29185e-19 $X=8.8 $Y=2.345
+ $X2=9.38 $Y2=1.93
cc_526 N_A_110_115#_c_467_n N_A_1084_115#_M1023_d 0.0051762f $X=8.715 $Y=1.22
+ $X2=5.42 $Y2=0.575
cc_527 N_A_110_115#_c_467_n N_A_1084_115#_c_1708_n 0.0119742f $X=8.715 $Y=1.22
+ $X2=7.685 $Y2=1.43
cc_528 N_A_110_115#_c_467_n N_A_1084_115#_c_1712_n 0.00328689f $X=8.715 $Y=1.22
+ $X2=7.685 $Y2=1.51
cc_529 N_A_110_115#_c_467_n N_A_1084_115#_c_1715_n 0.00616681f $X=8.715 $Y=1.22
+ $X2=5.065 $Y2=1.59
cc_530 N_A_110_115#_c_467_n N_A_1084_115#_c_1740_n 0.0536303f $X=8.715 $Y=1.22
+ $X2=5.475 $Y2=1.17
cc_531 N_A_110_115#_c_467_n N_A_1084_115#_c_1741_n 0.0129425f $X=8.715 $Y=1.22
+ $X2=5.15 $Y2=1.17
cc_532 N_A_110_115#_c_467_n N_A_1084_115#_c_1719_n 0.00241187f $X=8.715 $Y=1.22
+ $X2=7.595 $Y2=1.59
cc_533 N_A_110_115#_c_467_n N_A_1084_115#_c_1721_n 0.186671f $X=8.715 $Y=1.22
+ $X2=7.45 $Y2=1.59
cc_534 N_A_110_115#_c_467_n N_A_1084_115#_c_1724_n 0.0252354f $X=8.715 $Y=1.22
+ $X2=5.21 $Y2=1.59
cc_535 N_A_110_115#_c_467_n N_A_1084_115#_c_1725_n 0.0265552f $X=8.715 $Y=1.22
+ $X2=7.595 $Y2=1.59
cc_536 N_A_110_115#_c_441_n N_QN_c_1869_n 0.00557054f $X=8.535 $Y=1.205 $X2=9.28
+ $Y2=0.865
cc_537 N_A_110_115#_c_450_n N_QN_c_1869_n 0.0021703f $X=8.8 $Y=1.37 $X2=9.28
+ $Y2=0.865
cc_538 N_A_110_115#_c_465_n N_QN_c_1869_n 0.0193918f $X=8.86 $Y=1.22 $X2=9.28
+ $Y2=0.865
cc_539 N_A_110_115#_c_481_n N_QN_c_1869_n 0.00684422f $X=8.86 $Y=1.22 $X2=9.28
+ $Y2=0.865
cc_540 N_A_110_115#_c_446_n N_QN_c_1876_n 0.00202688f $X=8.8 $Y=2.345 $X2=9.365
+ $Y2=1.59
cc_541 N_A_110_115#_c_450_n N_QN_c_1876_n 8.42768e-19 $X=8.8 $Y=1.37 $X2=9.365
+ $Y2=1.59
cc_542 N_A_110_115#_c_452_n N_QN_c_1878_n 0.00115295f $X=8.545 $Y=2.49 $X2=9.365
+ $Y2=2.505
cc_543 N_A_110_115#_c_467_n A_400_115# 0.0100396f $X=8.715 $Y=1.22 $X2=2
+ $Y2=0.575
cc_544 N_A_110_115#_c_467_n A_662_115# 0.00911585f $X=8.715 $Y=1.22 $X2=3.31
+ $Y2=0.575
cc_545 N_A_110_115#_c_467_n A_854_115# 0.0100396f $X=8.715 $Y=1.22 $X2=4.27
+ $Y2=0.575
cc_546 N_A_110_115#_c_467_n A_1012_115# 0.00106636f $X=8.715 $Y=1.22 $X2=5.06
+ $Y2=0.575
cc_547 N_A_110_115#_c_467_n A_1204_115# 0.00917995f $X=8.715 $Y=1.22 $X2=6.02
+ $Y2=0.575
cc_548 N_A_110_115#_c_467_n A_1552_115# 0.0106361f $X=8.715 $Y=1.22 $X2=7.76
+ $Y2=0.575
cc_549 N_SN_M1011_g N_A_432_468#_M1000_g 0.103292f $X=1.925 $Y=0.945 $X2=2.285
+ $Y2=0.945
cc_550 N_SN_c_654_n N_A_432_468#_M1000_g 0.00875708f $X=1.855 $Y=2.11 $X2=2.285
+ $Y2=0.945
cc_551 N_SN_c_656_n N_A_432_468#_M1000_g 3.95753e-19 $X=1.71 $Y=2.7 $X2=2.285
+ $Y2=0.945
cc_552 N_SN_c_658_n N_A_432_468#_M1000_g 4.68111e-19 $X=1.71 $Y=2.11 $X2=2.285
+ $Y2=0.945
cc_553 N_SN_M1010_g N_A_432_468#_M1012_g 0.0530483f $X=1.855 $Y=3.825 $X2=2.285
+ $Y2=3.825
cc_554 N_SN_c_656_n N_A_432_468#_M1012_g 3.16831e-19 $X=1.71 $Y=2.7 $X2=2.285
+ $Y2=3.825
cc_555 N_SN_c_660_n N_A_432_468#_M1012_g 7.19848e-19 $X=7.79 $Y=2.7 $X2=2.285
+ $Y2=3.825
cc_556 N_SN_M1010_g N_A_432_468#_c_821_n 0.0179454f $X=1.855 $Y=3.825 $X2=2.295
+ $Y2=2.505
cc_557 N_SN_c_656_n N_A_432_468#_c_821_n 9.94587e-19 $X=1.71 $Y=2.7 $X2=2.295
+ $Y2=2.505
cc_558 N_SN_c_660_n N_A_432_468#_c_821_n 0.00593089f $X=7.79 $Y=2.7 $X2=2.295
+ $Y2=2.505
cc_559 N_SN_c_644_n N_A_432_468#_c_822_n 0.00268092f $X=1.89 $Y=1.625 $X2=2.295
+ $Y2=2.505
cc_560 N_SN_c_654_n N_A_432_468#_c_822_n 0.00272367f $X=1.855 $Y=2.11 $X2=2.295
+ $Y2=2.505
cc_561 N_SN_c_656_n N_A_432_468#_c_822_n 0.0170473f $X=1.71 $Y=2.7 $X2=2.295
+ $Y2=2.505
cc_562 N_SN_c_658_n N_A_432_468#_c_822_n 0.00704932f $X=1.71 $Y=2.11 $X2=2.295
+ $Y2=2.505
cc_563 N_SN_c_660_n N_A_432_468#_c_822_n 0.0236889f $X=7.79 $Y=2.7 $X2=2.295
+ $Y2=2.505
cc_564 N_SN_c_661_n N_A_432_468#_c_822_n 0.00164393f $X=1.855 $Y=2.7 $X2=2.295
+ $Y2=2.505
cc_565 N_SN_M1011_g N_A_432_468#_c_826_n 6.84827e-19 $X=1.925 $Y=0.945 $X2=2.38
+ $Y2=1.505
cc_566 N_SN_c_660_n N_A_432_468#_c_838_n 0.0775662f $X=7.79 $Y=2.7 $X2=3.725
+ $Y2=2.925
cc_567 N_SN_M1010_g N_A_432_468#_c_868_n 0.00105594f $X=1.855 $Y=3.825 $X2=2.38
+ $Y2=2.925
cc_568 N_SN_c_660_n N_D_M1014_g 0.00799543f $X=7.79 $Y=2.7 $X2=3.235 $Y2=3.825
cc_569 N_SN_c_660_n N_D_c_912_n 7.07415e-19 $X=7.79 $Y=2.7 $X2=3.295 $Y2=1.96
cc_570 N_SN_c_660_n N_D_c_913_n 0.00333216f $X=7.79 $Y=2.7 $X2=3.295 $Y2=1.96
cc_571 N_SN_c_660_n D 0.0134431f $X=7.79 $Y=2.7 $X2=3.295 $Y2=1.96
cc_572 N_SN_c_660_n N_CK_M1005_g 0.00294331f $X=7.79 $Y=2.7 $X2=3.595 $Y2=3.825
cc_573 N_SN_c_660_n N_CK_M1027_g 0.00796817f $X=7.79 $Y=2.7 $X2=5.945 $Y2=3.825
cc_574 N_SN_c_660_n N_CK_c_946_n 0.00448328f $X=7.79 $Y=2.7 $X2=6.735 $Y2=2.67
cc_575 N_SN_c_660_n N_CK_M1020_g 0.00909285f $X=7.79 $Y=2.7 $X2=6.735 $Y2=3.825
cc_576 N_SN_c_660_n N_CK_c_948_n 0.00264508f $X=7.79 $Y=2.7 $X2=3.655 $Y2=2.505
cc_577 N_SN_c_660_n N_CK_c_957_n 0.00264508f $X=7.79 $Y=2.7 $X2=5.885 $Y2=2.505
cc_578 N_SN_c_660_n N_CK_c_964_n 0.003555f $X=7.79 $Y=2.7 $X2=4.05 $Y2=2.33
cc_579 N_SN_c_660_n N_CK_c_967_n 0.00141703f $X=7.79 $Y=2.7 $X2=5.8 $Y2=2.33
cc_580 N_SN_c_660_n N_CK_c_968_n 9.71861e-19 $X=7.79 $Y=2.7 $X2=5.49 $Y2=2.33
cc_581 N_SN_c_660_n N_CK_c_969_n 0.00700078f $X=7.79 $Y=2.7 $X2=6.88 $Y2=2.33
cc_582 N_SN_c_660_n N_CK_c_970_n 0.00732128f $X=7.79 $Y=2.7 $X2=3.655 $Y2=2.33
cc_583 N_SN_c_660_n N_CK_c_971_n 0.00860578f $X=7.79 $Y=2.7 $X2=5.885 $Y2=2.33
cc_584 N_SN_c_660_n N_CK_c_972_n 0.15926f $X=7.79 $Y=2.7 $X2=5.74 $Y2=2.33
cc_585 N_SN_c_660_n N_CK_c_973_n 0.0251654f $X=7.79 $Y=2.7 $X2=3.8 $Y2=2.33
cc_586 N_SN_c_660_n N_CK_c_974_n 0.0598286f $X=7.79 $Y=2.7 $X2=6.735 $Y2=2.33
cc_587 N_SN_c_660_n N_CK_c_975_n 0.0251663f $X=7.79 $Y=2.7 $X2=6.03 $Y2=2.33
cc_588 N_SN_c_660_n CK 0.025144f $X=7.79 $Y=2.7 $X2=6.88 $Y2=2.33
cc_589 N_SN_c_660_n N_A_217_565#_M1030_g 0.00827407f $X=7.79 $Y=2.7 $X2=4.555
+ $Y2=3.825
cc_590 N_SN_c_660_n N_A_217_565#_c_1186_n 0.00177706f $X=7.79 $Y=2.7 $X2=4.91
+ $Y2=2.505
cc_591 N_SN_c_660_n N_A_217_565#_c_1187_n 0.00157006f $X=7.79 $Y=2.7 $X2=4.63
+ $Y2=2.505
cc_592 N_SN_c_660_n N_A_217_565#_M1032_g 0.00382698f $X=7.79 $Y=2.7 $X2=4.985
+ $Y2=3.825
cc_593 N_SN_c_645_n N_A_217_565#_c_1192_n 5.25241e-19 $X=1.89 $Y=1.945 $X2=1.21
+ $Y2=3.545
cc_594 N_SN_M1010_g N_A_217_565#_c_1192_n 3.2027e-19 $X=1.855 $Y=3.825 $X2=1.21
+ $Y2=3.545
cc_595 N_SN_c_654_n N_A_217_565#_c_1192_n 9.48304e-19 $X=1.855 $Y=2.11 $X2=1.21
+ $Y2=3.545
cc_596 N_SN_c_656_n N_A_217_565#_c_1192_n 0.0231905f $X=1.71 $Y=2.7 $X2=1.21
+ $Y2=3.545
cc_597 N_SN_c_658_n N_A_217_565#_c_1192_n 0.00963813f $X=1.71 $Y=2.11 $X2=1.21
+ $Y2=3.545
cc_598 N_SN_c_661_n N_A_217_565#_c_1192_n 0.00754015f $X=1.855 $Y=2.7 $X2=1.21
+ $Y2=3.545
cc_599 N_SN_c_645_n N_A_217_565#_c_1193_n 0.0055412f $X=1.89 $Y=1.945 $X2=1.625
+ $Y2=1.76
cc_600 N_SN_c_654_n N_A_217_565#_c_1193_n 0.00517882f $X=1.855 $Y=2.11 $X2=1.625
+ $Y2=1.76
cc_601 N_SN_c_658_n N_A_217_565#_c_1193_n 0.0186534f $X=1.71 $Y=2.11 $X2=1.625
+ $Y2=1.76
cc_602 N_SN_c_644_n N_A_217_565#_c_1195_n 0.00283874f $X=1.89 $Y=1.625 $X2=1.71
+ $Y2=0.865
cc_603 N_SN_c_645_n N_A_217_565#_c_1195_n 0.00108565f $X=1.89 $Y=1.945 $X2=1.71
+ $Y2=0.865
cc_604 N_SN_M1011_g N_A_217_565#_c_1195_n 0.0067599f $X=1.925 $Y=0.945 $X2=1.71
+ $Y2=0.865
cc_605 N_SN_c_660_n N_A_217_565#_c_1198_n 0.00880485f $X=7.79 $Y=2.7 $X2=4.725
+ $Y2=2.505
cc_606 N_SN_c_644_n N_A_217_565#_c_1201_n 0.00106358f $X=1.89 $Y=1.625 $X2=4.49
+ $Y2=1.59
cc_607 N_SN_c_645_n N_A_217_565#_c_1201_n 0.00565746f $X=1.89 $Y=1.945 $X2=4.49
+ $Y2=1.59
cc_608 N_SN_M1011_g N_A_217_565#_c_1201_n 0.00153565f $X=1.925 $Y=0.945 $X2=4.49
+ $Y2=1.59
cc_609 N_SN_c_658_n N_A_217_565#_c_1201_n 5.85585e-19 $X=1.71 $Y=2.11 $X2=4.49
+ $Y2=1.59
cc_610 N_SN_c_644_n N_A_217_565#_c_1202_n 4.80352e-19 $X=1.89 $Y=1.625 $X2=1.855
+ $Y2=1.59
cc_611 N_SN_c_645_n N_A_217_565#_c_1202_n 9.81257e-19 $X=1.89 $Y=1.945 $X2=1.855
+ $Y2=1.59
cc_612 N_SN_M1011_g N_A_217_565#_c_1202_n 5.70836e-19 $X=1.925 $Y=0.945
+ $X2=1.855 $Y2=1.59
cc_613 N_SN_c_658_n N_A_217_565#_c_1202_n 0.00329414f $X=1.71 $Y=2.11 $X2=1.855
+ $Y2=1.59
cc_614 N_SN_c_660_n N_A_704_89#_M1035_g 0.0108138f $X=7.79 $Y=2.7 $X2=4.195
+ $Y2=3.825
cc_615 N_SN_c_660_n N_A_704_89#_M1031_g 0.00578896f $X=7.79 $Y=2.7 $X2=5.345
+ $Y2=3.825
cc_616 N_SN_c_657_n N_A_704_89#_c_1370_n 0.00228032f $X=7.935 $Y=2.7 $X2=7.22
+ $Y2=2.84
cc_617 N_SN_c_660_n N_A_704_89#_c_1370_n 0.0163748f $X=7.79 $Y=2.7 $X2=7.22
+ $Y2=2.84
cc_618 SN N_A_704_89#_c_1370_n 0.00108239f $X=7.935 $Y=2.7 $X2=7.22 $Y2=2.84
cc_619 N_SN_c_660_n N_A_704_89#_c_1372_n 0.00232295f $X=7.79 $Y=2.7 $X2=7.22
+ $Y2=1.93
cc_620 N_SN_c_660_n N_A_704_89#_c_1383_n 0.0135346f $X=7.79 $Y=2.7 $X2=7.22
+ $Y2=2.925
cc_621 N_SN_c_660_n N_A_1246_89#_M1015_g 0.0105543f $X=7.79 $Y=2.7 $X2=6.305
+ $Y2=3.825
cc_622 N_SN_M1001_g N_A_1246_89#_c_1552_n 0.0089462f $X=8.045 $Y=0.945 $X2=8.26
+ $Y2=0.865
cc_623 N_SN_M1007_g N_A_1246_89#_c_1555_n 8.82733e-19 $X=8.115 $Y=3.825 $X2=8.76
+ $Y2=3.545
cc_624 N_SN_c_655_n N_A_1246_89#_c_1555_n 0.0019272f $X=8.025 $Y=1.995 $X2=8.76
+ $Y2=3.545
cc_625 N_SN_c_657_n N_A_1246_89#_c_1555_n 0.0144281f $X=7.935 $Y=2.7 $X2=8.76
+ $Y2=3.545
cc_626 N_SN_c_659_n N_A_1246_89#_c_1555_n 0.00492795f $X=8.025 $Y=1.995 $X2=8.76
+ $Y2=3.545
cc_627 SN N_A_1246_89#_c_1555_n 0.00496818f $X=7.935 $Y=2.7 $X2=8.76 $Y2=3.545
cc_628 N_SN_M1001_g N_A_1246_89#_c_1556_n 0.00483036f $X=8.045 $Y=0.945
+ $X2=8.845 $Y2=1.93
cc_629 N_SN_c_655_n N_A_1246_89#_c_1556_n 0.0026134f $X=8.025 $Y=1.995 $X2=8.845
+ $Y2=1.93
cc_630 N_SN_c_659_n N_A_1246_89#_c_1556_n 0.00832911f $X=8.025 $Y=1.995
+ $X2=8.845 $Y2=1.93
cc_631 N_SN_c_655_n N_A_1246_89#_c_1558_n 0.00614421f $X=8.025 $Y=1.995
+ $X2=9.235 $Y2=1.93
cc_632 N_SN_c_657_n N_A_1246_89#_c_1558_n 9.11589e-19 $X=7.935 $Y=2.7 $X2=9.235
+ $Y2=1.93
cc_633 N_SN_c_659_n N_A_1246_89#_c_1558_n 0.020493f $X=8.025 $Y=1.995 $X2=9.235
+ $Y2=1.93
cc_634 N_SN_M1001_g N_A_1084_115#_c_1707_n 0.00627778f $X=8.045 $Y=0.945
+ $X2=7.505 $Y2=2.37
cc_635 N_SN_M1007_g N_A_1084_115#_c_1707_n 0.00402616f $X=8.115 $Y=3.825
+ $X2=7.505 $Y2=2.37
cc_636 N_SN_c_655_n N_A_1084_115#_c_1707_n 0.0138276f $X=8.025 $Y=1.995
+ $X2=7.505 $Y2=2.37
cc_637 N_SN_c_657_n N_A_1084_115#_c_1707_n 5.97554e-19 $X=7.935 $Y=2.7 $X2=7.505
+ $Y2=2.37
cc_638 N_SN_c_659_n N_A_1084_115#_c_1707_n 6.33368e-19 $X=8.025 $Y=1.995
+ $X2=7.505 $Y2=2.37
cc_639 N_SN_M1001_g N_A_1084_115#_c_1708_n 0.0702195f $X=8.045 $Y=0.945
+ $X2=7.685 $Y2=1.43
cc_640 N_SN_c_660_n N_A_1084_115#_M1021_g 0.00486063f $X=7.79 $Y=2.7 $X2=7.685
+ $Y2=3.825
cc_641 SN N_A_1084_115#_M1021_g 5.06369e-19 $X=7.935 $Y=2.7 $X2=7.685 $Y2=3.825
cc_642 N_SN_M1007_g N_A_1084_115#_c_1714_n 0.0670991f $X=8.115 $Y=3.825
+ $X2=7.685 $Y2=2.505
cc_643 N_SN_c_657_n N_A_1084_115#_c_1714_n 0.00312462f $X=7.935 $Y=2.7 $X2=7.685
+ $Y2=2.505
cc_644 N_SN_c_660_n N_A_1084_115#_c_1714_n 0.00760041f $X=7.79 $Y=2.7 $X2=7.685
+ $Y2=2.505
cc_645 SN N_A_1084_115#_c_1714_n 5.28053e-19 $X=7.935 $Y=2.7 $X2=7.685 $Y2=2.505
cc_646 N_SN_c_660_n N_A_1084_115#_c_1715_n 0.0225202f $X=7.79 $Y=2.7 $X2=5.065
+ $Y2=1.59
cc_647 N_SN_c_660_n N_A_1084_115#_c_1759_n 0.0256731f $X=7.79 $Y=2.7 $X2=5.475
+ $Y2=2.925
cc_648 N_SN_M1001_g N_A_1084_115#_c_1719_n 0.00316718f $X=8.045 $Y=0.945
+ $X2=7.595 $Y2=1.59
cc_649 N_SN_c_655_n N_A_1084_115#_c_1719_n 0.00203974f $X=8.025 $Y=1.995
+ $X2=7.595 $Y2=1.59
cc_650 N_SN_c_657_n N_A_1084_115#_c_1719_n 0.0367765f $X=7.935 $Y=2.7 $X2=7.595
+ $Y2=1.59
cc_651 N_SN_c_659_n N_A_1084_115#_c_1719_n 0.0189565f $X=8.025 $Y=1.995
+ $X2=7.595 $Y2=1.59
cc_652 N_SN_c_660_n N_A_1084_115#_c_1719_n 0.0136826f $X=7.79 $Y=2.7 $X2=7.595
+ $Y2=1.59
cc_653 SN N_A_1084_115#_c_1719_n 9.02875e-19 $X=7.935 $Y=2.7 $X2=7.595 $Y2=1.59
cc_654 N_SN_M1001_g N_A_1084_115#_c_1725_n 0.00271237f $X=8.045 $Y=0.945
+ $X2=7.595 $Y2=1.59
cc_655 N_SN_M1010_g N_A_300_565#_c_1949_n 0.0147996f $X=1.855 $Y=3.825 $X2=2.415
+ $Y2=3.37
cc_656 N_SN_c_656_n N_A_300_565#_c_1949_n 8.68455e-19 $X=1.71 $Y=2.7 $X2=2.415
+ $Y2=3.37
cc_657 N_SN_c_660_n N_A_300_565#_c_1949_n 0.0122781f $X=7.79 $Y=2.7 $X2=2.415
+ $Y2=3.37
cc_658 N_SN_c_661_n N_A_300_565#_c_1949_n 0.00326201f $X=1.855 $Y=2.7 $X2=2.415
+ $Y2=3.37
cc_659 N_SN_c_656_n N_A_300_565#_c_1960_n 0.00230057f $X=1.71 $Y=2.7 $X2=1.725
+ $Y2=3.37
cc_660 N_SN_c_661_n N_A_300_565#_c_1960_n 0.00491504f $X=1.855 $Y=2.7 $X2=1.725
+ $Y2=3.37
cc_661 N_SN_M1007_g N_A_1469_565#_c_1973_n 0.0172185f $X=8.115 $Y=3.825
+ $X2=8.245 $Y2=3.37
cc_662 N_SN_c_657_n N_A_1469_565#_c_1973_n 0.0032182f $X=7.935 $Y=2.7 $X2=8.245
+ $Y2=3.37
cc_663 N_SN_c_660_n N_A_1469_565#_c_1973_n 0.0055835f $X=7.79 $Y=2.7 $X2=8.245
+ $Y2=3.37
cc_664 SN N_A_1469_565#_c_1973_n 0.00793147f $X=7.935 $Y=2.7 $X2=8.245 $Y2=3.37
cc_665 N_SN_c_660_n N_A_1469_565#_c_1982_n 0.00594846f $X=7.79 $Y=2.7 $X2=7.555
+ $Y2=3.37
cc_666 N_A_432_468#_c_823_n N_D_M1002_g 0.0123125f $X=3.71 $Y=1.505 $X2=3.235
+ $Y2=0.945
cc_667 N_A_432_468#_c_838_n N_D_M1014_g 0.0167212f $X=3.725 $Y=2.925 $X2=3.235
+ $Y2=3.825
cc_668 N_A_432_468#_c_823_n N_D_c_912_n 0.00207628f $X=3.71 $Y=1.505 $X2=3.295
+ $Y2=1.96
cc_669 N_A_432_468#_c_823_n N_D_c_913_n 0.0086486f $X=3.71 $Y=1.505 $X2=3.295
+ $Y2=1.96
cc_670 N_A_432_468#_c_823_n D 0.00200799f $X=3.71 $Y=1.505 $X2=3.295 $Y2=1.96
cc_671 N_A_432_468#_c_838_n N_CK_M1005_g 0.0150535f $X=3.725 $Y=2.925 $X2=3.595
+ $Y2=3.825
cc_672 N_A_432_468#_c_838_n N_CK_c_948_n 0.00123101f $X=3.725 $Y=2.925 $X2=3.655
+ $Y2=2.505
cc_673 N_A_432_468#_c_823_n N_CK_c_949_n 9.45214e-19 $X=3.71 $Y=1.505 $X2=4.135
+ $Y2=1.59
cc_674 N_A_432_468#_c_849_n N_CK_c_949_n 0.00168646f $X=3.887 $Y=1.155 $X2=4.135
+ $Y2=1.59
cc_675 N_A_432_468#_c_827_n N_CK_c_950_n 0.00464203f $X=3.795 $Y=1.42 $X2=4.135
+ $Y2=1.425
cc_676 N_A_432_468#_c_849_n N_CK_c_950_n 0.00381867f $X=3.887 $Y=1.155 $X2=4.135
+ $Y2=1.425
cc_677 N_A_432_468#_c_823_n N_CK_c_964_n 0.0019742f $X=3.71 $Y=1.505 $X2=4.05
+ $Y2=2.33
cc_678 N_A_432_468#_c_838_n N_CK_c_964_n 0.00786738f $X=3.725 $Y=2.925 $X2=4.05
+ $Y2=2.33
cc_679 N_A_432_468#_c_823_n N_CK_c_965_n 0.012316f $X=3.71 $Y=1.505 $X2=4.135
+ $Y2=1.59
cc_680 N_A_432_468#_c_849_n N_CK_c_965_n 5.27251e-19 $X=3.887 $Y=1.155 $X2=4.135
+ $Y2=1.59
cc_681 N_A_432_468#_c_823_n N_CK_c_970_n 0.00224444f $X=3.71 $Y=1.505 $X2=3.655
+ $Y2=2.33
cc_682 N_A_432_468#_c_838_n N_CK_c_970_n 0.0085861f $X=3.725 $Y=2.925 $X2=3.655
+ $Y2=2.33
cc_683 N_A_432_468#_M1000_g N_A_217_565#_c_1193_n 4.08059e-19 $X=2.285 $Y=0.945
+ $X2=1.625 $Y2=1.76
cc_684 N_A_432_468#_c_822_n N_A_217_565#_c_1193_n 0.00578447f $X=2.295 $Y=2.505
+ $X2=1.625 $Y2=1.76
cc_685 N_A_432_468#_M1000_g N_A_217_565#_c_1195_n 3.32429e-19 $X=2.285 $Y=0.945
+ $X2=1.71 $Y2=0.865
cc_686 N_A_432_468#_c_822_n N_A_217_565#_c_1195_n 0.00179268f $X=2.295 $Y=2.505
+ $X2=1.71 $Y2=0.865
cc_687 N_A_432_468#_c_826_n N_A_217_565#_c_1195_n 0.00488587f $X=2.38 $Y=1.505
+ $X2=1.71 $Y2=0.865
cc_688 N_A_432_468#_M1000_g N_A_217_565#_c_1201_n 8.36391e-19 $X=2.285 $Y=0.945
+ $X2=4.49 $Y2=1.59
cc_689 N_A_432_468#_c_822_n N_A_217_565#_c_1201_n 0.0151086f $X=2.295 $Y=2.505
+ $X2=4.49 $Y2=1.59
cc_690 N_A_432_468#_c_823_n N_A_217_565#_c_1201_n 0.0578899f $X=3.71 $Y=1.505
+ $X2=4.49 $Y2=1.59
cc_691 N_A_432_468#_c_826_n N_A_217_565#_c_1201_n 0.00475107f $X=2.38 $Y=1.505
+ $X2=4.49 $Y2=1.59
cc_692 N_A_432_468#_c_849_n N_A_217_565#_c_1201_n 8.67164e-19 $X=3.887 $Y=1.155
+ $X2=4.49 $Y2=1.59
cc_693 N_A_432_468#_c_822_n N_A_217_565#_c_1202_n 6.43558e-19 $X=2.295 $Y=2.505
+ $X2=1.855 $Y2=1.59
cc_694 N_A_432_468#_c_826_n N_A_217_565#_c_1202_n 6.84883e-19 $X=2.38 $Y=1.505
+ $X2=1.855 $Y2=1.59
cc_695 N_A_432_468#_c_823_n N_A_704_89#_c_1344_n 0.0022787f $X=3.71 $Y=1.505
+ $X2=3.595 $Y2=1.425
cc_696 N_A_432_468#_c_849_n N_A_704_89#_c_1344_n 0.0060945f $X=3.887 $Y=1.155
+ $X2=3.595 $Y2=1.425
cc_697 N_A_432_468#_c_823_n N_A_704_89#_c_1347_n 0.00324141f $X=3.71 $Y=1.505
+ $X2=3.715 $Y2=1.965
cc_698 N_A_432_468#_c_823_n N_A_704_89#_c_1355_n 0.00993431f $X=3.71 $Y=1.505
+ $X2=3.715 $Y2=1.5
cc_699 N_A_432_468#_c_838_n N_A_300_565#_M1012_d 0.00690809f $X=3.725 $Y=2.925
+ $X2=2.36 $Y2=2.825
cc_700 N_A_432_468#_M1012_g N_A_300_565#_c_1949_n 0.0146873f $X=2.285 $Y=3.825
+ $X2=2.415 $Y2=3.37
cc_701 N_A_432_468#_c_838_n N_A_300_565#_c_1949_n 0.00856071f $X=3.725 $Y=2.925
+ $X2=2.415 $Y2=3.37
cc_702 N_A_432_468#_c_868_n N_A_300_565#_c_1949_n 0.0070523f $X=2.38 $Y=2.925
+ $X2=2.415 $Y2=3.37
cc_703 N_A_432_468#_c_838_n A_662_565# 0.00481059f $X=3.725 $Y=2.925 $X2=3.31
+ $Y2=2.825
cc_704 N_D_M1014_g N_CK_c_948_n 0.158539f $X=3.235 $Y=3.825 $X2=3.655 $Y2=2.505
cc_705 N_D_c_912_n N_CK_c_965_n 2.89615e-19 $X=3.295 $Y=1.96 $X2=4.135 $Y2=1.59
cc_706 N_D_c_913_n N_CK_c_965_n 0.00478177f $X=3.295 $Y=1.96 $X2=4.135 $Y2=1.59
cc_707 D N_CK_c_965_n 0.00551577f $X=3.295 $Y=1.96 $X2=4.135 $Y2=1.59
cc_708 N_D_M1014_g N_CK_c_970_n 0.00512934f $X=3.235 $Y=3.825 $X2=3.655 $Y2=2.33
cc_709 N_D_M1014_g N_CK_c_973_n 0.00515433f $X=3.235 $Y=3.825 $X2=3.8 $Y2=2.33
cc_710 D N_CK_c_973_n 0.00375733f $X=3.295 $Y=1.96 $X2=3.8 $Y2=2.33
cc_711 N_D_M1002_g N_A_217_565#_c_1201_n 0.00303372f $X=3.235 $Y=0.945 $X2=4.49
+ $Y2=1.59
cc_712 N_D_c_912_n N_A_217_565#_c_1201_n 7.9412e-19 $X=3.295 $Y=1.96 $X2=4.49
+ $Y2=1.59
cc_713 N_D_c_913_n N_A_217_565#_c_1201_n 0.00111625f $X=3.295 $Y=1.96 $X2=4.49
+ $Y2=1.59
cc_714 D N_A_217_565#_c_1201_n 0.0353362f $X=3.295 $Y=1.96 $X2=4.49 $Y2=1.59
cc_715 N_D_M1002_g N_A_704_89#_c_1344_n 0.0695166f $X=3.235 $Y=0.945 $X2=3.595
+ $Y2=1.425
cc_716 N_D_M1002_g N_A_704_89#_c_1347_n 0.00932846f $X=3.235 $Y=0.945 $X2=3.715
+ $Y2=1.965
cc_717 N_D_c_912_n N_A_704_89#_c_1347_n 0.0210215f $X=3.295 $Y=1.96 $X2=3.715
+ $Y2=1.965
cc_718 N_D_c_913_n N_A_704_89#_c_1347_n 0.00164409f $X=3.295 $Y=1.96 $X2=3.715
+ $Y2=1.965
cc_719 D N_A_704_89#_c_1347_n 0.00342011f $X=3.295 $Y=1.96 $X2=3.715 $Y2=1.965
cc_720 D N_A_704_89#_c_1349_n 4.62757e-19 $X=3.295 $Y=1.96 $X2=3.79 $Y2=2.04
cc_721 N_CK_c_950_n N_A_217_565#_M1022_g 0.0406519f $X=4.135 $Y=1.425 $X2=4.555
+ $Y2=0.945
cc_722 N_CK_c_965_n N_A_217_565#_M1022_g 0.00109079f $X=4.135 $Y=1.59 $X2=4.555
+ $Y2=0.945
cc_723 N_CK_c_953_n N_A_217_565#_c_1183_n 0.0396058f $X=5.405 $Y=1.59 $X2=4.91
+ $Y2=1.59
cc_724 N_CK_c_949_n N_A_217_565#_c_1185_n 0.0406519f $X=4.135 $Y=1.59 $X2=4.63
+ $Y2=1.59
cc_725 N_CK_c_972_n N_A_217_565#_c_1186_n 0.00203319f $X=5.74 $Y=2.33 $X2=4.91
+ $Y2=2.505
cc_726 N_CK_c_972_n N_A_217_565#_c_1187_n 0.00203351f $X=5.74 $Y=2.33 $X2=4.63
+ $Y2=2.505
cc_727 N_CK_c_954_n N_A_217_565#_M1028_g 0.0396058f $X=5.405 $Y=1.425 $X2=4.985
+ $Y2=0.945
cc_728 N_CK_c_966_n N_A_217_565#_M1028_g 3.67139e-19 $X=5.405 $Y=1.59 $X2=4.985
+ $Y2=0.945
cc_729 N_CK_c_949_n N_A_217_565#_c_1198_n 7.30049e-19 $X=4.135 $Y=1.59 $X2=4.725
+ $Y2=2.505
cc_730 N_CK_c_964_n N_A_217_565#_c_1198_n 0.00401809f $X=4.05 $Y=2.33 $X2=4.725
+ $Y2=2.505
cc_731 N_CK_c_965_n N_A_217_565#_c_1198_n 0.0203851f $X=4.135 $Y=1.59 $X2=4.725
+ $Y2=2.505
cc_732 N_CK_c_972_n N_A_217_565#_c_1198_n 0.0154699f $X=5.74 $Y=2.33 $X2=4.725
+ $Y2=2.505
cc_733 N_CK_c_949_n N_A_217_565#_c_1199_n 7.18106e-19 $X=4.135 $Y=1.59 $X2=4.725
+ $Y2=1.59
cc_734 N_CK_c_965_n N_A_217_565#_c_1199_n 0.00742068f $X=4.135 $Y=1.59 $X2=4.725
+ $Y2=1.59
cc_735 N_CK_c_972_n N_A_217_565#_c_1199_n 0.00102309f $X=5.74 $Y=2.33 $X2=4.725
+ $Y2=1.59
cc_736 N_CK_c_949_n N_A_217_565#_c_1201_n 0.00383172f $X=4.135 $Y=1.59 $X2=4.49
+ $Y2=1.59
cc_737 N_CK_c_964_n N_A_217_565#_c_1201_n 0.00443421f $X=4.05 $Y=2.33 $X2=4.49
+ $Y2=1.59
cc_738 N_CK_c_965_n N_A_217_565#_c_1201_n 0.0149977f $X=4.135 $Y=1.59 $X2=4.49
+ $Y2=1.59
cc_739 N_CK_c_970_n N_A_217_565#_c_1201_n 7.12046e-19 $X=3.655 $Y=2.33 $X2=4.49
+ $Y2=1.59
cc_740 N_CK_c_973_n N_A_217_565#_c_1201_n 0.0126164f $X=3.8 $Y=2.33 $X2=4.49
+ $Y2=1.59
cc_741 N_CK_c_949_n N_A_217_565#_c_1252_n 3.3031e-19 $X=4.135 $Y=1.59 $X2=4.635
+ $Y2=1.59
cc_742 N_CK_c_965_n N_A_217_565#_c_1252_n 0.00143592f $X=4.135 $Y=1.59 $X2=4.635
+ $Y2=1.59
cc_743 N_CK_c_972_n N_A_217_565#_c_1252_n 0.0129652f $X=5.74 $Y=2.33 $X2=4.635
+ $Y2=1.59
cc_744 N_CK_c_950_n N_A_704_89#_c_1344_n 0.020867f $X=4.135 $Y=1.425 $X2=3.595
+ $Y2=1.425
cc_745 N_CK_c_965_n N_A_704_89#_c_1347_n 0.00613747f $X=4.135 $Y=1.59 $X2=3.715
+ $Y2=1.965
cc_746 N_CK_c_949_n N_A_704_89#_c_1348_n 0.0183603f $X=4.135 $Y=1.59 $X2=4.12
+ $Y2=2.04
cc_747 N_CK_c_965_n N_A_704_89#_c_1348_n 0.00630484f $X=4.135 $Y=1.59 $X2=4.12
+ $Y2=2.04
cc_748 N_CK_c_972_n N_A_704_89#_c_1348_n 0.00613485f $X=5.74 $Y=2.33 $X2=4.12
+ $Y2=2.04
cc_749 N_CK_c_948_n N_A_704_89#_c_1349_n 0.00904036f $X=3.655 $Y=2.505 $X2=3.79
+ $Y2=2.04
cc_750 N_CK_c_964_n N_A_704_89#_c_1349_n 0.00878348f $X=4.05 $Y=2.33 $X2=3.79
+ $Y2=2.04
cc_751 N_CK_c_970_n N_A_704_89#_c_1349_n 0.00109468f $X=3.655 $Y=2.33 $X2=3.79
+ $Y2=2.04
cc_752 N_CK_c_973_n N_A_704_89#_c_1349_n 0.00137501f $X=3.8 $Y=2.33 $X2=3.79
+ $Y2=2.04
cc_753 N_CK_M1005_g N_A_704_89#_M1035_g 0.0437214f $X=3.595 $Y=3.825 $X2=4.195
+ $Y2=3.825
cc_754 N_CK_c_948_n N_A_704_89#_M1035_g 0.0129692f $X=3.655 $Y=2.505 $X2=4.195
+ $Y2=3.825
cc_755 N_CK_c_964_n N_A_704_89#_M1035_g 0.0081071f $X=4.05 $Y=2.33 $X2=4.195
+ $Y2=3.825
cc_756 N_CK_c_965_n N_A_704_89#_M1035_g 0.00478024f $X=4.135 $Y=1.59 $X2=4.195
+ $Y2=3.825
cc_757 N_CK_c_970_n N_A_704_89#_M1035_g 0.00197555f $X=3.655 $Y=2.33 $X2=4.195
+ $Y2=3.825
cc_758 N_CK_c_972_n N_A_704_89#_M1035_g 0.00462358f $X=5.74 $Y=2.33 $X2=4.195
+ $Y2=3.825
cc_759 N_CK_c_973_n N_A_704_89#_M1035_g 4.2e-19 $X=3.8 $Y=2.33 $X2=4.195
+ $Y2=3.825
cc_760 N_CK_c_972_n N_A_704_89#_c_1351_n 0.00607908f $X=5.74 $Y=2.33 $X2=5.27
+ $Y2=2.04
cc_761 N_CK_M1027_g N_A_704_89#_M1031_g 0.0437279f $X=5.945 $Y=3.825 $X2=5.345
+ $Y2=3.825
cc_762 N_CK_c_957_n N_A_704_89#_M1031_g 0.0122143f $X=5.885 $Y=2.505 $X2=5.345
+ $Y2=3.825
cc_763 N_CK_c_966_n N_A_704_89#_M1031_g 0.00399495f $X=5.405 $Y=1.59 $X2=5.345
+ $Y2=3.825
cc_764 N_CK_c_968_n N_A_704_89#_M1031_g 0.00654233f $X=5.49 $Y=2.33 $X2=5.345
+ $Y2=3.825
cc_765 N_CK_c_971_n N_A_704_89#_M1031_g 0.00130061f $X=5.885 $Y=2.33 $X2=5.345
+ $Y2=3.825
cc_766 N_CK_c_972_n N_A_704_89#_M1031_g 0.00422185f $X=5.74 $Y=2.33 $X2=5.345
+ $Y2=3.825
cc_767 N_CK_c_975_n N_A_704_89#_M1031_g 4.2e-19 $X=6.03 $Y=2.33 $X2=5.345
+ $Y2=3.825
cc_768 N_CK_c_957_n N_A_704_89#_c_1353_n 0.00904036f $X=5.885 $Y=2.505 $X2=5.75
+ $Y2=2.04
cc_769 N_CK_c_966_n N_A_704_89#_c_1353_n 0.00909647f $X=5.405 $Y=1.59 $X2=5.75
+ $Y2=2.04
cc_770 N_CK_c_967_n N_A_704_89#_c_1353_n 0.00924811f $X=5.8 $Y=2.33 $X2=5.75
+ $Y2=2.04
cc_771 N_CK_c_971_n N_A_704_89#_c_1353_n 0.00102633f $X=5.885 $Y=2.33 $X2=5.75
+ $Y2=2.04
cc_772 N_CK_c_972_n N_A_704_89#_c_1353_n 0.00613485f $X=5.74 $Y=2.33 $X2=5.75
+ $Y2=2.04
cc_773 N_CK_c_975_n N_A_704_89#_c_1353_n 0.00137501f $X=6.03 $Y=2.33 $X2=5.75
+ $Y2=2.04
cc_774 N_CK_c_966_n N_A_704_89#_c_1354_n 0.00649764f $X=5.405 $Y=1.59 $X2=5.825
+ $Y2=1.965
cc_775 N_CK_c_949_n N_A_704_89#_c_1355_n 0.0216263f $X=4.135 $Y=1.59 $X2=3.715
+ $Y2=1.5
cc_776 N_CK_c_970_n N_A_704_89#_c_1355_n 2.45465e-19 $X=3.655 $Y=2.33 $X2=3.715
+ $Y2=1.5
cc_777 N_CK_c_965_n N_A_704_89#_c_1356_n 0.00568091f $X=4.135 $Y=1.59 $X2=4.195
+ $Y2=2.04
cc_778 N_CK_c_953_n N_A_704_89#_c_1357_n 0.0183603f $X=5.405 $Y=1.59 $X2=5.345
+ $Y2=2.04
cc_779 N_CK_c_966_n N_A_704_89#_c_1357_n 0.00436024f $X=5.405 $Y=1.59 $X2=5.345
+ $Y2=2.04
cc_780 N_CK_c_953_n N_A_704_89#_c_1358_n 0.0220721f $X=5.405 $Y=1.59 $X2=5.885
+ $Y2=1.59
cc_781 N_CK_c_957_n N_A_704_89#_c_1358_n 0.00227671f $X=5.885 $Y=2.505 $X2=5.885
+ $Y2=1.59
cc_782 N_CK_c_966_n N_A_704_89#_c_1358_n 0.00131283f $X=5.405 $Y=1.59 $X2=5.885
+ $Y2=1.59
cc_783 N_CK_c_971_n N_A_704_89#_c_1358_n 5.27321e-19 $X=5.885 $Y=2.33 $X2=5.885
+ $Y2=1.59
cc_784 N_CK_c_975_n N_A_704_89#_c_1358_n 8.78837e-19 $X=6.03 $Y=2.33 $X2=5.885
+ $Y2=1.59
cc_785 N_CK_c_954_n N_A_704_89#_c_1359_n 0.022472f $X=5.405 $Y=1.425 $X2=5.885
+ $Y2=1.425
cc_786 N_CK_c_947_n N_A_704_89#_c_1362_n 0.00592387f $X=6.79 $Y=2.34 $X2=6.865
+ $Y2=1.59
cc_787 N_CK_c_953_n N_A_704_89#_c_1362_n 8.05876e-19 $X=5.405 $Y=1.59 $X2=6.865
+ $Y2=1.59
cc_788 N_CK_c_957_n N_A_704_89#_c_1362_n 5.56676e-19 $X=5.885 $Y=2.505 $X2=6.865
+ $Y2=1.59
cc_789 N_CK_c_963_n N_A_704_89#_c_1362_n 0.00762848f $X=6.762 $Y=1.575 $X2=6.865
+ $Y2=1.59
cc_790 N_CK_c_966_n N_A_704_89#_c_1362_n 0.00853323f $X=5.405 $Y=1.59 $X2=6.865
+ $Y2=1.59
cc_791 N_CK_c_967_n N_A_704_89#_c_1362_n 0.00132011f $X=5.8 $Y=2.33 $X2=6.865
+ $Y2=1.59
cc_792 N_CK_c_969_n N_A_704_89#_c_1362_n 8.24249e-19 $X=6.88 $Y=2.33 $X2=6.865
+ $Y2=1.59
cc_793 N_CK_c_971_n N_A_704_89#_c_1362_n 0.00261697f $X=5.885 $Y=2.33 $X2=6.865
+ $Y2=1.59
cc_794 N_CK_c_972_n N_A_704_89#_c_1362_n 3.12599e-19 $X=5.74 $Y=2.33 $X2=6.865
+ $Y2=1.59
cc_795 N_CK_c_974_n N_A_704_89#_c_1362_n 0.00341454f $X=6.735 $Y=2.33 $X2=6.865
+ $Y2=1.59
cc_796 N_CK_c_975_n N_A_704_89#_c_1362_n 0.00221563f $X=6.03 $Y=2.33 $X2=6.865
+ $Y2=1.59
cc_797 N_CK_c_958_n N_A_704_89#_c_1364_n 0.0117675f $X=6.762 $Y=1.425 $X2=6.95
+ $Y2=0.865
cc_798 N_CK_c_963_n N_A_704_89#_c_1364_n 0.00243671f $X=6.762 $Y=1.575 $X2=6.95
+ $Y2=0.865
cc_799 N_CK_c_947_n N_A_704_89#_c_1369_n 0.00495963f $X=6.79 $Y=2.34 $X2=6.95
+ $Y2=1.845
cc_800 N_CK_c_946_n N_A_704_89#_c_1370_n 0.00262756f $X=6.735 $Y=2.67 $X2=7.22
+ $Y2=2.84
cc_801 N_CK_M1020_g N_A_704_89#_c_1370_n 0.00395773f $X=6.735 $Y=3.825 $X2=7.22
+ $Y2=2.84
cc_802 N_CK_c_947_n N_A_704_89#_c_1370_n 0.0049943f $X=6.79 $Y=2.34 $X2=7.22
+ $Y2=2.84
cc_803 N_CK_c_969_n N_A_704_89#_c_1370_n 0.0285927f $X=6.88 $Y=2.33 $X2=7.22
+ $Y2=2.84
cc_804 CK N_A_704_89#_c_1370_n 0.00851352f $X=6.88 $Y=2.33 $X2=7.22 $Y2=2.84
cc_805 N_CK_c_947_n N_A_704_89#_c_1371_n 0.00126782f $X=6.79 $Y=2.34 $X2=6.95
+ $Y2=1.59
cc_806 N_CK_c_963_n N_A_704_89#_c_1371_n 8.92648e-19 $X=6.762 $Y=1.575 $X2=6.95
+ $Y2=1.59
cc_807 N_CK_c_946_n N_A_704_89#_c_1372_n 0.001573f $X=6.735 $Y=2.67 $X2=7.22
+ $Y2=1.93
cc_808 N_CK_c_947_n N_A_704_89#_c_1372_n 0.00236123f $X=6.79 $Y=2.34 $X2=7.22
+ $Y2=1.93
cc_809 N_CK_c_969_n N_A_704_89#_c_1372_n 0.00528683f $X=6.88 $Y=2.33 $X2=7.22
+ $Y2=1.93
cc_810 CK N_A_704_89#_c_1372_n 8.7939e-19 $X=6.88 $Y=2.33 $X2=7.22 $Y2=1.93
cc_811 N_CK_c_946_n N_A_704_89#_c_1383_n 0.00233394f $X=6.735 $Y=2.67 $X2=7.22
+ $Y2=2.925
cc_812 N_CK_c_969_n N_A_704_89#_c_1383_n 0.00601935f $X=6.88 $Y=2.33 $X2=7.22
+ $Y2=2.925
cc_813 N_CK_c_947_n N_A_1246_89#_M1003_g 0.00697006f $X=6.79 $Y=2.34 $X2=6.305
+ $Y2=0.945
cc_814 N_CK_c_958_n N_A_1246_89#_M1003_g 0.0315481f $X=6.762 $Y=1.425 $X2=6.305
+ $Y2=0.945
cc_815 N_CK_c_946_n N_A_1246_89#_M1015_g 0.029689f $X=6.735 $Y=2.67 $X2=6.305
+ $Y2=3.825
cc_816 N_CK_c_947_n N_A_1246_89#_M1015_g 0.0175925f $X=6.79 $Y=2.34 $X2=6.305
+ $Y2=3.825
cc_817 N_CK_c_957_n N_A_1246_89#_M1015_g 0.157364f $X=5.885 $Y=2.505 $X2=6.305
+ $Y2=3.825
cc_818 N_CK_c_969_n N_A_1246_89#_M1015_g 0.00276527f $X=6.88 $Y=2.33 $X2=6.305
+ $Y2=3.825
cc_819 N_CK_c_971_n N_A_1246_89#_M1015_g 0.00472186f $X=5.885 $Y=2.33 $X2=6.305
+ $Y2=3.825
cc_820 N_CK_c_974_n N_A_1246_89#_M1015_g 0.00672311f $X=6.735 $Y=2.33 $X2=6.305
+ $Y2=3.825
cc_821 N_CK_c_975_n N_A_1246_89#_M1015_g 0.00113587f $X=6.03 $Y=2.33 $X2=6.305
+ $Y2=3.825
cc_822 CK N_A_1246_89#_M1015_g 3.05655e-19 $X=6.88 $Y=2.33 $X2=6.305 $Y2=3.825
cc_823 N_CK_c_947_n N_A_1246_89#_c_1540_n 0.0213817f $X=6.79 $Y=2.34 $X2=6.365
+ $Y2=1.93
cc_824 N_CK_c_974_n N_A_1246_89#_c_1540_n 0.00185875f $X=6.735 $Y=2.33 $X2=6.365
+ $Y2=1.93
cc_825 N_CK_c_947_n N_A_1246_89#_c_1551_n 8.95026e-19 $X=6.79 $Y=2.34 $X2=6.365
+ $Y2=1.93
cc_826 N_CK_c_974_n N_A_1246_89#_c_1551_n 0.00488871f $X=6.735 $Y=2.33 $X2=6.365
+ $Y2=1.93
cc_827 N_CK_c_946_n N_A_1246_89#_c_1558_n 2.34467e-19 $X=6.735 $Y=2.67 $X2=9.235
+ $Y2=1.93
cc_828 N_CK_c_947_n N_A_1246_89#_c_1558_n 0.0033485f $X=6.79 $Y=2.34 $X2=9.235
+ $Y2=1.93
cc_829 N_CK_c_969_n N_A_1246_89#_c_1558_n 8.38639e-19 $X=6.88 $Y=2.33 $X2=9.235
+ $Y2=1.93
cc_830 N_CK_c_974_n N_A_1246_89#_c_1558_n 0.0179446f $X=6.735 $Y=2.33 $X2=9.235
+ $Y2=1.93
cc_831 CK N_A_1246_89#_c_1558_n 0.0248956f $X=6.88 $Y=2.33 $X2=9.235 $Y2=1.93
cc_832 N_CK_c_947_n N_A_1246_89#_c_1559_n 8.66236e-19 $X=6.79 $Y=2.34 $X2=6.51
+ $Y2=1.93
cc_833 N_CK_c_974_n N_A_1246_89#_c_1559_n 0.0247156f $X=6.735 $Y=2.33 $X2=6.51
+ $Y2=1.93
cc_834 N_CK_c_946_n N_A_1084_115#_c_1707_n 0.00744372f $X=6.735 $Y=2.67
+ $X2=7.505 $Y2=2.37
cc_835 N_CK_c_947_n N_A_1084_115#_c_1707_n 0.00688829f $X=6.79 $Y=2.34 $X2=7.505
+ $Y2=2.37
cc_836 N_CK_c_946_n N_A_1084_115#_M1021_g 5.00344e-19 $X=6.735 $Y=2.67 $X2=7.685
+ $Y2=3.825
cc_837 N_CK_c_963_n N_A_1084_115#_c_1712_n 0.00688829f $X=6.762 $Y=1.575
+ $X2=7.685 $Y2=1.51
cc_838 N_CK_c_954_n N_A_1084_115#_c_1715_n 0.00554221f $X=5.405 $Y=1.425
+ $X2=5.065 $Y2=1.59
cc_839 N_CK_c_966_n N_A_1084_115#_c_1715_n 0.057541f $X=5.405 $Y=1.59 $X2=5.065
+ $Y2=1.59
cc_840 N_CK_c_968_n N_A_1084_115#_c_1715_n 0.0116326f $X=5.49 $Y=2.33 $X2=5.065
+ $Y2=1.59
cc_841 N_CK_c_971_n N_A_1084_115#_c_1715_n 0.00539276f $X=5.885 $Y=2.33
+ $X2=5.065 $Y2=1.59
cc_842 N_CK_c_972_n N_A_1084_115#_c_1715_n 0.0139004f $X=5.74 $Y=2.33 $X2=5.065
+ $Y2=1.59
cc_843 N_CK_c_975_n N_A_1084_115#_c_1715_n 6.61118e-19 $X=6.03 $Y=2.33 $X2=5.065
+ $Y2=1.59
cc_844 N_CK_c_953_n N_A_1084_115#_c_1740_n 0.00227142f $X=5.405 $Y=1.59
+ $X2=5.475 $Y2=1.17
cc_845 N_CK_c_954_n N_A_1084_115#_c_1740_n 0.0147334f $X=5.405 $Y=1.425
+ $X2=5.475 $Y2=1.17
cc_846 N_CK_c_966_n N_A_1084_115#_c_1740_n 0.0103267f $X=5.405 $Y=1.59 $X2=5.475
+ $Y2=1.17
cc_847 N_CK_c_957_n N_A_1084_115#_c_1759_n 0.00123101f $X=5.885 $Y=2.505
+ $X2=5.475 $Y2=2.925
cc_848 N_CK_c_967_n N_A_1084_115#_c_1759_n 0.00729874f $X=5.8 $Y=2.33 $X2=5.475
+ $Y2=2.925
cc_849 N_CK_c_968_n N_A_1084_115#_c_1759_n 0.00292714f $X=5.49 $Y=2.33 $X2=5.475
+ $Y2=2.925
cc_850 N_CK_c_971_n N_A_1084_115#_c_1759_n 8.86954e-19 $X=5.885 $Y=2.33
+ $X2=5.475 $Y2=2.925
cc_851 N_CK_c_947_n N_A_1084_115#_c_1719_n 2.89967e-19 $X=6.79 $Y=2.34 $X2=7.595
+ $Y2=1.59
cc_852 N_CK_c_963_n N_A_1084_115#_c_1719_n 2.26851e-19 $X=6.762 $Y=1.575
+ $X2=7.595 $Y2=1.59
cc_853 N_CK_c_947_n N_A_1084_115#_c_1721_n 0.00128484f $X=6.79 $Y=2.34 $X2=7.45
+ $Y2=1.59
cc_854 N_CK_c_953_n N_A_1084_115#_c_1721_n 0.00362401f $X=5.405 $Y=1.59 $X2=7.45
+ $Y2=1.59
cc_855 N_CK_c_963_n N_A_1084_115#_c_1721_n 0.00179204f $X=6.762 $Y=1.575
+ $X2=7.45 $Y2=1.59
cc_856 N_CK_c_966_n N_A_1084_115#_c_1721_n 0.0127028f $X=5.405 $Y=1.59 $X2=7.45
+ $Y2=1.59
cc_857 N_CK_c_967_n N_A_1084_115#_c_1721_n 0.00451177f $X=5.8 $Y=2.33 $X2=7.45
+ $Y2=1.59
cc_858 N_CK_c_971_n N_A_1084_115#_c_1721_n 6.39375e-19 $X=5.885 $Y=2.33 $X2=7.45
+ $Y2=1.59
cc_859 N_CK_c_975_n N_A_1084_115#_c_1721_n 0.0144351f $X=6.03 $Y=2.33 $X2=7.45
+ $Y2=1.59
cc_860 N_CK_c_953_n N_A_1084_115#_c_1724_n 9.79344e-19 $X=5.405 $Y=1.59 $X2=5.21
+ $Y2=1.59
cc_861 N_CK_c_966_n N_A_1084_115#_c_1724_n 0.00180575f $X=5.405 $Y=1.59 $X2=5.21
+ $Y2=1.59
cc_862 N_CK_c_972_n N_A_1084_115#_c_1724_n 0.0128239f $X=5.74 $Y=2.33 $X2=5.21
+ $Y2=1.59
cc_863 N_A_217_565#_c_1201_n N_A_704_89#_c_1347_n 0.00253253f $X=4.49 $Y=1.59
+ $X2=3.715 $Y2=1.965
cc_864 N_A_217_565#_c_1201_n N_A_704_89#_c_1348_n 0.00296105f $X=4.49 $Y=1.59
+ $X2=4.12 $Y2=2.04
cc_865 N_A_217_565#_c_1187_n N_A_704_89#_M1035_g 0.157715f $X=4.63 $Y=2.505
+ $X2=4.195 $Y2=3.825
cc_866 N_A_217_565#_c_1198_n N_A_704_89#_M1035_g 0.00493295f $X=4.725 $Y=2.505
+ $X2=4.195 $Y2=3.825
cc_867 N_A_217_565#_c_1185_n N_A_704_89#_c_1351_n 0.0342351f $X=4.63 $Y=1.59
+ $X2=5.27 $Y2=2.04
cc_868 N_A_217_565#_c_1187_n N_A_704_89#_c_1351_n 0.0307748f $X=4.63 $Y=2.505
+ $X2=5.27 $Y2=2.04
cc_869 N_A_217_565#_c_1198_n N_A_704_89#_c_1351_n 0.0113171f $X=4.725 $Y=2.505
+ $X2=5.27 $Y2=2.04
cc_870 N_A_217_565#_c_1199_n N_A_704_89#_c_1351_n 8.69982e-19 $X=4.725 $Y=1.59
+ $X2=5.27 $Y2=2.04
cc_871 N_A_217_565#_c_1201_n N_A_704_89#_c_1351_n 0.00486036f $X=4.49 $Y=1.59
+ $X2=5.27 $Y2=2.04
cc_872 N_A_217_565#_c_1252_n N_A_704_89#_c_1351_n 4.12801e-19 $X=4.635 $Y=1.59
+ $X2=5.27 $Y2=2.04
cc_873 N_A_217_565#_c_1186_n N_A_704_89#_M1031_g 0.155112f $X=4.91 $Y=2.505
+ $X2=5.345 $Y2=3.825
cc_874 N_A_217_565#_M1022_g N_A_1084_115#_c_1715_n 0.001069f $X=4.555 $Y=0.945
+ $X2=5.065 $Y2=1.59
cc_875 N_A_217_565#_M1030_g N_A_1084_115#_c_1715_n 0.0012608f $X=4.555 $Y=3.825
+ $X2=5.065 $Y2=1.59
cc_876 N_A_217_565#_c_1183_n N_A_1084_115#_c_1715_n 0.0061959f $X=4.91 $Y=1.59
+ $X2=5.065 $Y2=1.59
cc_877 N_A_217_565#_c_1186_n N_A_1084_115#_c_1715_n 0.00723389f $X=4.91 $Y=2.505
+ $X2=5.065 $Y2=1.59
cc_878 N_A_217_565#_M1028_g N_A_1084_115#_c_1715_n 0.00502021f $X=4.985 $Y=0.945
+ $X2=5.065 $Y2=1.59
cc_879 N_A_217_565#_M1032_g N_A_1084_115#_c_1715_n 0.0051844f $X=4.985 $Y=3.825
+ $X2=5.065 $Y2=1.59
cc_880 N_A_217_565#_c_1198_n N_A_1084_115#_c_1715_n 0.0700853f $X=4.725 $Y=2.505
+ $X2=5.065 $Y2=1.59
cc_881 N_A_217_565#_c_1199_n N_A_1084_115#_c_1715_n 0.0157315f $X=4.725 $Y=1.59
+ $X2=5.065 $Y2=1.59
cc_882 N_A_217_565#_c_1252_n N_A_1084_115#_c_1715_n 4.18442e-19 $X=4.635 $Y=1.59
+ $X2=5.065 $Y2=1.59
cc_883 N_A_217_565#_M1022_g N_A_1084_115#_c_1741_n 0.00136315f $X=4.555 $Y=0.945
+ $X2=5.15 $Y2=1.17
cc_884 N_A_217_565#_M1028_g N_A_1084_115#_c_1741_n 0.00979345f $X=4.985 $Y=0.945
+ $X2=5.15 $Y2=1.17
cc_885 N_A_217_565#_M1030_g N_A_1084_115#_c_1807_n 9.13132e-19 $X=4.555 $Y=3.825
+ $X2=5.15 $Y2=2.925
cc_886 N_A_217_565#_M1032_g N_A_1084_115#_c_1807_n 0.0096885f $X=4.985 $Y=3.825
+ $X2=5.15 $Y2=2.925
cc_887 N_A_217_565#_c_1183_n N_A_1084_115#_c_1724_n 0.00229064f $X=4.91 $Y=1.59
+ $X2=5.21 $Y2=1.59
cc_888 N_A_217_565#_c_1199_n N_A_1084_115#_c_1724_n 0.0012094f $X=4.725 $Y=1.59
+ $X2=5.21 $Y2=1.59
cc_889 N_A_217_565#_c_1252_n N_A_1084_115#_c_1724_n 0.0241863f $X=4.635 $Y=1.59
+ $X2=5.21 $Y2=1.59
cc_890 N_A_704_89#_c_1354_n N_A_1246_89#_M1003_g 0.0073696f $X=5.825 $Y=1.965
+ $X2=6.305 $Y2=0.945
cc_891 N_A_704_89#_c_1359_n N_A_1246_89#_M1003_g 0.0823485f $X=5.885 $Y=1.425
+ $X2=6.305 $Y2=0.945
cc_892 N_A_704_89#_c_1362_n N_A_1246_89#_M1003_g 0.0107575f $X=6.865 $Y=1.59
+ $X2=6.305 $Y2=0.945
cc_893 N_A_704_89#_c_1353_n N_A_1246_89#_c_1540_n 0.0073696f $X=5.75 $Y=2.04
+ $X2=6.365 $Y2=1.93
cc_894 N_A_704_89#_c_1362_n N_A_1246_89#_c_1540_n 0.00290516f $X=6.865 $Y=1.59
+ $X2=6.365 $Y2=1.93
cc_895 N_A_704_89#_c_1372_n N_A_1246_89#_c_1540_n 2.96928e-19 $X=7.22 $Y=1.93
+ $X2=6.365 $Y2=1.93
cc_896 N_A_704_89#_c_1354_n N_A_1246_89#_c_1551_n 0.0035305f $X=5.825 $Y=1.965
+ $X2=6.365 $Y2=1.93
cc_897 N_A_704_89#_c_1362_n N_A_1246_89#_c_1551_n 0.0219931f $X=6.865 $Y=1.59
+ $X2=6.365 $Y2=1.93
cc_898 N_A_704_89#_c_1372_n N_A_1246_89#_c_1551_n 0.00559532f $X=7.22 $Y=1.93
+ $X2=6.365 $Y2=1.93
cc_899 N_A_704_89#_c_1362_n N_A_1246_89#_c_1558_n 0.00314603f $X=6.865 $Y=1.59
+ $X2=9.235 $Y2=1.93
cc_900 N_A_704_89#_c_1369_n N_A_1246_89#_c_1558_n 6.94255e-19 $X=6.95 $Y=1.845
+ $X2=9.235 $Y2=1.93
cc_901 N_A_704_89#_c_1370_n N_A_1246_89#_c_1558_n 0.00464833f $X=7.22 $Y=2.84
+ $X2=9.235 $Y2=1.93
cc_902 N_A_704_89#_c_1372_n N_A_1246_89#_c_1558_n 0.0207528f $X=7.22 $Y=1.93
+ $X2=9.235 $Y2=1.93
cc_903 N_A_704_89#_c_1354_n N_A_1246_89#_c_1559_n 9.14174e-19 $X=5.825 $Y=1.965
+ $X2=6.51 $Y2=1.93
cc_904 N_A_704_89#_c_1362_n N_A_1246_89#_c_1559_n 0.0010261f $X=6.865 $Y=1.59
+ $X2=6.51 $Y2=1.93
cc_905 N_A_704_89#_c_1369_n N_A_1246_89#_c_1559_n 0.00122156f $X=6.95 $Y=1.845
+ $X2=6.51 $Y2=1.93
cc_906 N_A_704_89#_c_1369_n N_A_1084_115#_c_1707_n 0.00130229f $X=6.95 $Y=1.845
+ $X2=7.505 $Y2=2.37
cc_907 N_A_704_89#_c_1370_n N_A_1084_115#_c_1707_n 0.00568165f $X=7.22 $Y=2.84
+ $X2=7.505 $Y2=2.37
cc_908 N_A_704_89#_c_1372_n N_A_1084_115#_c_1707_n 0.00134862f $X=7.22 $Y=1.93
+ $X2=7.505 $Y2=2.37
cc_909 N_A_704_89#_c_1364_n N_A_1084_115#_c_1708_n 0.00595822f $X=6.95 $Y=0.865
+ $X2=7.685 $Y2=1.43
cc_910 N_A_704_89#_c_1379_n N_A_1084_115#_M1021_g 0.00666412f $X=6.95 $Y=3.205
+ $X2=7.685 $Y2=3.825
cc_911 N_A_704_89#_c_1370_n N_A_1084_115#_M1021_g 0.00331798f $X=7.22 $Y=2.84
+ $X2=7.685 $Y2=3.825
cc_912 N_A_704_89#_c_1383_n N_A_1084_115#_M1021_g 0.00560488f $X=7.22 $Y=2.925
+ $X2=7.685 $Y2=3.825
cc_913 N_A_704_89#_c_1364_n N_A_1084_115#_c_1712_n 0.00137598f $X=6.95 $Y=0.865
+ $X2=7.685 $Y2=1.51
cc_914 N_A_704_89#_c_1371_n N_A_1084_115#_c_1712_n 9.86466e-19 $X=6.95 $Y=1.59
+ $X2=7.685 $Y2=1.51
cc_915 N_A_704_89#_c_1351_n N_A_1084_115#_c_1715_n 0.0124213f $X=5.27 $Y=2.04
+ $X2=5.065 $Y2=1.59
cc_916 N_A_704_89#_M1031_g N_A_1084_115#_c_1715_n 0.0105859f $X=5.345 $Y=3.825
+ $X2=5.065 $Y2=1.59
cc_917 N_A_704_89#_c_1358_n N_A_1084_115#_c_1740_n 0.00174653f $X=5.885 $Y=1.59
+ $X2=5.475 $Y2=1.17
cc_918 N_A_704_89#_c_1359_n N_A_1084_115#_c_1740_n 0.00205316f $X=5.885 $Y=1.425
+ $X2=5.475 $Y2=1.17
cc_919 N_A_704_89#_c_1362_n N_A_1084_115#_c_1740_n 0.00436807f $X=6.865 $Y=1.59
+ $X2=5.475 $Y2=1.17
cc_920 N_A_704_89#_M1031_g N_A_1084_115#_c_1759_n 0.0157833f $X=5.345 $Y=3.825
+ $X2=5.475 $Y2=2.925
cc_921 N_A_704_89#_c_1369_n N_A_1084_115#_c_1719_n 0.00520507f $X=6.95 $Y=1.845
+ $X2=7.595 $Y2=1.59
cc_922 N_A_704_89#_c_1370_n N_A_1084_115#_c_1719_n 0.039533f $X=7.22 $Y=2.84
+ $X2=7.595 $Y2=1.59
cc_923 N_A_704_89#_c_1371_n N_A_1084_115#_c_1719_n 0.00358095f $X=6.95 $Y=1.59
+ $X2=7.595 $Y2=1.59
cc_924 N_A_704_89#_c_1372_n N_A_1084_115#_c_1719_n 0.00955403f $X=7.22 $Y=1.93
+ $X2=7.595 $Y2=1.59
cc_925 N_A_704_89#_c_1351_n N_A_1084_115#_c_1721_n 0.00156696f $X=5.27 $Y=2.04
+ $X2=7.45 $Y2=1.59
cc_926 N_A_704_89#_c_1353_n N_A_1084_115#_c_1721_n 0.00244106f $X=5.75 $Y=2.04
+ $X2=7.45 $Y2=1.59
cc_927 N_A_704_89#_c_1357_n N_A_1084_115#_c_1721_n 5.19983e-19 $X=5.345 $Y=2.04
+ $X2=7.45 $Y2=1.59
cc_928 N_A_704_89#_c_1358_n N_A_1084_115#_c_1721_n 0.00455939f $X=5.885 $Y=1.59
+ $X2=7.45 $Y2=1.59
cc_929 N_A_704_89#_c_1362_n N_A_1084_115#_c_1721_n 0.0492477f $X=6.865 $Y=1.59
+ $X2=7.45 $Y2=1.59
cc_930 N_A_704_89#_c_1371_n N_A_1084_115#_c_1721_n 0.0117855f $X=6.95 $Y=1.59
+ $X2=7.45 $Y2=1.59
cc_931 N_A_704_89#_c_1372_n N_A_1084_115#_c_1721_n 0.00219678f $X=7.22 $Y=1.93
+ $X2=7.45 $Y2=1.59
cc_932 N_A_704_89#_c_1351_n N_A_1084_115#_c_1724_n 0.00120486f $X=5.27 $Y=2.04
+ $X2=5.21 $Y2=1.59
cc_933 N_A_704_89#_c_1364_n N_A_1084_115#_c_1725_n 0.0010241f $X=6.95 $Y=0.865
+ $X2=7.595 $Y2=1.59
cc_934 N_A_704_89#_c_1369_n N_A_1084_115#_c_1725_n 6.33705e-19 $X=6.95 $Y=1.845
+ $X2=7.595 $Y2=1.59
cc_935 N_A_704_89#_c_1379_n N_A_1469_565#_c_1970_n 0.0585029f $X=6.95 $Y=3.205
+ $X2=7.47 $Y2=3.545
cc_936 N_A_704_89#_c_1379_n N_A_1469_565#_c_1982_n 0.00811594f $X=6.95 $Y=3.205
+ $X2=7.555 $Y2=3.37
cc_937 N_A_1246_89#_c_1558_n N_A_1084_115#_c_1707_n 0.00586968f $X=9.235 $Y=1.93
+ $X2=7.505 $Y2=2.37
cc_938 N_A_1246_89#_c_1558_n N_A_1084_115#_c_1712_n 6.8924e-19 $X=9.235 $Y=1.93
+ $X2=7.685 $Y2=1.51
cc_939 N_A_1246_89#_c_1558_n N_A_1084_115#_c_1714_n 0.00207076f $X=9.235 $Y=1.93
+ $X2=7.685 $Y2=2.505
cc_940 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1719_n 0.0010677f $X=8.26 $Y=0.865
+ $X2=7.595 $Y2=1.59
cc_941 N_A_1246_89#_c_1556_n N_A_1084_115#_c_1719_n 0.00422342f $X=8.845 $Y=1.93
+ $X2=7.595 $Y2=1.59
cc_942 N_A_1246_89#_c_1558_n N_A_1084_115#_c_1719_n 0.0169834f $X=9.235 $Y=1.93
+ $X2=7.595 $Y2=1.59
cc_943 N_A_1246_89#_M1003_g N_A_1084_115#_c_1721_n 0.00231271f $X=6.305 $Y=0.945
+ $X2=7.45 $Y2=1.59
cc_944 N_A_1246_89#_c_1540_n N_A_1084_115#_c_1721_n 0.00187603f $X=6.365 $Y=1.93
+ $X2=7.45 $Y2=1.59
cc_945 N_A_1246_89#_c_1551_n N_A_1084_115#_c_1721_n 0.00166223f $X=6.365 $Y=1.93
+ $X2=7.45 $Y2=1.59
cc_946 N_A_1246_89#_c_1558_n N_A_1084_115#_c_1721_n 0.0841111f $X=9.235 $Y=1.93
+ $X2=7.45 $Y2=1.59
cc_947 N_A_1246_89#_c_1559_n N_A_1084_115#_c_1721_n 0.0289631f $X=6.51 $Y=1.93
+ $X2=7.45 $Y2=1.59
cc_948 N_A_1246_89#_c_1552_n N_A_1084_115#_c_1725_n 0.00247064f $X=8.26 $Y=0.865
+ $X2=7.595 $Y2=1.59
cc_949 N_A_1246_89#_c_1556_n N_A_1084_115#_c_1725_n 0.00385422f $X=8.845 $Y=1.93
+ $X2=7.595 $Y2=1.59
cc_950 N_A_1246_89#_c_1558_n N_A_1084_115#_c_1725_n 0.027605f $X=9.235 $Y=1.93
+ $X2=7.595 $Y2=1.59
cc_951 N_A_1246_89#_c_1542_n N_QN_M1006_g 0.0153129f $X=9.382 $Y=1.765 $X2=9.925
+ $Y2=0.945
cc_952 N_A_1246_89#_c_1543_n N_QN_M1006_g 0.0276883f $X=9.47 $Y=1.39 $X2=9.925
+ $Y2=0.945
cc_953 N_A_1246_89#_c_1557_n N_QN_M1006_g 4.79563e-19 $X=9.38 $Y=1.93 $X2=9.925
+ $Y2=0.945
cc_954 N_A_1246_89#_c_1549_n N_QN_M1019_g 0.0102953f $X=9.47 $Y=2.595 $X2=9.925
+ $Y2=3.825
cc_955 N_A_1246_89#_c_1550_n N_QN_M1019_g 0.0240292f $X=9.47 $Y=2.745 $X2=9.925
+ $Y2=3.825
cc_956 N_A_1246_89#_c_1541_n N_QN_c_1868_n 0.021196f $X=9.38 $Y=1.93 $X2=9.865
+ $Y2=2.135
cc_957 N_A_1246_89#_c_1557_n N_QN_c_1868_n 3.0115e-19 $X=9.38 $Y=1.93 $X2=9.865
+ $Y2=2.135
cc_958 N_A_1246_89#_c_1560_n N_QN_c_1868_n 4.60229e-19 $X=9.38 $Y=1.93 $X2=9.865
+ $Y2=2.135
cc_959 N_A_1246_89#_c_1543_n N_QN_c_1869_n 0.00715777f $X=9.47 $Y=1.39 $X2=9.28
+ $Y2=0.865
cc_960 N_A_1246_89#_c_1548_n N_QN_c_1869_n 0.00310506f $X=9.47 $Y=1.54 $X2=9.28
+ $Y2=0.865
cc_961 N_A_1246_89#_c_1549_n N_QN_c_1873_n 0.00521938f $X=9.47 $Y=2.595 $X2=9.28
+ $Y2=2.7
cc_962 N_A_1246_89#_c_1550_n N_QN_c_1873_n 0.00746388f $X=9.47 $Y=2.745 $X2=9.28
+ $Y2=2.7
cc_963 N_A_1246_89#_c_1555_n N_QN_c_1873_n 0.0926802f $X=8.76 $Y=3.545 $X2=9.28
+ $Y2=2.7
cc_964 N_A_1246_89#_c_1542_n N_QN_c_1874_n 0.00722072f $X=9.382 $Y=1.765
+ $X2=9.78 $Y2=1.59
cc_965 N_A_1246_89#_c_1548_n N_QN_c_1874_n 0.0107741f $X=9.47 $Y=1.54 $X2=9.78
+ $Y2=1.59
cc_966 N_A_1246_89#_c_1557_n N_QN_c_1874_n 0.0110498f $X=9.38 $Y=1.93 $X2=9.78
+ $Y2=1.59
cc_967 N_A_1246_89#_c_1560_n N_QN_c_1874_n 0.00387586f $X=9.38 $Y=1.93 $X2=9.78
+ $Y2=1.59
cc_968 N_A_1246_89#_c_1541_n N_QN_c_1876_n 0.00308111f $X=9.38 $Y=1.93 $X2=9.365
+ $Y2=1.59
cc_969 N_A_1246_89#_c_1556_n N_QN_c_1876_n 0.00372477f $X=8.845 $Y=1.93
+ $X2=9.365 $Y2=1.59
cc_970 N_A_1246_89#_c_1557_n N_QN_c_1876_n 0.0120703f $X=9.38 $Y=1.93 $X2=9.365
+ $Y2=1.59
cc_971 N_A_1246_89#_c_1558_n N_QN_c_1876_n 0.0010572f $X=9.235 $Y=1.93 $X2=9.365
+ $Y2=1.59
cc_972 N_A_1246_89#_c_1560_n N_QN_c_1876_n 0.00336135f $X=9.38 $Y=1.93 $X2=9.365
+ $Y2=1.59
cc_973 N_A_1246_89#_c_1549_n N_QN_c_1877_n 0.0152835f $X=9.47 $Y=2.595 $X2=9.78
+ $Y2=2.505
cc_974 N_A_1246_89#_c_1550_n N_QN_c_1877_n 0.00248624f $X=9.47 $Y=2.745 $X2=9.78
+ $Y2=2.505
cc_975 N_A_1246_89#_c_1557_n N_QN_c_1877_n 0.00426371f $X=9.38 $Y=1.93 $X2=9.78
+ $Y2=2.505
cc_976 N_A_1246_89#_c_1560_n N_QN_c_1877_n 0.00253233f $X=9.38 $Y=1.93 $X2=9.78
+ $Y2=2.505
cc_977 N_A_1246_89#_c_1541_n N_QN_c_1878_n 0.00265611f $X=9.38 $Y=1.93 $X2=9.365
+ $Y2=2.505
cc_978 N_A_1246_89#_c_1555_n N_QN_c_1878_n 0.00826781f $X=8.76 $Y=3.545
+ $X2=9.365 $Y2=2.505
cc_979 N_A_1246_89#_c_1557_n N_QN_c_1878_n 0.00471962f $X=9.38 $Y=1.93 $X2=9.365
+ $Y2=2.505
cc_980 N_A_1246_89#_c_1558_n N_QN_c_1878_n 9.40773e-19 $X=9.235 $Y=1.93
+ $X2=9.365 $Y2=2.505
cc_981 N_A_1246_89#_c_1560_n N_QN_c_1878_n 0.00140341f $X=9.38 $Y=1.93 $X2=9.365
+ $Y2=2.505
cc_982 N_A_1246_89#_c_1541_n N_QN_c_1879_n 0.00216137f $X=9.38 $Y=1.93 $X2=9.865
+ $Y2=2.135
cc_983 N_A_1246_89#_c_1542_n N_QN_c_1879_n 0.00323473f $X=9.382 $Y=1.765
+ $X2=9.865 $Y2=2.135
cc_984 N_A_1246_89#_c_1549_n N_QN_c_1879_n 0.00226435f $X=9.47 $Y=2.595
+ $X2=9.865 $Y2=2.135
cc_985 N_A_1246_89#_c_1557_n N_QN_c_1879_n 0.00987106f $X=9.38 $Y=1.93 $X2=9.865
+ $Y2=2.135
cc_986 N_A_1246_89#_c_1560_n N_QN_c_1879_n 0.00377439f $X=9.38 $Y=1.93 $X2=9.865
+ $Y2=2.135
cc_987 N_A_1246_89#_c_1550_n QN 0.00718989f $X=9.47 $Y=2.745 $X2=9.285 $Y2=2.7
cc_988 N_A_1246_89#_c_1555_n QN 0.00721908f $X=8.76 $Y=3.545 $X2=9.285 $Y2=2.7
cc_989 N_A_1246_89#_c_1557_n QN 0.00359685f $X=9.38 $Y=1.93 $X2=9.285 $Y2=2.7
cc_990 N_A_1246_89#_c_1560_n QN 0.00842298f $X=9.38 $Y=1.93 $X2=9.285 $Y2=2.7
cc_991 N_A_1084_115#_c_1759_n A_1012_565# 0.00310684f $X=5.475 $Y=2.925 $X2=5.06
+ $Y2=2.825
cc_992 N_A_1084_115#_c_1807_n A_1012_565# 0.00144354f $X=5.15 $Y=2.925 $X2=5.06
+ $Y2=2.825
cc_993 N_A_1084_115#_M1021_g N_A_1469_565#_c_1973_n 0.0157576f $X=7.685 $Y=3.825
+ $X2=8.245 $Y2=3.37
cc_994 N_A_1084_115#_c_1719_n N_A_1469_565#_c_1973_n 0.00125278f $X=7.595
+ $Y=1.59 $X2=8.245 $Y2=3.37
cc_995 N_A_1084_115#_c_1714_n N_A_1469_565#_c_1982_n 0.0020255f $X=7.685
+ $Y=2.505 $X2=7.555 $Y2=3.37
cc_996 N_A_1084_115#_c_1719_n N_A_1469_565#_c_1982_n 7.57421e-19 $X=7.595
+ $Y=1.59 $X2=7.555 $Y2=3.37
cc_997 N_A_1084_115#_c_1715_n A_1012_115# 9.4749e-19 $X=5.065 $Y=1.59 $X2=5.06
+ $Y2=0.575
cc_998 N_A_1084_115#_c_1740_n A_1012_115# 0.00337089f $X=5.475 $Y=1.17 $X2=5.06
+ $Y2=0.575
cc_999 N_A_1084_115#_c_1741_n A_1012_115# 0.00148865f $X=5.15 $Y=1.17 $X2=5.06
+ $Y2=0.575
cc_1000 N_QN_M1019_g N_Q_c_1993_n 0.00331568f $X=9.925 $Y=3.825 $X2=10.14
+ $Y2=3.07
cc_1001 N_QN_M1006_g N_Q_c_1991_n 0.0330655f $X=9.925 $Y=0.945 $X2=10.255
+ $Y2=2.745
cc_1002 N_QN_c_1874_n N_Q_c_1991_n 0.0111776f $X=9.78 $Y=1.59 $X2=10.255
+ $Y2=2.745
cc_1003 N_QN_c_1877_n N_Q_c_1991_n 0.0111776f $X=9.78 $Y=2.505 $X2=10.255
+ $Y2=2.745
cc_1004 N_QN_c_1879_n N_Q_c_1991_n 0.0438362f $X=9.865 $Y=2.135 $X2=10.255
+ $Y2=2.745
cc_1005 N_QN_M1006_g N_Q_c_1992_n 0.00373219f $X=9.925 $Y=0.945 $X2=10.255
+ $Y2=1.255
cc_1006 N_QN_M1019_g N_Q_c_1997_n 0.00495318f $X=9.925 $Y=3.825 $X2=10.255
+ $Y2=2.83
cc_1007 N_QN_M1019_g Q 0.0105324f $X=9.925 $Y=3.825 $X2=10.14 $Y2=3.07
cc_1008 N_QN_c_1877_n Q 0.00228117f $X=9.78 $Y=2.505 $X2=10.14 $Y2=3.07
