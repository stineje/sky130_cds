* File: sky130_osu_sc_15T_ls__oai21_l.spice
* Created: Fri Nov 12 14:58:55 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__oai21_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__oai21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_A0_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_115#_M1000_d N_A1_M1000_g N_GND_M1003_d N_GND_M1003_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_115#_M1000_d N_GND_M1003_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_110_565# N_A0_M1001_g N_Y_M1001_s N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.9 A=0.3 P=4.3 MULT=1
MM1005 N_VDD_M1005_d N_A1_M1005_g A_110_565# N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.383129 AS=0.21 PD=2.87117 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333
+ SA=75000.5 SB=75000.5 A=0.3 P=4.3 MULT=1
MM1004 N_Y_M1004_d N_B0_M1004_g N_VDD_M1005_d N_VDD_M1001_b PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.241371 PD=3.05 PS=1.80883 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75001 SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1001_b NWDIODE A=5.64925 P=9.73
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__oai21_l.pxi.spice"
*
.ends
*
*
