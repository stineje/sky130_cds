* File: sky130_osu_sc_18T_ls__and2_6.pex.spice
* Created: Fri Nov 12 13:39:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__AND2_6%GND 1 2 3 4 47 49 57 59 66 68 75 77 85
+ 95 97
r105 95 97 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.06 $Y2=0.152
r106 83 85 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.825
r107 78 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r108 77 83 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=3.615 $Y=0.152
+ $X2=3.7 $Y2=0.305
r109 73 91 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r110 73 75 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.825
r111 69 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r112 68 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r113 64 90 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r114 64 66 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r115 59 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r116 55 57 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r117 47 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=0.19
+ $X2=3.06 $Y2=0.19
r118 47 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r119 47 55 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r120 47 49 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r121 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r122 47 77 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r123 47 78 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r124 47 68 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r125 47 69 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r126 47 59 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r127 47 60 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r128 47 49 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r129 4 85 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.825
r130 3 75 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r131 2 66 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r132 1 57 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_6%VDD 1 2 3 4 5 41 45 49 55 59 65 69 75 79
+ 86 97 101
r70 97 101 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.06 $Y2=6.507
r71 91 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r72 86 89 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.7 $Y=3.455
+ $X2=3.7 $Y2=5.835
r73 84 89 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.7 $Y=6.355 $X2=3.7
+ $Y2=5.835
r74 82 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=6.47
+ $X2=3.06 $Y2=6.47
r75 80 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=6.507
+ $X2=2.84 $Y2=6.507
r76 80 82 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=6.507
+ $X2=3.06 $Y2=6.507
r77 79 84 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=3.615 $Y=6.507
+ $X2=3.7 $Y2=6.355
r78 79 82 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=6.507
+ $X2=3.06 $Y2=6.507
r79 75 78 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r80 73 95 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.84 $Y2=6.507
r81 73 78 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.84 $Y2=5.835
r82 70 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=1.98 $Y2=6.507
r83 70 72 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=2.38 $Y2=6.507
r84 69 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.84 $Y2=6.507
r85 69 72 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.38 $Y2=6.507
r86 65 68 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r87 63 94 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=6.507
r88 63 68 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r89 60 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r90 60 62 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r91 59 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.98 $Y2=6.507
r92 59 62 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r93 55 58 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r94 53 93 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r95 53 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r96 50 91 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r97 50 52 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r98 49 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r99 49 52 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r100 45 48 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r101 43 91 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r102 43 48 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r103 41 82 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r104 41 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r105 41 62 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r106 41 52 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r107 41 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r108 5 89 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=5.835
r109 5 86 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=3.455
r110 4 78 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r111 4 75 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r112 3 68 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r113 3 65 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r114 2 58 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r115 2 55 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r116 1 48 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r117 1 45 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_6%A 3 7 12 15 23
r29 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=3.33
+ $X2=0.235 $Y2=3.33
r31 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.235 $Y=2.765
+ $X2=0.235 $Y2=3.33
r32 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.235
+ $Y=2.765 $X2=0.235 $Y2=2.765
r33 10 12 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.235 $Y=2.765
+ $X2=0.475 $Y2=2.765
r34 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=2.765
r35 5 7 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=4.585
r36 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=2.765
r37 1 3 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_6%B 3 7 10 13 21
c38 7 0 1.42883e-19 $X=0.905 $Y=4.585
r39 19 21 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.915 $Y=2.96
+ $X2=0.92 $Y2=2.96
r40 16 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.915 $Y=2.96
+ $X2=0.915 $Y2=2.96
r41 13 16 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.915 $Y=2.425
+ $X2=0.915 $Y2=2.96
r42 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=2.425 $X2=0.915 $Y2=2.425
r43 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.425
+ $X2=0.905 $Y2=2.26
r44 5 10 49.0931 $w=2.9e-07 $l=1.7e-07 $layer=POLY_cond $X=0.905 $Y=2.595
+ $X2=0.905 $Y2=2.425
r45 5 7 1020.4 $w=1.5e-07 $l=1.99e-06 $layer=POLY_cond $X=0.905 $Y=2.595
+ $X2=0.905 $Y2=4.585
r46 3 11 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_6%A_27_115# 1 3 11 14 15 17 18 20 24 26 28
+ 29 31 35 37 39 40 42 46 48 50 51 53 57 60 61 63 64 66 70 72 74 75 80 81 82 83
+ 84 85 86 87 88 91 94 97 101 103 110
c188 57 0 1.33323e-19 $X=3.055 $Y=1.075
c189 46 0 1.33323e-19 $X=2.625 $Y=1.075
c190 35 0 1.33323e-19 $X=2.195 $Y=1.075
c191 24 0 1.33323e-19 $X=1.765 $Y=1.075
r192 108 110 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.575 $Y=3.63
+ $X2=0.69 $Y2=3.63
r193 105 107 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=1.935
+ $X2=0.575 $Y2=1.935
r194 101 107 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=1.935
+ $X2=0.575 $Y2=1.935
r195 101 103 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.66 $Y=1.935
+ $X2=1.395 $Y2=1.935
r196 97 99 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.69 $Y=3.795
+ $X2=0.69 $Y2=5.835
r197 95 110 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.715
+ $X2=0.69 $Y2=3.63
r198 95 97 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.715
+ $X2=0.69 $Y2=3.795
r199 94 108 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.575 $Y=3.545
+ $X2=0.575 $Y2=3.63
r200 93 107 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.575 $Y=2.02
+ $X2=0.575 $Y2=1.935
r201 93 94 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.575 $Y=2.02
+ $X2=0.575 $Y2=3.545
r202 89 105 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=1.935
r203 89 91 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r204 78 103 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.935 $X2=1.395 $Y2=1.935
r205 78 79 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.935
+ $X2=1.395 $Y2=2.1
r206 75 78 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.395 $Y=1.845
+ $X2=1.395 $Y2=1.935
r207 75 76 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=1.845
+ $X2=1.395 $Y2=1.77
r208 72 74 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=3.485 $Y=2.96
+ $X2=3.485 $Y2=4.585
r209 68 70 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.075
r210 67 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.885
+ $X2=3.055 $Y2=2.885
r211 66 72 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=2.885
+ $X2=3.485 $Y2=2.96
r212 66 67 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.885
+ $X2=3.13 $Y2=2.885
r213 65 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.845
+ $X2=3.055 $Y2=1.845
r214 64 68 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.485 $Y2=1.77
r215 64 65 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.13 $Y2=1.845
r216 61 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.96
+ $X2=3.055 $Y2=2.885
r217 61 63 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=3.055 $Y=2.96
+ $X2=3.055 $Y2=4.585
r218 60 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.81
+ $X2=3.055 $Y2=2.885
r219 59 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.92
+ $X2=3.055 $Y2=1.845
r220 59 60 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.055 $Y=1.92
+ $X2=3.055 $Y2=2.81
r221 55 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.845
r222 55 57 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.075
r223 54 86 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.885
+ $X2=2.625 $Y2=2.885
r224 53 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.885
+ $X2=3.055 $Y2=2.885
r225 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.885
+ $X2=2.7 $Y2=2.885
r226 52 85 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.845
+ $X2=2.625 $Y2=1.845
r227 51 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=3.055 $Y2=1.845
r228 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=2.7 $Y2=1.845
r229 48 86 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.96
+ $X2=2.625 $Y2=2.885
r230 48 50 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.625 $Y=2.96
+ $X2=2.625 $Y2=4.585
r231 44 85 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.845
r232 44 46 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.075
r233 43 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.885
+ $X2=2.195 $Y2=2.885
r234 42 86 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.625 $Y2=2.885
r235 42 43 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.27 $Y2=2.885
r236 41 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.195 $Y2=1.845
r237 40 85 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.625 $Y2=1.845
r238 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.27 $Y2=1.845
r239 37 84 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=2.885
r240 37 39 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=4.585
r241 33 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.845
r242 33 35 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r243 32 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.885
+ $X2=1.765 $Y2=2.885
r244 31 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=2.195 $Y2=2.885
r245 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=1.84 $Y2=2.885
r246 30 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.765 $Y2=1.845
r247 29 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.845
r248 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r249 26 82 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=2.885
r250 26 28 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r251 22 81 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.845
r252 22 24 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r253 21 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.53 $Y=1.845
+ $X2=1.395 $Y2=1.845
r254 20 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.765 $Y2=1.845
r255 20 21 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.53 $Y2=1.845
r256 19 80 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.885
+ $X2=1.335 $Y2=2.885
r257 18 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.885
r258 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.41 $Y2=2.885
r259 15 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=2.885
r260 15 17 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r261 14 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.81
+ $X2=1.335 $Y2=2.885
r262 14 79 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.335 $Y=2.81
+ $X2=1.335 $Y2=2.1
r263 11 76 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=1.77
r264 3 99 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r265 3 97 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.795
r266 1 91 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_6%Y 1 2 3 7 8 9 26 32 40 46 54 60 67 68 70
+ 72 74 77 78 79 80 81 82 83
c124 82 0 1.33323e-19 $X=3.27 $Y=1.595
c125 79 0 2.66647e-19 $X=2.555 $Y=1.48
c126 67 0 1.33323e-19 $X=1.55 $Y=1.595
c127 32 0 1.42883e-19 $X=1.55 $Y=2.59
r128 83 95 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.475
+ $X2=3.27 $Y2=2.59
r129 82 93 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.595
+ $X2=3.27 $Y2=1.48
r130 82 83 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=3.27 $Y=1.595
+ $X2=3.27 $Y2=2.475
r131 81 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.59
+ $X2=2.41 $Y2=2.59
r132 80 95 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.59
+ $X2=3.27 $Y2=2.59
r133 80 81 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.59
+ $X2=2.555 $Y2=2.59
r134 79 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.48
+ $X2=2.41 $Y2=1.48
r135 78 93 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.48
+ $X2=3.27 $Y2=1.48
r136 78 79 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.48
+ $X2=2.555 $Y2=1.48
r137 77 91 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.475
+ $X2=2.41 $Y2=2.59
r138 76 89 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=1.48
r139 76 77 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=2.475
r140 75 87 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.59
+ $X2=1.55 $Y2=2.59
r141 74 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.59
+ $X2=2.41 $Y2=2.59
r142 74 75 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.59
+ $X2=1.695 $Y2=2.59
r143 73 85 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.48
+ $X2=1.55 $Y2=1.48
r144 72 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=2.41 $Y2=1.48
r145 72 73 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=1.695 $Y2=1.48
r146 68 87 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r147 68 70 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r148 67 85 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r149 67 70 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r150 63 65 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.27 $Y=3.455
+ $X2=3.27 $Y2=5.835
r151 60 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.59
+ $X2=3.27 $Y2=2.59
r152 60 63 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.27 $Y=2.59
+ $X2=3.27 $Y2=3.455
r153 57 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.48
+ $X2=3.27 $Y2=1.48
r154 54 57 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.27 $Y=0.825
+ $X2=3.27 $Y2=1.48
r155 49 51 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r156 46 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.59
+ $X2=2.41 $Y2=2.59
r157 46 49 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.41 $Y=2.59
+ $X2=2.41 $Y2=3.455
r158 43 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.48
+ $X2=2.41 $Y2=1.48
r159 40 43 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.41 $Y=0.825
+ $X2=2.41 $Y2=1.48
r160 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r161 32 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r162 32 35 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r163 29 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r164 26 29 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r165 9 65 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=5.835
r166 9 63 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=3.455
r167 8 51 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r168 8 49 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r169 7 37 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r170 7 35 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r171 3 54 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.825
r172 2 40 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r173 1 26 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

