* File: sky130_osu_sc_12T_hs__and2_1.pxi.spice
* Created: Fri Nov 12 15:06:44 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__AND2_1%GND N_GND_M1002_d N_GND_M1003_b N_GND_c_2_p
+ N_GND_c_8_p GND N_GND_c_3_p PM_SKY130_OSU_SC_12T_HS__AND2_1%GND
x_PM_SKY130_OSU_SC_12T_HS__AND2_1%VDD N_VDD_M1000_s N_VDD_M1004_d N_VDD_M1000_b
+ N_VDD_c_38_p N_VDD_c_39_p N_VDD_c_50_p N_VDD_c_57_p VDD N_VDD_c_40_p
+ PM_SKY130_OSU_SC_12T_HS__AND2_1%VDD
x_PM_SKY130_OSU_SC_12T_HS__AND2_1%A N_A_M1003_g N_A_M1000_g N_A_c_69_n
+ N_A_c_70_n A PM_SKY130_OSU_SC_12T_HS__AND2_1%A
x_PM_SKY130_OSU_SC_12T_HS__AND2_1%B N_B_M1002_g N_B_M1004_g N_B_c_103_n
+ N_B_c_104_n B PM_SKY130_OSU_SC_12T_HS__AND2_1%B
x_PM_SKY130_OSU_SC_12T_HS__AND2_1%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1000_d N_A_27_115#_M1001_g N_A_27_115#_M1005_g
+ N_A_27_115#_c_142_n N_A_27_115#_c_143_n N_A_27_115#_c_144_n
+ N_A_27_115#_c_145_n N_A_27_115#_c_148_n N_A_27_115#_c_149_n
+ N_A_27_115#_c_158_n N_A_27_115#_c_150_n N_A_27_115#_c_152_n
+ N_A_27_115#_c_153_n N_A_27_115#_c_174_n
+ PM_SKY130_OSU_SC_12T_HS__AND2_1%A_27_115#
x_PM_SKY130_OSU_SC_12T_HS__AND2_1%Y N_Y_M1001_d N_Y_M1005_d N_Y_c_208_n
+ N_Y_c_211_n Y N_Y_c_213_n N_Y_c_215_n PM_SKY130_OSU_SC_12T_HS__AND2_1%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.079001f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_A_M1003_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_A_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.85
cc_4 N_GND_M1003_b N_A_c_69_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.285
cc_5 N_GND_M1003_b N_A_c_70_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.285
cc_6 N_GND_M1003_b N_B_M1002_g 0.0444472f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.85
cc_7 N_GND_c_2_p N_B_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.85
cc_8 N_GND_c_8_p N_B_M1002_g 0.00319969f $X=1.05 $Y=0.755 $X2=0.835 $Y2=0.85
cc_9 N_GND_c_3_p N_B_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.85
cc_10 N_GND_M1003_b N_B_M1004_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_11 N_GND_M1003_b N_B_c_103_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.945
cc_12 N_GND_M1003_b N_B_c_104_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.945
cc_13 N_GND_M1003_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.48
cc_14 N_GND_M1003_b N_A_27_115#_M1001_g 0.0324724f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.85
cc_15 N_GND_c_8_p N_A_27_115#_M1001_g 0.00610843f $X=1.05 $Y=0.755 $X2=1.335
+ $Y2=0.85
cc_16 N_GND_c_3_p N_A_27_115#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=0.85
cc_17 N_GND_M1003_b N_A_27_115#_c_142_n 0.0373102f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=1.62
cc_18 N_GND_M1003_b N_A_27_115#_c_143_n 0.0470206f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.33
cc_19 N_GND_M1003_b N_A_27_115#_c_144_n 0.0076653f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.48
cc_20 N_GND_M1003_b N_A_27_115#_c_145_n 0.0128494f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_21 N_GND_c_2_p N_A_27_115#_c_145_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_22 N_GND_c_3_p N_A_27_115#_c_145_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_23 N_GND_M1003_b N_A_27_115#_c_148_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.455
cc_24 N_GND_M1003_b N_A_27_115#_c_149_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.455
cc_25 N_GND_M1003_b N_A_27_115#_c_150_n 0.0240789f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_26 N_GND_c_8_p N_A_27_115#_c_150_n 0.00704977f $X=1.05 $Y=0.755 $X2=1.43
+ $Y2=1.455
cc_27 N_GND_M1003_b N_A_27_115#_c_152_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.455
cc_28 N_GND_M1003_b N_A_27_115#_c_153_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.065
cc_29 N_GND_M1003_b N_Y_c_208_n 0.00897448f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_30 N_GND_c_8_p N_Y_c_208_n 0.00806382f $X=1.05 $Y=0.755 $X2=1.55 $Y2=0.755
cc_31 N_GND_c_3_p N_Y_c_208_n 0.00471849f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.755
cc_32 N_GND_M1003_b N_Y_c_211_n 0.0163869f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_33 N_GND_M1003_b Y 0.0396622f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.74
cc_34 N_GND_M1003_b N_Y_c_213_n 0.0122717f $X=-0.045 $Y=0 $X2=1.55 $Y2=1
cc_35 N_GND_c_8_p N_Y_c_213_n 0.00119317f $X=1.05 $Y=0.755 $X2=1.55 $Y2=1
cc_36 N_GND_M1003_b N_Y_c_215_n 0.0141689f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_37 N_VDD_M1000_b N_A_M1000_g 0.0189471f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_38 N_VDD_c_38_p N_A_M1000_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=3.235
cc_39 N_VDD_c_39_p N_A_M1000_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.235
cc_40 N_VDD_c_40_p N_A_M1000_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.235
cc_41 N_VDD_M1000_b N_A_c_69_n 0.0111025f $X=-0.045 $Y=2.425 $X2=0.475 $Y2=2.285
cc_42 N_VDD_M1000_s N_A_c_70_n 0.0127298f $X=0.135 $Y=2.605 $X2=0.27 $Y2=2.285
cc_43 N_VDD_M1000_b N_A_c_70_n 0.00612103f $X=-0.045 $Y=2.425 $X2=0.27 $Y2=2.285
cc_44 N_VDD_c_38_p N_A_c_70_n 0.00370742f $X=0.26 $Y=3.635 $X2=0.27 $Y2=2.285
cc_45 N_VDD_M1000_s A 0.00742066f $X=0.135 $Y=2.605 $X2=0.275 $Y2=2.85
cc_46 N_VDD_M1000_b A 0.00970321f $X=-0.045 $Y=2.425 $X2=0.275 $Y2=2.85
cc_47 N_VDD_c_38_p A 0.00434783f $X=0.26 $Y=3.635 $X2=0.275 $Y2=2.85
cc_48 N_VDD_M1000_b N_B_M1004_g 0.0187476f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_49 N_VDD_c_39_p N_B_M1004_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.235
cc_50 N_VDD_c_50_p N_B_M1004_g 0.00337744f $X=1.12 $Y=3.295 $X2=0.905 $Y2=3.235
cc_51 N_VDD_c_40_p N_B_M1004_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.905 $Y2=3.235
cc_52 N_VDD_M1000_b N_B_c_104_n 0.00170274f $X=-0.045 $Y=2.425 $X2=0.95
+ $Y2=1.945
cc_53 N_VDD_M1000_b B 0.00856863f $X=-0.045 $Y=2.425 $X2=0.955 $Y2=2.48
cc_54 N_VDD_c_50_p B 0.00240671f $X=1.12 $Y=3.295 $X2=0.955 $Y2=2.48
cc_55 N_VDD_M1000_b N_A_27_115#_c_144_n 0.0267233f $X=-0.045 $Y=2.425 $X2=1.352
+ $Y2=2.48
cc_56 N_VDD_c_50_p N_A_27_115#_c_144_n 0.00337744f $X=1.12 $Y=3.295 $X2=1.352
+ $Y2=2.48
cc_57 N_VDD_c_57_p N_A_27_115#_c_144_n 0.00606474f $X=1.12 $Y=4.287 $X2=1.352
+ $Y2=2.48
cc_58 N_VDD_c_40_p N_A_27_115#_c_144_n 0.00468827f $X=1.02 $Y=4.25 $X2=1.352
+ $Y2=2.48
cc_59 N_VDD_M1000_b N_A_27_115#_c_158_n 0.00155118f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=3.295
cc_60 N_VDD_c_39_p N_A_27_115#_c_158_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69
+ $Y2=3.295
cc_61 N_VDD_c_40_p N_A_27_115#_c_158_n 0.00475776f $X=1.02 $Y=4.25 $X2=0.69
+ $Y2=3.295
cc_62 N_VDD_M1000_b N_A_27_115#_c_153_n 8.22047e-19 $X=-0.045 $Y=2.425 $X2=0.65
+ $Y2=3.065
cc_63 N_VDD_M1000_b N_Y_c_211_n 0.0100094f $X=-0.045 $Y=2.425 $X2=1.55 $Y2=2.11
cc_64 N_VDD_c_57_p N_Y_c_211_n 0.00757793f $X=1.12 $Y=4.287 $X2=1.55 $Y2=2.11
cc_65 N_VDD_c_40_p N_Y_c_211_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.55 $Y2=2.11
cc_66 N_A_M1003_g N_B_M1002_g 0.101204f $X=0.475 $Y=0.85 $X2=0.835 $Y2=0.85
cc_67 N_A_M1003_g N_B_M1004_g 0.048305f $X=0.475 $Y=0.85 $X2=0.905 $Y2=3.235
cc_68 N_A_M1003_g N_B_c_104_n 7.8234e-19 $X=0.475 $Y=0.85 $X2=0.95 $Y2=1.945
cc_69 N_A_M1003_g N_A_27_115#_c_145_n 0.0128217f $X=0.475 $Y=0.85 $X2=0.26
+ $Y2=0.755
cc_70 N_A_M1003_g N_A_27_115#_c_148_n 0.0160984f $X=0.475 $Y=0.85 $X2=0.525
+ $Y2=1.455
cc_71 N_A_c_69_n N_A_27_115#_c_148_n 0.00117122f $X=0.475 $Y=2.285 $X2=0.525
+ $Y2=1.455
cc_72 N_A_c_70_n N_A_27_115#_c_148_n 2.65873e-19 $X=0.27 $Y=2.285 $X2=0.525
+ $Y2=1.455
cc_73 N_A_c_69_n N_A_27_115#_c_149_n 0.00133457f $X=0.475 $Y=2.285 $X2=0.345
+ $Y2=1.455
cc_74 N_A_c_70_n N_A_27_115#_c_149_n 0.0055861f $X=0.27 $Y=2.285 $X2=0.345
+ $Y2=1.455
cc_75 N_A_M1003_g N_A_27_115#_c_152_n 0.00322084f $X=0.475 $Y=0.85 $X2=0.61
+ $Y2=1.455
cc_76 N_A_M1003_g N_A_27_115#_c_153_n 0.0265302f $X=0.475 $Y=0.85 $X2=0.65
+ $Y2=3.065
cc_77 N_A_M1000_g N_A_27_115#_c_153_n 0.0140172f $X=0.475 $Y=3.235 $X2=0.65
+ $Y2=3.065
cc_78 N_A_c_69_n N_A_27_115#_c_153_n 0.00766302f $X=0.475 $Y=2.285 $X2=0.65
+ $Y2=3.065
cc_79 N_A_c_70_n N_A_27_115#_c_153_n 0.0456533f $X=0.27 $Y=2.285 $X2=0.65
+ $Y2=3.065
cc_80 A N_A_27_115#_c_153_n 0.00758489f $X=0.275 $Y=2.85 $X2=0.65 $Y2=3.065
cc_81 N_A_M1000_g N_A_27_115#_c_174_n 0.00865855f $X=0.475 $Y=3.235 $X2=0.65
+ $Y2=3.235
cc_82 N_B_M1002_g N_A_27_115#_M1001_g 0.0269401f $X=0.835 $Y=0.85 $X2=1.335
+ $Y2=0.85
cc_83 N_B_M1002_g N_A_27_115#_c_142_n 0.0104742f $X=0.835 $Y=0.85 $X2=1.37
+ $Y2=1.62
cc_84 N_B_M1004_g N_A_27_115#_c_143_n 0.00773101f $X=0.905 $Y=3.235 $X2=1.352
+ $Y2=2.33
cc_85 N_B_c_103_n N_A_27_115#_c_143_n 0.0206104f $X=0.95 $Y=1.945 $X2=1.352
+ $Y2=2.33
cc_86 N_B_c_104_n N_A_27_115#_c_143_n 0.0033451f $X=0.95 $Y=1.945 $X2=1.352
+ $Y2=2.33
cc_87 N_B_M1004_g N_A_27_115#_c_144_n 0.0381253f $X=0.905 $Y=3.235 $X2=1.352
+ $Y2=2.48
cc_88 N_B_c_104_n N_A_27_115#_c_144_n 0.00156524f $X=0.95 $Y=1.945 $X2=1.352
+ $Y2=2.48
cc_89 B N_A_27_115#_c_144_n 0.0037561f $X=0.955 $Y=2.48 $X2=1.352 $Y2=2.48
cc_90 N_B_M1002_g N_A_27_115#_c_150_n 0.0182215f $X=0.835 $Y=0.85 $X2=1.43
+ $Y2=1.455
cc_91 N_B_c_103_n N_A_27_115#_c_150_n 0.00258465f $X=0.95 $Y=1.945 $X2=1.43
+ $Y2=1.455
cc_92 N_B_c_104_n N_A_27_115#_c_150_n 0.0101796f $X=0.95 $Y=1.945 $X2=1.43
+ $Y2=1.455
cc_93 N_B_M1002_g N_A_27_115#_c_153_n 0.00755919f $X=0.835 $Y=0.85 $X2=0.65
+ $Y2=3.065
cc_94 N_B_M1004_g N_A_27_115#_c_153_n 0.0133197f $X=0.905 $Y=3.235 $X2=0.65
+ $Y2=3.065
cc_95 N_B_c_104_n N_A_27_115#_c_153_n 0.0541375f $X=0.95 $Y=1.945 $X2=0.65
+ $Y2=3.065
cc_96 B N_A_27_115#_c_153_n 0.00866797f $X=0.955 $Y=2.48 $X2=0.65 $Y2=3.065
cc_97 B N_A_27_115#_c_174_n 0.00286715f $X=0.955 $Y=2.48 $X2=0.65 $Y2=3.235
cc_98 N_B_c_104_n N_Y_c_211_n 0.0153635f $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_99 B N_Y_c_211_n 0.00659455f $X=0.955 $Y=2.48 $X2=1.55 $Y2=2.11
cc_100 N_B_M1002_g Y 6.71108e-19 $X=0.835 $Y=0.85 $X2=1.555 $Y2=1.74
cc_101 N_B_c_104_n Y 0.00695761f $X=0.95 $Y=1.945 $X2=1.555 $Y2=1.74
cc_102 N_B_M1002_g N_Y_c_213_n 7.71626e-19 $X=0.835 $Y=0.85 $X2=1.55 $Y2=1
cc_103 N_B_c_103_n N_Y_c_215_n 5.70769e-19 $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_104 N_B_c_104_n N_Y_c_215_n 0.00532157f $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_105 N_A_27_115#_M1001_g N_Y_c_208_n 0.00358423f $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=0.755
cc_106 N_A_27_115#_c_142_n N_Y_c_208_n 0.00166765f $X=1.37 $Y=1.62 $X2=1.55
+ $Y2=0.755
cc_107 N_A_27_115#_c_150_n N_Y_c_208_n 0.00508629f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_108 N_A_27_115#_c_142_n N_Y_c_211_n 0.00125776f $X=1.37 $Y=1.62 $X2=1.55
+ $Y2=2.11
cc_109 N_A_27_115#_c_143_n N_Y_c_211_n 0.0115869f $X=1.352 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_110 N_A_27_115#_c_144_n N_Y_c_211_n 0.00731267f $X=1.352 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_111 N_A_27_115#_c_150_n N_Y_c_211_n 0.00273485f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_112 N_A_27_115#_M1001_g Y 0.00406656f $X=1.335 $Y=0.85 $X2=1.555 $Y2=1.74
cc_113 N_A_27_115#_c_142_n Y 0.00711756f $X=1.37 $Y=1.62 $X2=1.555 $Y2=1.74
cc_114 N_A_27_115#_c_143_n Y 0.00892438f $X=1.352 $Y=2.33 $X2=1.555 $Y2=1.74
cc_115 N_A_27_115#_c_150_n Y 0.0152626f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_116 N_A_27_115#_M1001_g N_Y_c_213_n 0.00579788f $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=1
cc_117 N_A_27_115#_c_142_n N_Y_c_213_n 0.00154864f $X=1.37 $Y=1.62 $X2=1.55
+ $Y2=1
cc_118 N_A_27_115#_c_150_n N_Y_c_213_n 0.00238892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1
cc_119 N_A_27_115#_c_142_n N_Y_c_215_n 4.58687e-19 $X=1.37 $Y=1.62 $X2=1.55
+ $Y2=2.11
cc_120 N_A_27_115#_c_143_n N_Y_c_215_n 0.00721849f $X=1.352 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_121 N_A_27_115#_c_150_n N_Y_c_215_n 0.00181779f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
