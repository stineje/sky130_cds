* File: sky130_osu_sc_15T_hs__dffsr_1.spice
* Created: Fri Nov 12 14:29:44 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__dffsr_1.pex.spice"
.subckt sky130_osu_sc_15T_hs__dffsr_1  GND VDD RN SN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* RN	RN
* VDD	VDD
* GND	GND
MM1019 N_A_110_115#_M1019_d N_RN_M1019_g N_GND_M1019_s N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1034 N_A_217_565#_M1034_d N_A_110_115#_M1034_g N_GND_M1034_s N_GND_M1019_b
+ NLOWVT L=0.15 W=0.42 AD=0.0796811 AS=0.1113 PD=0.776604 PS=1.37 NRD=17.136
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1016 A_400_115# N_SN_M1016_g N_A_217_565#_M1034_d N_GND_M1019_b NLOWVT L=0.15
+ W=0.64 AD=0.0672 AS=0.121419 PD=0.85 PS=1.1834 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75000.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_GND_M1001_d N_A_432_468#_M1001_g A_400_115# N_GND_M1019_b NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 A_662_115# N_D_M1004_g N_GND_M1004_s N_GND_M1019_b NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1035 N_A_432_468#_M1035_d N_A_704_89#_M1035_g A_662_115# N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.144 AS=0.0672 PD=1.09 PS=0.85 NRD=15.936 NRS=9.372 M=1
+ R=4.26667 SA=75000.6 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1029 A_854_115# N_CK_M1029_g N_A_432_468#_M1035_d N_GND_M1019_b NLOWVT L=0.15
+ W=0.64 AD=0.0672 AS=0.144 PD=0.85 PS=1.09 NRD=9.372 NRS=15.936 M=1 R=4.26667
+ SA=75001.1 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1025 N_GND_M1025_d N_A_217_565#_M1025_g A_854_115# N_GND_M1019_b NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75001.5 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1028 A_1012_115# N_A_217_565#_M1028_g N_GND_M1025_d N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=9.372 NRS=0 M=1
+ R=4.26667 SA=75001.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_1084_115#_M1026_d N_CK_M1026_g A_1012_115# N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.144 AS=0.0672 PD=1.09 PS=0.85 NRD=15.936 NRS=9.372 M=1
+ R=4.26667 SA=75002.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1020 A_1204_115# N_A_704_89#_M1020_g N_A_1084_115#_M1026_d N_GND_M1019_b
+ NLOWVT L=0.15 W=0.64 AD=0.0672 AS=0.144 PD=0.85 PS=1.09 NRD=9.372 NRS=15.936
+ M=1 R=4.26667 SA=75002.9 SB=75001 A=0.096 P=1.58 MULT=1
MM1005 N_GND_M1005_d N_A_1246_89#_M1005_g A_1204_115# N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=9.372 M=1
+ R=4.26667 SA=75003.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_704_89#_M1008_d N_CK_M1008_g N_GND_M1005_d N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 A_1552_115# N_A_1084_115#_M1009_g N_GND_M1009_s N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1002 N_A_1246_89#_M1002_d N_SN_M1002_g A_1552_115# N_GND_M1019_b NLOWVT L=0.15
+ W=0.64 AD=0.121419 AS=0.0672 PD=1.1834 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1027 N_GND_M1027_d N_A_110_115#_M1027_g N_A_1246_89#_M1002_d N_GND_M1019_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0796811 PD=1.37 PS=0.776604 NRD=0
+ NRS=17.136 M=1 R=2.8 SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_GND_M1006_d N_A_1246_89#_M1006_g N_QN_M1006_s N_GND_M1019_b NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_Q_M1007_d N_QN_M1007_g N_GND_M1006_d N_GND_M1019_b NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_110_115#_M1023_d N_RN_M1023_g N_VDD_M1023_s N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1022 N_A_300_565#_M1022_d N_A_110_115#_M1022_g N_A_217_565#_M1022_s
+ N_VDD_M1023_b PSHORT L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0
+ M=1 R=13.3333 SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1010 N_VDD_M1010_d N_SN_M1010_g N_A_300_565#_M1022_d N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1011 N_A_300_565#_M1011_d N_A_432_468#_M1011_g N_VDD_M1010_d N_VDD_M1023_b
+ PSHORT L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1013 A_662_565# N_D_M1013_g N_VDD_M1013_s N_VDD_M1023_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75003.7 A=0.3 P=4.3 MULT=1
MM1000 N_A_432_468#_M1000_d N_CK_M1000_g A_662_565# N_VDD_M1023_b PSHORT L=0.15
+ W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75000.5 SB=75003.3 A=0.3 P=4.3 MULT=1
MM1033 A_854_565# N_A_704_89#_M1033_g N_A_432_468#_M1000_d N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75001.1 SB=75002.7 A=0.3 P=4.3 MULT=1
MM1030 N_VDD_M1030_d N_A_217_565#_M1030_g A_854_565# N_VDD_M1023_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001.5
+ SB=75002.4 A=0.3 P=4.3 MULT=1
MM1032 A_1012_565# N_A_217_565#_M1032_g N_VDD_M1030_d N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333
+ SA=75001.9 SB=75001.9 A=0.3 P=4.3 MULT=1
MM1031 N_A_1084_115#_M1031_d N_A_704_89#_M1031_g A_1012_565# N_VDD_M1023_b
+ PSHORT L=0.15 W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1
+ R=13.3333 SA=75002.3 SB=75001.6 A=0.3 P=4.3 MULT=1
MM1024 A_1204_565# N_CK_M1024_g N_A_1084_115#_M1031_d N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75002.9 SB=75001 A=0.3 P=4.3 MULT=1
MM1014 N_VDD_M1014_d N_A_1246_89#_M1014_g A_1204_565# N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333
+ SA=75003.3 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1018 N_A_704_89#_M1018_d N_CK_M1018_g N_VDD_M1014_d N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.7 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1021 N_VDD_M1021_d N_A_1084_115#_M1021_g N_A_1469_565#_M1021_s N_VDD_M1023_b
+ PSHORT L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1003 N_A_1469_565#_M1003_d N_SN_M1003_g N_VDD_M1021_d N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1012 N_A_1246_89#_M1012_d N_A_110_115#_M1012_g N_A_1469_565#_M1003_d
+ N_VDD_M1023_b PSHORT L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0
+ M=1 R=13.3333 SA=75001 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1015 N_VDD_M1015_d N_A_1246_89#_M1015_g N_QN_M1015_s N_VDD_M1023_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1017 N_Q_M1017_d N_QN_M1017_g N_VDD_M1015_d N_VDD_M1023_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX36_noxref N_GND_M1019_b N_VDD_M1023_b NWDIODE A=30.975 P=26.9
pX37_noxref noxref_27 RN RN PROBETYPE=1
pX38_noxref noxref_28 D D PROBETYPE=1
pX39_noxref noxref_29 CK CK PROBETYPE=1
pX40_noxref noxref_30 SN SN PROBETYPE=1
pX41_noxref noxref_31 QN QN PROBETYPE=1
pX42_noxref noxref_32 Q Q PROBETYPE=1
c_1971 A_1012_565# 0 1.57671e-19 $X=5.06 $Y=2.825
*
.include "sky130_osu_sc_15T_hs__dffsr_1.pxi.spice"
*
.ends
*
*
