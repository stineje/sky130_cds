* File: sky130_osu_sc_12T_hs__dff_l.pex.spice
* Created: Fri Nov 12 15:09:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%GND 1 2 3 4 5 81 83 91 93 103 105 115 117
+ 124 126 133 152 154
c181 115 0 1.61426e-19 $X=4.215 $Y=0.755
c182 81 0 1.27355e-19 $X=-0.045 $Y=0
r183 152 154 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r184 131 133 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.545 $Y=0.305
+ $X2=6.545 $Y2=0.74
r185 122 124 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.165 $Y=0.305
+ $X2=5.165 $Y2=0.755
r186 118 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.152
+ $X2=4.215 $Y2=0.152
r187 113 141 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.152
r188 113 115 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.755
r189 105 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.152
+ $X2=4.215 $Y2=0.152
r190 101 103 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.465 $Y=0.305
+ $X2=2.465 $Y2=0.74
r191 94 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.152
+ $X2=0.715 $Y2=0.152
r192 89 137 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.152
r193 89 91 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.755
r194 83 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.152
+ $X2=0.715 $Y2=0.152
r195 81 154 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r196 81 152 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r197 81 131 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.545 $Y2=0.305
r198 81 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.46 $Y2=0.152
r199 81 122 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.165 $Y2=0.305
r200 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.08 $Y2=0.152
r201 81 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.25 $Y2=0.152
r202 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.465 $Y2=0.305
r203 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.38 $Y2=0.152
r204 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.55 $Y2=0.152
r205 81 126 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.46 $Y2=0.152
r206 81 127 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.25 $Y2=0.152
r207 81 117 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=5.08 $Y2=0.152
r208 81 118 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.3 $Y2=0.152
r209 81 105 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.13 $Y2=0.152
r210 81 106 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.55 $Y2=0.152
r211 81 93 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.38 $Y2=0.152
r212 81 94 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.8 $Y2=0.152
r213 81 83 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.63 $Y2=0.152
r214 5 133 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.405
+ $Y=0.575 $X2=6.545 $Y2=0.74
r215 4 124 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.575 $X2=5.165 $Y2=0.755
r216 3 115 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.575 $X2=4.215 $Y2=0.755
r217 2 103 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.74
r218 1 91 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.575 $X2=0.715 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%VDD 1 2 3 4 5 61 63 70 72 80 82 90 92 98
+ 100 106 117 120 124
c104 70 0 5.41559e-20 $X=0.715 $Y=3.295
c105 1 0 1.59851e-19 $X=0.575 $Y=2.605
r106 120 124 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=6.46 $Y2=4.287
r107 117 124 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=4.25
+ $X2=6.46 $Y2=4.25
r108 104 117 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=4.135
+ $X2=6.545 $Y2=4.287
r109 104 106 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.545 $Y=4.135
+ $X2=6.545 $Y2=3.615
r110 101 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.25 $Y=4.287
+ $X2=5.165 $Y2=4.287
r111 101 103 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.25 $Y=4.287
+ $X2=5.78 $Y2=4.287
r112 100 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=4.287
+ $X2=6.545 $Y2=4.287
r113 100 103 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.46 $Y=4.287
+ $X2=5.78 $Y2=4.287
r114 96 115 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.165 $Y=4.135
+ $X2=5.165 $Y2=4.287
r115 96 98 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.165 $Y=4.135
+ $X2=5.165 $Y2=3.295
r116 93 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=4.287
+ $X2=4.215 $Y2=4.287
r117 93 95 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.3 $Y=4.287
+ $X2=4.42 $Y2=4.287
r118 92 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=4.287
+ $X2=5.165 $Y2=4.287
r119 92 95 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.08 $Y=4.287
+ $X2=4.42 $Y2=4.287
r120 88 113 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.215 $Y=4.135
+ $X2=4.215 $Y2=4.287
r121 88 90 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.215 $Y=4.135
+ $X2=4.215 $Y2=3.21
r122 85 87 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=4.287
+ $X2=3.74 $Y2=4.287
r123 83 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=4.287
+ $X2=2.465 $Y2=4.287
r124 83 85 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=2.55 $Y=4.287
+ $X2=3.06 $Y2=4.287
r125 82 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=4.287
+ $X2=4.215 $Y2=4.287
r126 82 87 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=4.13 $Y=4.287
+ $X2=3.74 $Y2=4.287
r127 78 112 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.465 $Y=4.135
+ $X2=2.465 $Y2=4.287
r128 78 80 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.465 $Y=4.135
+ $X2=2.465 $Y2=3.295
r129 75 77 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r130 73 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=4.287
+ $X2=0.715 $Y2=4.287
r131 73 75 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=0.8 $Y=4.287
+ $X2=1.02 $Y2=4.287
r132 72 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=4.287
+ $X2=2.465 $Y2=4.287
r133 72 77 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=4.287
+ $X2=1.7 $Y2=4.287
r134 68 110 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=4.287
r135 68 70 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=3.295
r136 65 120 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r137 63 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=4.287
+ $X2=0.715 $Y2=4.287
r138 63 65 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.63 $Y=4.287
+ $X2=0.34 $Y2=4.287
r139 61 117 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=4.135 $X2=6.46 $Y2=4.22
r140 61 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=4.135 $X2=5.78 $Y2=4.22
r141 61 115 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=4.135 $X2=5.1 $Y2=4.22
r142 61 95 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=4.135 $X2=4.42 $Y2=4.22
r143 61 87 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r144 61 85 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r145 61 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r146 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r147 61 75 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r148 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r149 5 106 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=3.025 $X2=6.545 $Y2=3.615
r150 4 98 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=2.605 $X2=5.165 $Y2=3.295
r151 3 90 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=4.075
+ $Y=2.605 $X2=4.215 $Y2=3.21
r152 2 80 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=2.605 $X2=2.465 $Y2=3.295
r153 1 70 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.605 $X2=0.715 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%A_75_248# 1 3 13 16 18 19 21 22 27 28 29
+ 30 31 33 36 41 42 44
c89 27 0 1.59851e-19 $X=0.625 $Y=2.62
c90 21 0 5.41559e-20 $X=0.51 $Y=2.285
r91 44 46 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=1.49 $Y=0.755 $X2=1.59
+ $Y2=0.755
r92 41 43 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.285
+ $X2=0.567 $Y2=2.45
r93 41 42 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.285
+ $X2=0.567 $Y2=2.12
r94 36 38 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=1.59 $Y=2.955
+ $X2=1.59 $Y2=3.635
r95 34 36 2.03372 $w=3.38e-07 $l=6e-08 $layer=LI1_cond $X=1.59 $Y=2.895 $X2=1.59
+ $Y2=2.955
r96 32 44 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.49 $Y=0.935
+ $X2=1.49 $Y2=0.755
r97 32 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.49 $Y=0.935
+ $X2=1.49 $Y2=1.2
r98 30 34 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=1.42 $Y=2.705
+ $X2=1.59 $Y2=2.895
r99 30 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.42 $Y=2.705
+ $X2=0.71 $Y2=2.705
r100 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.285
+ $X2=1.49 $Y2=1.2
r101 28 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.405 $Y=1.285
+ $X2=0.71 $Y2=1.285
r102 27 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=2.62
+ $X2=0.71 $Y2=2.705
r103 27 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.625 $Y=2.62
+ $X2=0.625 $Y2=2.45
r104 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.37
+ $X2=0.71 $Y2=1.285
r105 24 42 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.625 $Y=1.37
+ $X2=0.625 $Y2=2.12
r106 21 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=2.285 $X2=0.51 $Y2=2.285
r107 21 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.285
+ $X2=0.51 $Y2=2.45
r108 21 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.285
+ $X2=0.51 $Y2=2.12
r109 19 22 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.45 $Y=1.39
+ $X2=0.45 $Y2=2.12
r110 18 19 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.475 $Y=1.24
+ $X2=0.475 $Y2=1.39
r111 16 23 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.5 $Y=3.235
+ $X2=0.5 $Y2=2.45
r112 13 18 125.32 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.5 $Y=0.85 $X2=0.5
+ $Y2=1.24
r113 3 38 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.605 $X2=1.59 $Y2=3.635
r114 3 36 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.605 $X2=1.59 $Y2=2.955
r115 1 46 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.575 $X2=1.59 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%D 3 7 10 14 19
c43 19 0 1.36979e-19 $X=0.99 $Y=1.74
c44 10 0 1.98306e-19 $X=0.99 $Y=1.74
r45 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=1.74
+ $X2=0.99 $Y2=1.74
r46 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.74 $X2=0.99 $Y2=1.74
r47 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.74
+ $X2=0.99 $Y2=1.905
r48 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.74
+ $X2=0.99 $Y2=1.575
r49 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.93 $Y=3.235
+ $X2=0.93 $Y2=1.905
r50 3 11 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=0.93 $Y=0.85
+ $X2=0.93 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 67 70 71 72 73 80
c228 73 0 1.48522e-19 $X=3.725 $Y=2.11
c229 71 0 1.48522e-19 $X=1.495 $Y=2.11
c230 70 0 9.35091e-20 $X=3.435 $Y=2.11
c231 57 0 1.35605e-19 $X=4.575 $Y=2.11
c232 55 0 6.91727e-20 $X=3.185 $Y=2.11
c233 54 0 3.00693e-19 $X=3.465 $Y=2.11
c234 52 0 1.54708e-19 $X=3.1 $Y=1.4
c235 48 0 3.67809e-19 $X=1.83 $Y=1.4
c236 44 0 1.89329e-19 $X=1.745 $Y=2.11
c237 37 0 1.18241e-19 $X=3.55 $Y=2.285
c238 34 0 1.46493e-19 $X=3.1 $Y=1.235
c239 33 0 8.96132e-20 $X=3.1 $Y=1.4
c240 25 0 1.36979e-19 $X=1.38 $Y=2.285
r241 73 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.725 $Y=2.11
+ $X2=3.58 $Y2=2.11
r242 72 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.43 $Y=2.11
+ $X2=4.575 $Y2=2.11
r243 72 73 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=4.43 $Y=2.11
+ $X2=3.725 $Y2=2.11
r244 71 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.495 $Y=2.11
+ $X2=1.35 $Y2=2.11
r245 70 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.435 $Y=2.11
+ $X2=3.58 $Y2=2.11
r246 70 71 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=3.435 $Y=2.11
+ $X2=1.495 $Y2=2.11
r247 67 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.11
+ $X2=3.58 $Y2=2.11
r248 67 69 11.7308 $w=1.82e-07 $l=1.75e-07 $layer=LI1_cond $X=3.565 $Y=2.11
+ $X2=3.565 $Y2=2.285
r249 63 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.35 $Y=2.11
+ $X2=1.35 $Y2=2.11
r250 63 65 11.7308 $w=1.82e-07 $l=1.75e-07 $layer=LI1_cond $X=1.365 $Y=2.11
+ $X2=1.365 $Y2=2.285
r251 57 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.575 $Y=2.11
+ $X2=4.575 $Y2=2.11
r252 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.11
+ $X2=4.575 $Y2=2.285
r253 54 67 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.465 $Y=2.11 $X2=3.565
+ $Y2=2.11
r254 54 55 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.465 $Y=2.11
+ $X2=3.185 $Y2=2.11
r255 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.025
+ $X2=3.185 $Y2=2.11
r256 50 52 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.1 $Y=2.025
+ $X2=3.1 $Y2=1.4
r257 46 48 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.83 $Y=2.025
+ $X2=1.83 $Y2=1.4
r258 45 63 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.465 $Y=2.11 $X2=1.365
+ $Y2=2.11
r259 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=2.11
+ $X2=1.83 $Y2=2.025
r260 44 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.745 $Y=2.11
+ $X2=1.465 $Y2=2.11
r261 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=2.285 $X2=4.575 $Y2=2.285
r262 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=4.457 $Y=1.205
+ $X2=4.457 $Y2=1.355
r263 37 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=2.285 $X2=3.55 $Y2=2.285
r264 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=2.285
+ $X2=3.55 $Y2=2.45
r265 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.4 $X2=3.1 $Y2=1.4
r266 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.4 $X2=3.1
+ $Y2=1.235
r267 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.4 $X2=1.83 $Y2=1.4
r268 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.4
+ $X2=1.83 $Y2=1.235
r269 25 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.38
+ $Y=2.285 $X2=1.38 $Y2=2.285
r270 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=2.285
+ $X2=1.38 $Y2=2.45
r271 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=4.485 $Y=2.12
+ $X2=4.532 $Y2=2.285
r272 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.485 $Y=2.12
+ $X2=4.485 $Y2=1.355
r273 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=4.43 $Y=2.45
+ $X2=4.532 $Y2=2.285
r274 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=4.43 $Y=2.45
+ $X2=4.43 $Y2=3.235
r275 17 40 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.43 $Y=0.85
+ $X2=4.43 $Y2=1.205
r276 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.64 $Y=3.235
+ $X2=3.64 $Y2=2.45
r277 10 34 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.04 $Y=0.85
+ $X2=3.04 $Y2=1.235
r278 7 30 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.89 $Y=0.85
+ $X2=1.89 $Y2=1.235
r279 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.29 $Y=3.235
+ $X2=1.29 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%A_32_115# 1 3 11 15 17 18 21 22 27 31 34
+ 37 41 47 52 56 61 62 63 68
c115 61 0 8.96132e-20 $X=2.42 $Y=1.4
c116 47 0 1.5821e-19 $X=2.42 $Y=2.285
c117 31 0 6.36774e-20 $X=2.68 $Y=3.235
c118 27 0 1.54708e-19 $X=2.68 $Y=0.85
c119 22 0 1.89329e-19 $X=2.325 $Y=2.285
c120 21 0 6.91727e-20 $X=2.605 $Y=2.285
c121 15 0 6.36774e-20 $X=2.25 $Y=3.235
r122 63 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.43 $Y=1.37
+ $X2=0.285 $Y2=1.37
r123 62 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.185 $Y=1.37
+ $X2=2.33 $Y2=1.37
r124 62 63 1.68986 $w=1.7e-07 $l=1.755e-06 $layer=MET1_cond $X=2.185 $Y=1.37
+ $X2=0.43 $Y2=1.37
r125 59 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.33 $Y=1.37
+ $X2=2.33 $Y2=1.37
r126 59 61 5.43564 $w=2.02e-07 $l=9e-08 $layer=LI1_cond $X=2.33 $Y=1.345
+ $X2=2.42 $Y2=1.345
r127 54 56 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=2.78
+ $X2=0.285 $Y2=2.78
r128 52 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.285 $Y=1.37
+ $X2=0.285 $Y2=1.37
r129 49 52 4.81931 $w=2.73e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=1.317
+ $X2=0.285 $Y2=1.317
r130 45 61 1.74864 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.42 $Y=1.455
+ $X2=2.42 $Y2=1.345
r131 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.42 $Y=1.455
+ $X2=2.42 $Y2=2.285
r132 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.285 $Y=2.955
+ $X2=0.285 $Y2=3.635
r133 39 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.865
+ $X2=0.285 $Y2=2.78
r134 39 41 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.285 $Y=2.865
+ $X2=0.285 $Y2=2.955
r135 35 52 3.55113 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.285 $Y=1.18
+ $X2=0.285 $Y2=1.317
r136 35 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.285 $Y=1.18
+ $X2=0.285 $Y2=0.755
r137 34 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=2.695
+ $X2=0.17 $Y2=2.78
r138 33 49 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=1.317
r139 33 34 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=2.695
r140 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.68 $Y=2.42
+ $X2=2.68 $Y2=3.235
r141 25 27 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=2.68 $Y=1.265
+ $X2=2.68 $Y2=0.85
r142 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=2.285 $X2=2.42 $Y2=2.285
r143 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=2.285
+ $X2=2.42 $Y2=2.285
r144 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=2.285
+ $X2=2.68 $Y2=2.42
r145 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=2.285
+ $X2=2.42 $Y2=2.285
r146 20 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.4 $X2=2.42 $Y2=1.4
r147 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=1.4
+ $X2=2.42 $Y2=1.4
r148 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=1.4
+ $X2=2.68 $Y2=1.265
r149 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=1.4
+ $X2=2.42 $Y2=1.4
r150 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=2.42
+ $X2=2.325 $Y2=2.285
r151 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.25 $Y=2.42
+ $X2=2.25 $Y2=3.235
r152 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=1.265
+ $X2=2.325 $Y2=1.4
r153 9 11 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=2.25 $Y=1.265
+ $X2=2.25 $Y2=0.85
r154 3 43 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.605 $X2=0.285 $Y2=3.635
r155 3 41 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.605 $X2=0.285 $Y2=2.955
r156 1 37 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%A_243_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 50 54 59 63 67 70 74 75
c193 75 0 1.35605e-19 $X=4.5 $Y=1.74
c194 70 0 1.95058e-19 $X=3.725 $Y=1.725
c195 44 0 9.35091e-20 $X=3.58 $Y=1.74
c196 34 0 1.69503e-19 $X=1.41 $Y=1.28
c197 24 0 1.48522e-19 $X=3.04 $Y=3.235
c198 18 0 1.48522e-19 $X=1.89 $Y=3.235
r199 74 75 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.645 $Y=1.74
+ $X2=4.5 $Y2=1.74
r200 70 72 0.0981889 $w=2.26e-07 $l=1.52315e-07 $layer=MET1_cond $X=3.725
+ $Y=1.725 $X2=3.58 $Y2=1.74
r201 70 75 0.959157 $w=1.4e-07 $l=7.75e-07 $layer=MET1_cond $X=3.725 $Y=1.725
+ $X2=4.5 $Y2=1.725
r202 65 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=2.705
+ $X2=4.915 $Y2=2.705
r203 62 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.645 $Y=1.74
+ $X2=4.645 $Y2=1.74
r204 62 63 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=1.755
+ $X2=4.915 $Y2=1.755
r205 59 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.62
+ $X2=4.915 $Y2=2.705
r206 58 63 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.915 $Y=1.855
+ $X2=4.915 $Y2=1.755
r207 58 59 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.915 $Y=1.855
+ $X2=4.915 $Y2=2.62
r208 54 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.645 $Y=2.955
+ $X2=4.645 $Y2=3.635
r209 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=2.79
+ $X2=4.645 $Y2=2.705
r210 52 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=2.79
+ $X2=4.645 $Y2=2.955
r211 48 62 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.645 $Y=1.655
+ $X2=4.645 $Y2=1.755
r212 48 50 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.645 $Y=1.655
+ $X2=4.645 $Y2=0.755
r213 44 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=1.74
+ $X2=3.58 $Y2=1.74
r214 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.74 $X2=3.58 $Y2=1.74
r215 39 41 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=3.58 $Y=1.74
+ $X2=3.58 $Y2=1.85
r216 39 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.74
+ $X2=3.58 $Y2=1.575
r217 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.29 $Y=1.28
+ $X2=1.41 $Y2=1.28
r218 30 40 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=3.64 $Y=0.85
+ $X2=3.64 $Y2=1.575
r219 27 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.115 $Y=1.85
+ $X2=3.04 $Y2=1.85
r220 26 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.445 $Y=1.85
+ $X2=3.58 $Y2=1.85
r221 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.445 $Y=1.85
+ $X2=3.115 $Y2=1.85
r222 22 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.04 $Y=1.925
+ $X2=3.04 $Y2=1.85
r223 22 24 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=3.04 $Y=1.925
+ $X2=3.04 $Y2=3.235
r224 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=1.85
+ $X2=1.89 $Y2=1.85
r225 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.965 $Y=1.85
+ $X2=3.04 $Y2=1.85
r226 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.965 $Y=1.85
+ $X2=1.965 $Y2=1.85
r227 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=1.925
+ $X2=1.89 $Y2=1.85
r228 16 18 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=1.89 $Y=1.925
+ $X2=1.89 $Y2=3.235
r229 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=1.85
+ $X2=1.89 $Y2=1.85
r230 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.815 $Y=1.85
+ $X2=1.485 $Y2=1.85
r231 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.775
+ $X2=1.485 $Y2=1.85
r232 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.355
+ $X2=1.41 $Y2=1.28
r233 12 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.41 $Y=1.355
+ $X2=1.41 $Y2=1.775
r234 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.205
+ $X2=1.29 $Y2=1.28
r235 9 11 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=1.29 $Y=1.205
+ $X2=1.29 $Y2=0.85
r236 3 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.605 $X2=4.645 $Y2=3.635
r237 3 54 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.605 $X2=4.645 $Y2=2.955
r238 1 50 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.575 $X2=4.645 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%A_785_89# 1 3 11 15 17 21 25 28 31 32 35
+ 37 41 45 51 56 57 58 60 61 62 67
c167 67 0 7.28655e-20 $X=6.215 $Y=1.74
c168 61 0 1.62658e-19 $X=6.08 $Y=1.74
c169 35 0 1.61426e-19 $X=4.062 $Y=1.812
c170 11 0 1.35097e-19 $X=4 $Y=0.85
r171 61 67 0.0969593 $w=2.3e-07 $l=1.35e-07 $layer=MET1_cond $X=6.08 $Y=1.74
+ $X2=6.215 $Y2=1.74
r172 61 62 0.962882 $w=1.7e-07 $l=1e-06 $layer=MET1_cond $X=6.08 $Y=1.74
+ $X2=5.08 $Y2=1.74
r173 59 62 0.0704148 $w=1.7e-07 $l=1.15888e-07 $layer=MET1_cond $X=5.007
+ $Y=1.825 $X2=5.08 $Y2=1.74
r174 59 60 0.664026 $w=1.45e-07 $l=5.7e-07 $layer=MET1_cond $X=5.007 $Y=1.825
+ $X2=5.007 $Y2=2.395
r175 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.205 $Y=2.48
+ $X2=4.06 $Y2=2.48
r176 57 60 0.0704148 $w=1.7e-07 $l=1.15521e-07 $layer=MET1_cond $X=4.935 $Y=2.48
+ $X2=5.007 $Y2=2.395
r177 57 58 0.702904 $w=1.7e-07 $l=7.3e-07 $layer=MET1_cond $X=4.935 $Y=2.48
+ $X2=4.205 $Y2=2.48
r178 51 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=1.74
+ $X2=6.215 $Y2=1.74
r179 49 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=1.74
+ $X2=5.595 $Y2=1.74
r180 49 51 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.68 $Y=1.74
+ $X2=6.215 $Y2=1.74
r181 45 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.595 $Y=2.955
+ $X2=5.595 $Y2=3.635
r182 43 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.825
+ $X2=5.595 $Y2=1.74
r183 43 45 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=5.595 $Y=1.825
+ $X2=5.595 $Y2=2.955
r184 39 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.655
+ $X2=5.595 $Y2=1.74
r185 39 41 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.595 $Y=1.655
+ $X2=5.595 $Y2=0.755
r186 37 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.06 $Y=2.48
+ $X2=4.06 $Y2=2.48
r187 35 55 5.01943 $w=1.75e-07 $l=7.2e-08 $layer=LI1_cond $X=4.062 $Y=1.812
+ $X2=4.062 $Y2=1.74
r188 35 37 42.3356 $w=1.73e-07 $l=6.68e-07 $layer=LI1_cond $X=4.062 $Y=1.812
+ $X2=4.062 $Y2=2.48
r189 34 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.74 $X2=6.215 $Y2=1.74
r190 31 32 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=2.475
+ $X2=6.305 $Y2=2.625
r191 28 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.74 $X2=4.06 $Y2=1.74
r192 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.74
+ $X2=4.06 $Y2=1.905
r193 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.74
+ $X2=4.06 $Y2=1.575
r194 25 32 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.33 $Y=3.445
+ $X2=6.33 $Y2=2.625
r195 19 34 105.348 $w=2.27e-07 $l=5.12113e-07 $layer=POLY_cond $X=6.33 $Y=1.27
+ $X2=6.242 $Y2=1.74
r196 19 21 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.33 $Y=1.27
+ $X2=6.33 $Y2=0.785
r197 17 34 40.5863 $w=2.27e-07 $l=1.83016e-07 $layer=POLY_cond $X=6.28 $Y=1.905
+ $X2=6.242 $Y2=1.74
r198 17 31 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.28 $Y=1.905
+ $X2=6.28 $Y2=2.475
r199 15 30 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=4 $Y=3.235 $X2=4
+ $Y2=1.905
r200 11 29 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=4 $Y=0.85 $X2=4
+ $Y2=1.575
r201 3 47 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=2.605 $X2=5.595 $Y2=3.635
r202 3 45 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=2.605 $X2=5.595 $Y2=2.955
r203 1 41 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.575 $X2=5.595 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%A_623_115# 1 3 9 11 14 19 23 25 26 29 33
+ 36 40 43 44 45 46 53
c123 46 0 4.30668e-19 $X=3.585 $Y=1.37
c124 44 0 1.5821e-19 $X=2.905 $Y=1.37
c125 33 0 7.47985e-20 $X=3.44 $Y=1.34
c126 23 0 1.57671e-19 $X=2.76 $Y=1.37
r127 46 51 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=3.585
+ $Y=1.37 $X2=3.44 $Y2=1.34
r128 45 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.37
+ $X2=5.175 $Y2=1.37
r129 45 46 1.39137 $w=1.7e-07 $l=1.445e-06 $layer=MET1_cond $X=5.03 $Y=1.37
+ $X2=3.585 $Y2=1.37
r130 44 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.905 $Y=1.37
+ $X2=2.76 $Y2=1.37
r131 43 51 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=3.295
+ $Y=1.37 $X2=3.44 $Y2=1.34
r132 43 44 0.375524 $w=1.7e-07 $l=3.9e-07 $layer=MET1_cond $X=3.295 $Y=1.37
+ $X2=2.905 $Y2=1.37
r133 40 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.37
+ $X2=5.175 $Y2=1.37
r134 40 42 1.19608 $w=3.06e-07 $l=3e-08 $layer=LI1_cond $X=5.175 $Y=1.37
+ $X2=5.175 $Y2=1.4
r135 36 38 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=3.347 $Y=0.755
+ $X2=3.347 $Y2=1.035
r136 33 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.44 $Y=1.34
+ $X2=3.44 $Y2=1.34
r137 33 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.44 $Y=1.34
+ $X2=3.44 $Y2=1.035
r138 27 29 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=3.34 $Y=2.79
+ $X2=3.34 $Y2=3.295
r139 25 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=2.705
+ $X2=3.34 $Y2=2.79
r140 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=2.705
+ $X2=2.845 $Y2=2.705
r141 23 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.76 $Y=1.37
+ $X2=2.76 $Y2=1.37
r142 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=2.62
+ $X2=2.845 $Y2=2.705
r143 21 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.76 $Y=2.62
+ $X2=2.76 $Y2=1.37
r144 17 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.4 $X2=5.175 $Y2=1.4
r145 17 19 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.175 $Y=1.4
+ $X2=5.38 $Y2=1.4
r146 12 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.565
+ $X2=5.38 $Y2=1.4
r147 12 14 856.319 $w=1.5e-07 $l=1.67e-06 $layer=POLY_cond $X=5.38 $Y=1.565
+ $X2=5.38 $Y2=3.235
r148 9 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.235
+ $X2=5.38 $Y2=1.4
r149 9 11 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.38 $Y=1.235
+ $X2=5.38 $Y2=0.85
r150 3 29 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=3.115
+ $Y=2.605 $X2=3.34 $Y2=3.295
r151 1 36 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.575 $X2=3.34 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%ON 1 3 11 15 18 23 25 27 29 30 31 34 38
+ 41 43
c76 25 0 1.62658e-19 $X=6.115 $Y=2.195
c77 18 0 7.28655e-20 $X=6.7 $Y=2.015
r78 40 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.115 $Y=2.11
+ $X2=6.115 $Y2=2.11
r79 38 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.7 $Y=2.015 $X2=6.7
+ $Y2=1.745
r80 36 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.7 $Y=2.025 $X2=6.7
+ $Y2=2.015
r81 34 41 5.51377 $w=1.73e-07 $l=8.7e-08 $layer=LI1_cond $X=6.702 $Y=1.658
+ $X2=6.702 $Y2=1.745
r82 33 34 10.9642 $w=1.73e-07 $l=1.73e-07 $layer=LI1_cond $X=6.702 $Y=1.485
+ $X2=6.702 $Y2=1.658
r83 32 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=2.11 $X2=6.115
+ $Y2=2.11
r84 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=2.11
+ $X2=6.7 $Y2=2.025
r85 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=2.11
+ $X2=6.2 $Y2=2.11
r86 29 33 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=6.615 $Y=1.4
+ $X2=6.702 $Y2=1.485
r87 29 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=1.4
+ $X2=6.2 $Y2=1.4
r88 25 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=2.195
+ $X2=6.115 $Y2=2.11
r89 25 27 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=6.115 $Y=2.195
+ $X2=6.115 $Y2=3.615
r90 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=1.315
+ $X2=6.2 $Y2=1.4
r91 21 23 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.115 $Y=1.315
+ $X2=6.115 $Y2=0.74
r92 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=2.015 $X2=6.7 $Y2=2.015
r93 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.015
+ $X2=6.7 $Y2=2.18
r94 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.015
+ $X2=6.7 $Y2=1.85
r95 15 20 648.649 $w=1.5e-07 $l=1.265e-06 $layer=POLY_cond $X=6.76 $Y=3.445
+ $X2=6.76 $Y2=2.18
r96 11 19 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=6.76 $Y=0.785
+ $X2=6.76 $Y2=1.85
r97 3 27 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=3.025 $X2=6.115 $Y2=3.615
r98 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.575 $X2=6.115 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFF_L%Q 1 3 13 17 20 24 26 27 30 33
r26 28 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=1.07
+ $X2=7.09 $Y2=1.07
r27 26 27 18.6961 $w=1.73e-07 $l=2.95e-07 $layer=LI1_cond $X=6.972 $Y=2.88
+ $X2=6.972 $Y2=3.175
r28 22 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.97 $Y=2.48
+ $X2=6.97 $Y2=2.48
r29 22 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.97 $Y=2.48
+ $X2=7.09 $Y2=2.48
r30 20 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=2.395
+ $X2=7.09 $Y2=2.48
r31 19 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.155
+ $X2=7.09 $Y2=1.07
r32 19 20 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.09 $Y=1.155
+ $X2=7.09 $Y2=2.395
r33 17 27 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.975 $Y=3.615
+ $X2=6.975 $Y2=3.175
r34 11 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=0.985
+ $X2=6.975 $Y2=1.07
r35 11 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.975 $Y=0.985
+ $X2=6.975 $Y2=0.74
r36 9 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=2.565
+ $X2=6.97 $Y2=2.48
r37 9 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.97 $Y=2.565
+ $X2=6.97 $Y2=2.88
r38 3 17 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=6.835
+ $Y=3.025 $X2=6.975 $Y2=3.615
r39 1 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.575 $X2=6.975 $Y2=0.74
.ends

