magic
tech sky130A
magscale 1 2
timestamp 1606864598
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 374 1341
<< nmos >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
<< pmoshvt >>
rect 80 617 110 1217
rect 152 617 182 1217
rect 250 817 280 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 199 166 315
rect 110 131 121 199
rect 155 131 166 199
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 266 335 315
rect 282 131 293 266
rect 327 131 335 266
rect 282 115 335 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 617 152 1217
rect 182 1201 250 1217
rect 182 861 193 1201
rect 227 861 250 1201
rect 182 817 250 861
rect 280 1201 333 1217
rect 280 861 291 1201
rect 325 861 333 1201
rect 280 817 333 861
rect 182 617 235 817
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 199
rect 207 131 241 267
rect 293 131 327 266
<< pdiffc >>
rect 35 793 69 1201
rect 193 861 227 1201
rect 291 861 325 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 152 1217 182 1243
rect 250 1217 280 1243
rect 80 585 110 617
rect 56 569 110 585
rect 56 535 66 569
rect 100 535 110 569
rect 56 519 110 535
rect 56 370 86 519
rect 152 471 182 617
rect 136 461 202 471
rect 136 427 152 461
rect 186 427 202 461
rect 136 417 202 427
rect 56 340 110 370
rect 80 315 110 340
rect 166 315 196 417
rect 250 409 280 817
rect 250 393 306 409
rect 252 359 262 393
rect 296 359 306 393
rect 252 343 306 359
rect 252 315 282 343
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
<< polycont >>
rect 66 535 100 569
rect 152 427 186 461
rect 262 359 296 393
<< locali >>
rect 0 1311 374 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 374 1311
rect 35 1201 69 1217
rect 193 1201 227 1271
rect 193 845 227 861
rect 291 1201 325 1217
rect 35 751 69 793
rect 291 751 325 861
rect 35 717 325 751
rect 66 569 100 649
rect 66 519 100 535
rect 152 575 162 609
rect 152 461 186 575
rect 152 411 186 427
rect 223 393 257 501
rect 291 461 325 717
rect 223 359 262 393
rect 296 359 312 393
rect 35 267 241 301
rect 35 115 69 131
rect 121 199 155 215
rect 121 61 155 131
rect 207 115 241 131
rect 293 266 327 279
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 66 649 100 683
rect 162 575 196 609
rect 223 501 257 535
rect 291 427 325 461
rect 293 279 327 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 374 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 374 1311
rect 0 1271 374 1277
rect 54 683 112 689
rect 54 649 66 683
rect 100 649 134 683
rect 54 643 112 649
rect 150 609 208 615
rect 150 575 162 609
rect 196 575 230 609
rect 150 569 208 575
rect 211 535 269 541
rect 189 501 223 535
rect 257 501 269 535
rect 211 495 269 501
rect 279 461 337 467
rect 279 427 291 461
rect 325 427 337 461
rect 279 421 337 427
rect 293 319 327 421
rect 281 313 339 319
rect 281 279 293 313
rect 327 279 339 313
rect 281 273 339 279
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 83 666 83 666 1 A0
port 1 n
rlabel metal1 179 592 179 592 1 A1
port 2 n
rlabel metal1 308 444 308 444 1 Y
port 3 n
rlabel metal1 240 518 240 518 1 B0
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
