magic
tech sky130A
magscale 1 2
timestamp 1612372036
<< nwell >>
rect -9 529 288 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
<< ndiff >>
rect 27 228 80 243
rect 27 131 35 228
rect 69 131 80 228
rect 27 115 80 131
rect 110 228 166 243
rect 110 131 121 228
rect 155 131 166 228
rect 110 115 166 131
rect 196 228 249 243
rect 196 131 207 228
rect 241 131 249 228
rect 196 115 249 131
<< pdiff >>
rect 27 949 80 965
rect 27 609 35 949
rect 69 609 80 949
rect 27 565 80 609
rect 110 949 166 965
rect 110 745 121 949
rect 155 745 166 949
rect 110 565 166 745
rect 196 949 249 965
rect 196 609 207 949
rect 241 609 249 949
rect 196 565 249 609
<< ndiffc >>
rect 35 131 69 228
rect 121 131 155 228
rect 207 131 241 228
<< pdiffc >>
rect 35 609 69 949
rect 121 745 155 949
rect 207 609 241 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 80 477 110 565
rect 166 550 196 565
rect 166 520 251 550
rect 80 461 154 477
rect 80 427 110 461
rect 144 427 154 461
rect 80 411 154 427
rect 80 243 110 411
rect 221 368 251 520
rect 166 352 251 368
rect 166 318 176 352
rect 210 318 251 352
rect 166 302 251 318
rect 166 243 196 302
rect 80 89 110 115
rect 166 89 196 115
<< polycont >>
rect 110 427 144 461
rect 176 318 210 352
<< locali >>
rect 0 1089 286 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 286 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 729 155 745
rect 207 949 241 965
rect 35 352 69 609
rect 110 461 144 597
rect 207 557 241 609
rect 110 411 144 427
rect 176 352 210 368
rect 35 318 176 352
rect 35 228 69 318
rect 176 302 210 318
rect 35 115 69 131
rect 121 228 155 249
rect 121 61 155 131
rect 207 115 241 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 110 597 144 631
rect 207 523 241 557
rect 207 228 241 261
rect 207 227 241 228
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 286 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 286 1089
rect 0 1049 286 1055
rect 98 631 156 637
rect 64 597 110 631
rect 144 597 156 631
rect 98 591 156 597
rect 195 557 253 563
rect 195 523 207 557
rect 241 523 253 557
rect 195 517 253 523
rect 207 267 241 517
rect 195 261 253 267
rect 195 227 207 261
rect 241 227 253 261
rect 195 221 253 227
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 213 403 213 403 1 Y
port 2 n
rlabel viali 127 614 127 614 1 A
port 1 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
