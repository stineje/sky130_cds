magic
tech sky130A
magscale 1 2
timestamp 1612373916
<< nwell >>
rect -9 529 638 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 238 115 268 243
rect 358 115 388 243
rect 430 115 460 243
rect 516 115 546 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 238 565 268 965
rect 358 565 388 965
rect 430 565 460 965
rect 516 565 546 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 166 243
rect 110 131 121 215
rect 155 131 166 215
rect 110 115 166 131
rect 196 115 238 243
rect 268 215 358 243
rect 268 131 279 215
rect 347 131 358 215
rect 268 115 358 131
rect 388 115 430 243
rect 460 215 516 243
rect 460 131 471 215
rect 505 131 516 215
rect 460 115 516 131
rect 546 215 599 243
rect 546 131 557 215
rect 591 131 599 215
rect 546 115 599 131
<< pdiff >>
rect 27 949 80 965
rect 27 605 35 949
rect 69 605 80 949
rect 27 565 80 605
rect 110 949 166 965
rect 110 741 121 949
rect 155 741 166 949
rect 110 565 166 741
rect 196 565 238 965
rect 268 949 358 965
rect 268 605 279 949
rect 347 605 358 949
rect 268 565 358 605
rect 388 565 430 965
rect 460 949 516 965
rect 460 741 471 949
rect 505 741 516 949
rect 460 565 516 741
rect 546 949 599 965
rect 546 606 557 949
rect 591 606 599 949
rect 546 565 599 606
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 279 131 347 215
rect 471 131 505 215
rect 557 131 591 215
<< pdiffc >>
rect 35 605 69 949
rect 121 741 155 949
rect 279 605 347 949
rect 471 741 505 949
rect 557 606 591 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 238 965 268 991
rect 358 965 388 991
rect 430 965 460 991
rect 516 965 546 991
rect 80 550 110 565
rect 166 550 196 565
rect 70 520 196 550
rect 70 303 100 520
rect 142 518 196 520
rect 142 484 152 518
rect 186 484 196 518
rect 142 468 196 484
rect 142 410 196 426
rect 142 376 152 410
rect 186 376 196 410
rect 142 360 196 376
rect 70 278 110 303
rect 80 243 110 278
rect 166 243 196 360
rect 238 351 268 565
rect 358 534 388 565
rect 334 518 388 534
rect 430 550 460 565
rect 516 550 546 565
rect 430 520 546 550
rect 334 484 344 518
rect 378 484 388 518
rect 334 468 388 484
rect 479 518 546 520
rect 479 484 489 518
rect 523 484 546 518
rect 479 468 546 484
rect 420 409 474 425
rect 420 380 430 409
rect 358 375 430 380
rect 464 375 474 409
rect 238 335 292 351
rect 238 301 248 335
rect 282 301 292 335
rect 238 285 292 301
rect 358 350 474 375
rect 238 243 268 285
rect 358 243 388 350
rect 516 308 546 468
rect 430 278 546 308
rect 430 243 460 278
rect 516 243 546 278
rect 80 89 110 115
rect 166 89 196 115
rect 238 89 268 115
rect 358 89 388 115
rect 430 89 460 115
rect 516 89 546 115
<< polycont >>
rect 152 484 186 518
rect 152 376 186 410
rect 344 484 378 518
rect 489 484 523 518
rect 430 375 464 409
rect 248 301 282 335
<< locali >>
rect 0 1089 638 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 638 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 725 155 741
rect 279 949 347 965
rect 35 410 69 605
rect 152 597 200 631
rect 268 605 279 623
rect 471 949 505 1049
rect 471 725 505 741
rect 557 949 591 965
rect 152 518 186 597
rect 268 589 347 605
rect 136 484 152 518
rect 186 484 202 518
rect 268 483 302 589
rect 344 518 378 534
rect 344 410 378 484
rect 35 376 152 410
rect 186 376 378 410
rect 412 409 446 597
rect 489 518 523 523
rect 489 468 523 484
rect 35 215 69 376
rect 412 375 430 409
rect 464 375 480 409
rect 557 335 591 606
rect 232 301 248 335
rect 282 301 591 335
rect 35 115 69 131
rect 121 215 155 231
rect 121 61 155 131
rect 279 227 296 231
rect 330 227 347 231
rect 279 215 347 227
rect 279 115 347 131
rect 471 215 505 231
rect 471 61 505 131
rect 557 215 591 301
rect 557 115 591 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 638 61
rect 0 0 638 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 200 597 234 631
rect 412 597 446 631
rect 268 449 302 483
rect 489 523 523 557
rect 296 227 330 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1089 638 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 638 1089
rect 0 1049 638 1055
rect 188 631 246 637
rect 400 631 458 637
rect 188 597 200 631
rect 234 597 412 631
rect 446 597 458 631
rect 188 591 246 597
rect 400 591 458 597
rect 477 557 535 563
rect 455 523 489 557
rect 523 523 535 557
rect 477 517 535 523
rect 256 483 314 489
rect 256 449 268 483
rect 302 449 314 483
rect 256 443 314 449
rect 268 267 302 443
rect 268 261 342 267
rect 268 227 296 261
rect 330 227 342 261
rect 284 221 342 227
rect 0 55 638 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 638 55
rect 0 0 638 21
<< labels >>
rlabel viali 218 614 218 614 1 A
port 1 n
rlabel metal1 285 434 285 434 1 Y
port 2 n
rlabel viali 506 540 506 540 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
