* File: sky130_osu_sc_18T_ms__addf_l.spice
* Created: Fri Nov 12 13:59:49 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_ms__addf_l.pex.spice"
.subckt sky130_osu_sc_18T_ms__addf_l  GND VDD A B CI CON S CO
* 
* CO	CO
* S	S
* CON	CON
* CI	CI
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1010 N_GND_M1010_d N_A_M1010_g N_A_27_115#_M1010_s N_GND_M1010_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_27_115#_M1000_d N_B_M1000_g N_GND_M1010_d N_GND_M1010_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.7 A=0.15 P=2.3 MULT=1
MM1003 N_CON_M1003_d N_CI_M1003_g N_A_27_115#_M1000_d N_GND_M1010_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75004.3 A=0.15 P=2.3 MULT=1
MM1024 A_368_115# N_B_M1024_g N_CON_M1003_d N_GND_M1010_b NSHORT L=0.15 W=1
+ AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75003.9 A=0.15 P=2.3 MULT=1
MM1026 N_GND_M1026_d N_A_M1026_g A_368_115# N_GND_M1010_b NSHORT L=0.15 W=1
+ AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.8
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1019 N_A_526_115#_M1019_d N_A_M1019_g N_GND_M1026_d N_GND_M1010_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1022 N_GND_M1022_d N_B_M1022_g N_A_526_115#_M1019_d N_GND_M1010_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_526_115#_M1012_d N_CI_M1012_g N_GND_M1022_d N_GND_M1010_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.1 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_784_115#_M1014_d N_CON_M1014_g N_A_526_115#_M1012_d N_GND_M1010_b
+ NSHORT L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.6 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1016 A_870_115# N_B_M1016_g N_A_784_115#_M1014_d N_GND_M1010_b NSHORT L=0.15
+ W=1 AD=0.13 AS=0.14 PD=1.26 PS=1.28 NRD=8.988 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 A_952_115# N_CI_M1007_g A_870_115# N_GND_M1010_b NSHORT L=0.15 W=1
+ AD=0.13 AS=0.13 PD=1.26 PS=1.26 NRD=8.988 NRS=8.988 M=1 R=6.66667 SA=75004.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_GND_M1004_d N_A_M1004_g A_952_115# N_GND_M1010_b NSHORT L=0.15 W=1
+ AD=0.184195 AS=0.13 PD=1.54023 PS=1.26 NRD=0 NRS=8.988 M=1 R=6.66667
+ SA=75004.8 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_S_M1017_d N_A_784_115#_M1017_g N_GND_M1004_d N_GND_M1010_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.136305 PD=2.01 PS=1.13977 NRD=0 NRS=9.72 M=1
+ R=4.93333 SA=75005.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_CO_M1020_d N_CON_M1020_g N_GND_M1020_s N_GND_M1010_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VDD_M1011_d N_A_M1011_g N_A_27_617#_M1011_s N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75005.1 A=0.45 P=6.3 MULT=1
MM1001 N_A_27_617#_M1001_d N_B_M1001_g N_VDD_M1011_d N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75004.7
+ A=0.45 P=6.3 MULT=1
MM1006 N_CON_M1006_d N_CI_M1006_g N_A_27_617#_M1001_d N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001
+ SB=75004.3 A=0.45 P=6.3 MULT=1
MM1025 A_368_617# N_B_M1025_g N_CON_M1006_d N_VDD_M1011_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75001.5
+ SB=75003.8 A=0.45 P=6.3 MULT=1
MM1027 N_VDD_M1027_d N_A_M1027_g A_368_617# N_VDD_M1011_b PSHORT L=0.15 W=3
+ AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.8
+ SB=75003.5 A=0.45 P=6.3 MULT=1
MM1021 N_A_526_617#_M1021_d N_A_M1021_g N_VDD_M1027_d N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.3
+ SB=75003.1 A=0.45 P=6.3 MULT=1
MM1023 N_VDD_M1023_d N_B_M1023_g N_A_526_617#_M1021_d N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.7
+ SB=75002.6 A=0.45 P=6.3 MULT=1
MM1013 N_A_526_617#_M1013_d N_CI_M1013_g N_VDD_M1023_d N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.1
+ SB=75002.2 A=0.45 P=6.3 MULT=1
MM1015 N_A_784_115#_M1015_d N_CON_M1015_g N_A_526_617#_M1013_d N_VDD_M1011_b
+ PSHORT L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20
+ SA=75003.6 SB=75001.8 A=0.45 P=6.3 MULT=1
MM1018 A_870_617# N_B_M1018_g N_A_784_115#_M1015_d N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.39 AS=0.42 PD=3.26 PS=3.28 NRD=4.9053 NRS=0 M=1 R=20 SA=75004
+ SB=75001.3 A=0.45 P=6.3 MULT=1
MM1008 A_952_617# N_CI_M1008_g A_870_617# N_VDD_M1011_b PSHORT L=0.15 W=3
+ AD=0.39 AS=0.39 PD=3.26 PS=3.26 NRD=4.9053 NRS=4.9053 M=1 R=20 SA=75004.4
+ SB=75000.9 A=0.45 P=6.3 MULT=1
MM1005 N_VDD_M1005_d N_A_M1005_g A_952_617# N_VDD_M1011_b PSHORT L=0.15 W=3
+ AD=0.567 AS=0.39 PD=4.008 PS=3.26 NRD=0 NRS=4.9053 M=1 R=20 SA=75004.8
+ SB=75000.5 A=0.45 P=6.3 MULT=1
MM1002 N_S_M1002_d N_A_784_115#_M1002_g N_VDD_M1005_d N_VDD_M1011_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.378 PD=4.53 PS=2.672 NRD=0 NRS=5.9888 M=1 R=13.3333
+ SA=75005.3 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1009 N_CO_M1009_d N_CON_M1009_g N_VDD_M1009_s N_VDD_M1011_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX28_noxref N_GND_M1010_b N_VDD_M1011_b NWDIODE A=27.436 P=22.04
pX29_noxref noxref_20 A A PROBETYPE=1
pX30_noxref noxref_21 B B PROBETYPE=1
pX31_noxref noxref_22 CI CI PROBETYPE=1
pX32_noxref noxref_23 S S PROBETYPE=1
pX33_noxref noxref_24 CON CON PROBETYPE=1
pX34_noxref noxref_25 CO CO PROBETYPE=1
*
.include "sky130_osu_sc_18T_ms__addf_l.pxi.spice"
*
.ends
*
*
