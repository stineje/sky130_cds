* File: sky130_osu_sc_15T_hs__tnbufi_l.pxi.spice
* Created: Fri Nov 12 14:33:55 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_6_p
+ N_GND_c_2_p GND N_GND_c_3_p PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%GND
x_PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_33_p
+ N_VDD_c_38_p N_VDD_c_42_p VDD N_VDD_c_34_p
+ PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%VDD
x_PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_c_57_n N_A_27_115#_c_58_n
+ N_A_27_115#_c_61_n N_A_27_115#_c_62_n N_A_27_115#_c_63_n N_A_27_115#_c_64_n
+ PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%A_27_115#
x_PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%OE N_OE_M1002_g N_OE_c_101_n N_OE_M1001_g
+ N_OE_M1005_g N_OE_c_102_n N_OE_c_103_n OE PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%OE
x_PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%A N_A_M1004_g N_A_M1003_g N_A_c_146_n
+ N_A_c_147_n N_A_c_148_n A PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%A
x_PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%Y N_Y_M1004_d N_Y_M1003_d N_Y_c_190_n
+ N_Y_c_192_n Y N_Y_c_194_n N_Y_c_195_n PM_SKY130_OSU_SC_15T_HS__TNBUFI_L%Y
cc_1 N_GND_M1002_b N_A_27_115#_M1000_g 0.0501862f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.85
cc_2 N_GND_c_2_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905
+ $Y2=0.85
cc_3 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=0.85
cc_4 N_GND_M1002_b N_A_27_115#_c_57_n 0.0434193f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=1.915
cc_5 N_GND_M1002_b N_A_27_115#_c_58_n 0.0286712f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_6 N_GND_c_6_p N_A_27_115#_c_58_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_7 N_GND_c_3_p N_A_27_115#_c_58_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_8 N_GND_M1002_b N_A_27_115#_c_61_n 0.0221237f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=4.225
cc_9 N_GND_M1002_b N_A_27_115#_c_62_n 0.00872418f $X=-0.045 $Y=0 $X2=0.605
+ $Y2=1.915
cc_10 N_GND_M1002_b N_A_27_115#_c_63_n 0.00647094f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.915
cc_11 N_GND_M1002_b N_A_27_115#_c_64_n 0.00739462f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=1.915
cc_12 N_GND_M1002_b N_OE_M1002_g 0.0293808f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_13 N_GND_c_6_p N_OE_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.85
cc_14 N_GND_c_2_p N_OE_M1002_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.85
cc_15 N_GND_c_3_p N_OE_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.85
cc_16 N_GND_M1002_b N_OE_c_101_n 0.102331f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.75
cc_17 N_GND_M1002_b N_OE_c_102_n 0.0253119f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.465
cc_18 N_GND_M1002_b N_OE_c_103_n 0.00123196f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.505
cc_19 N_GND_M1002_b OE 5.10551e-19 $X=-0.045 $Y=0 $X2=0.69 $Y2=2.7
cc_20 N_GND_M1002_b N_A_M1004_g 0.0556043f $X=-0.045 $Y=0 $X2=1.265 $Y2=0.85
cc_21 N_GND_c_3_p N_A_M1004_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.265 $Y2=0.85
cc_22 N_GND_M1002_b N_A_M1003_g 0.0426097f $X=-0.045 $Y=0 $X2=1.265 $Y2=4.195
cc_23 N_GND_M1002_b N_A_c_146_n 0.031953f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.83
cc_24 N_GND_M1002_b N_A_c_147_n 0.0125638f $X=-0.045 $Y=0 $X2=1.14 $Y2=3.07
cc_25 N_GND_M1002_b N_A_c_148_n 0.00872469f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.83
cc_26 N_GND_M1002_b N_Y_c_190_n 0.0164997f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.74
cc_27 N_GND_c_3_p N_Y_c_190_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.48 $Y2=0.74
cc_28 N_GND_M1002_b N_Y_c_192_n 0.0151339f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.33
cc_29 N_GND_M1002_b Y 0.0395158f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.56
cc_30 N_GND_M1002_b N_Y_c_194_n 0.0122638f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.22
cc_31 N_GND_M1002_b N_Y_c_195_n 0.0157299f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.33
cc_32 N_VDD_M1001_b N_A_27_115#_c_61_n 0.0438222f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=4.225
cc_33 N_VDD_c_33_p N_A_27_115#_c_61_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=4.225
cc_34 N_VDD_c_34_p N_A_27_115#_c_61_n 0.00435496f $X=1.02 $Y=5.36 $X2=0.26
+ $Y2=4.225
cc_35 N_VDD_M1001_b N_OE_c_101_n 0.0237235f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=2.75
cc_36 N_VDD_M1001_b N_OE_M1001_g 0.0588985f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=4.195
cc_37 N_VDD_c_33_p N_OE_M1001_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475
+ $Y2=4.195
cc_38 N_VDD_c_38_p N_OE_M1001_g 0.00362996f $X=0.69 $Y=4.225 $X2=0.475 $Y2=4.195
cc_39 N_VDD_c_34_p N_OE_M1001_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=4.195
cc_40 N_VDD_M1001_b N_OE_M1005_g 0.0498873f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=4.195
cc_41 N_VDD_c_38_p N_OE_M1005_g 0.00362996f $X=0.69 $Y=4.225 $X2=0.905 $Y2=4.195
cc_42 N_VDD_c_42_p N_OE_M1005_g 0.00496961f $X=1.02 $Y=5.33 $X2=0.905 $Y2=4.195
cc_43 N_VDD_c_34_p N_OE_M1005_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.905 $Y2=4.195
cc_44 N_VDD_M1001_b N_OE_c_103_n 0.00252354f $X=-0.045 $Y=2.645 $X2=0.69
+ $Y2=2.505
cc_45 N_VDD_M1001_b OE 0.0104205f $X=-0.045 $Y=2.645 $X2=0.69 $Y2=2.7
cc_46 N_VDD_M1001_b N_A_M1003_g 0.0605315f $X=-0.045 $Y=2.645 $X2=1.265
+ $Y2=4.195
cc_47 N_VDD_c_42_p N_A_M1003_g 0.00496961f $X=1.02 $Y=5.33 $X2=1.265 $Y2=4.195
cc_48 N_VDD_c_34_p N_A_M1003_g 0.00429146f $X=1.02 $Y=5.36 $X2=1.265 $Y2=4.195
cc_49 N_VDD_M1001_b N_A_c_147_n 0.00640673f $X=-0.045 $Y=2.645 $X2=1.14 $Y2=3.07
cc_50 N_VDD_M1001_b A 0.011498f $X=-0.045 $Y=2.645 $X2=1.14 $Y2=3.07
cc_51 N_VDD_M1001_b N_Y_c_192_n 0.045274f $X=-0.045 $Y=2.645 $X2=1.48 $Y2=2.33
cc_52 N_VDD_c_42_p N_Y_c_192_n 0.00477009f $X=1.02 $Y=5.33 $X2=1.48 $Y2=2.33
cc_53 N_VDD_c_34_p N_Y_c_192_n 0.00435496f $X=1.02 $Y=5.36 $X2=1.48 $Y2=2.33
cc_54 N_A_27_115#_M1000_g N_OE_M1002_g 0.0330955f $X=0.905 $Y=0.85 $X2=0.475
+ $Y2=0.85
cc_55 N_A_27_115#_c_58_n N_OE_M1002_g 0.0138858f $X=0.26 $Y=0.74 $X2=0.475
+ $Y2=0.85
cc_56 N_A_27_115#_M1000_g N_OE_c_101_n 0.00301188f $X=0.905 $Y=0.85 $X2=0.475
+ $Y2=2.75
cc_57 N_A_27_115#_c_57_n N_OE_c_101_n 0.0400875f $X=0.905 $Y=1.915 $X2=0.475
+ $Y2=2.75
cc_58 N_A_27_115#_c_58_n N_OE_c_101_n 0.0121188f $X=0.26 $Y=0.74 $X2=0.475
+ $Y2=2.75
cc_59 N_A_27_115#_c_61_n N_OE_c_101_n 0.04195f $X=0.26 $Y=4.225 $X2=0.475
+ $Y2=2.75
cc_60 N_A_27_115#_c_62_n N_OE_c_101_n 0.00111679f $X=0.605 $Y=1.915 $X2=0.475
+ $Y2=2.75
cc_61 N_A_27_115#_c_63_n N_OE_c_101_n 0.00632922f $X=0.26 $Y=1.915 $X2=0.475
+ $Y2=2.75
cc_62 N_A_27_115#_c_64_n N_OE_c_101_n 7.56328e-19 $X=0.69 $Y=1.915 $X2=0.475
+ $Y2=2.75
cc_63 N_A_27_115#_c_61_n N_OE_M1001_g 0.0411995f $X=0.26 $Y=4.225 $X2=0.475
+ $Y2=4.195
cc_64 N_A_27_115#_c_58_n N_OE_c_102_n 0.0104429f $X=0.26 $Y=0.74 $X2=0.475
+ $Y2=1.465
cc_65 N_A_27_115#_c_62_n N_OE_c_102_n 0.00711711f $X=0.605 $Y=1.915 $X2=0.475
+ $Y2=1.465
cc_66 N_A_27_115#_c_57_n N_OE_c_103_n 2.15234e-19 $X=0.905 $Y=1.915 $X2=0.69
+ $Y2=2.505
cc_67 N_A_27_115#_c_61_n N_OE_c_103_n 0.0193056f $X=0.26 $Y=4.225 $X2=0.69
+ $Y2=2.505
cc_68 N_A_27_115#_c_64_n N_OE_c_103_n 0.00847614f $X=0.69 $Y=1.915 $X2=0.69
+ $Y2=2.505
cc_69 N_A_27_115#_c_57_n OE 0.00125736f $X=0.905 $Y=1.915 $X2=0.69 $Y2=2.7
cc_70 N_A_27_115#_c_61_n OE 0.00651113f $X=0.26 $Y=4.225 $X2=0.69 $Y2=2.7
cc_71 N_A_27_115#_c_62_n OE 0.00158904f $X=0.605 $Y=1.915 $X2=0.69 $Y2=2.7
cc_72 N_A_27_115#_c_64_n OE 7.36678e-19 $X=0.69 $Y=1.915 $X2=0.69 $Y2=2.7
cc_73 N_A_27_115#_M1000_g N_A_M1004_g 0.0509405f $X=0.905 $Y=0.85 $X2=1.265
+ $Y2=0.85
cc_74 N_A_27_115#_c_57_n N_A_c_146_n 0.0509405f $X=0.905 $Y=1.915 $X2=1.325
+ $Y2=1.83
cc_75 N_A_27_115#_c_64_n N_A_c_146_n 2.55709e-19 $X=0.69 $Y=1.915 $X2=1.325
+ $Y2=1.83
cc_76 N_A_27_115#_c_57_n N_A_c_147_n 0.00134082f $X=0.905 $Y=1.915 $X2=1.14
+ $Y2=3.07
cc_77 N_A_27_115#_c_64_n N_A_c_147_n 0.00813625f $X=0.69 $Y=1.915 $X2=1.14
+ $Y2=3.07
cc_78 N_A_27_115#_M1000_g N_A_c_148_n 0.00160395f $X=0.905 $Y=0.85 $X2=1.325
+ $Y2=1.83
cc_79 N_A_27_115#_c_64_n N_A_c_148_n 0.00878007f $X=0.69 $Y=1.915 $X2=1.325
+ $Y2=1.83
cc_80 N_A_27_115#_c_61_n A 0.00539687f $X=0.26 $Y=4.225 $X2=1.14 $Y2=3.07
cc_81 N_A_27_115#_M1000_g Y 3.32545e-19 $X=0.905 $Y=0.85 $X2=1.525 $Y2=1.56
cc_82 N_A_27_115#_M1000_g N_Y_c_194_n 0.00101819f $X=0.905 $Y=0.85 $X2=1.48
+ $Y2=1.22
cc_83 N_OE_c_101_n N_A_M1003_g 0.151072f $X=0.475 $Y=2.75 $X2=1.265 $Y2=4.195
cc_84 N_OE_c_103_n N_A_M1003_g 4.61952e-19 $X=0.69 $Y=2.505 $X2=1.265 $Y2=4.195
cc_85 N_OE_c_101_n N_A_c_147_n 0.0110152f $X=0.475 $Y=2.75 $X2=1.14 $Y2=3.07
cc_86 N_OE_c_103_n N_A_c_147_n 0.0187675f $X=0.69 $Y=2.505 $X2=1.14 $Y2=3.07
cc_87 OE N_A_c_147_n 0.007197f $X=0.69 $Y=2.7 $X2=1.14 $Y2=3.07
cc_88 N_OE_M1001_g A 8.46663e-19 $X=0.475 $Y=4.195 $X2=1.14 $Y2=3.07
cc_89 N_OE_M1005_g A 0.0104662f $X=0.905 $Y=4.195 $X2=1.14 $Y2=3.07
cc_90 OE A 0.004991f $X=0.69 $Y=2.7 $X2=1.14 $Y2=3.07
cc_91 N_A_M1004_g N_Y_c_190_n 0.00971844f $X=1.265 $Y=0.85 $X2=1.48 $Y2=0.74
cc_92 N_A_c_146_n N_Y_c_190_n 8.70049e-19 $X=1.325 $Y=1.83 $X2=1.48 $Y2=0.74
cc_93 N_A_c_148_n N_Y_c_190_n 0.00231567f $X=1.325 $Y=1.83 $X2=1.48 $Y2=0.74
cc_94 N_A_M1003_g N_Y_c_192_n 0.0453863f $X=1.265 $Y=4.195 $X2=1.48 $Y2=2.33
cc_95 N_A_c_146_n N_Y_c_192_n 0.00102058f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
cc_96 N_A_c_147_n N_Y_c_192_n 0.0606572f $X=1.14 $Y=3.07 $X2=1.48 $Y2=2.33
cc_97 N_A_c_148_n N_Y_c_192_n 0.00330615f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
cc_98 A N_Y_c_192_n 0.00706656f $X=1.14 $Y=3.07 $X2=1.48 $Y2=2.33
cc_99 N_A_M1004_g Y 0.00768908f $X=1.265 $Y=0.85 $X2=1.525 $Y2=1.56
cc_100 N_A_M1003_g Y 0.00511826f $X=1.265 $Y=4.195 $X2=1.525 $Y2=1.56
cc_101 N_A_c_146_n Y 0.00539093f $X=1.325 $Y=1.83 $X2=1.525 $Y2=1.56
cc_102 N_A_c_147_n Y 0.012418f $X=1.14 $Y=3.07 $X2=1.525 $Y2=1.56
cc_103 N_A_c_148_n Y 0.0130872f $X=1.325 $Y=1.83 $X2=1.525 $Y2=1.56
cc_104 N_A_M1004_g N_Y_c_194_n 0.00707709f $X=1.265 $Y=0.85 $X2=1.48 $Y2=1.22
cc_105 N_A_c_146_n N_Y_c_194_n 0.00129509f $X=1.325 $Y=1.83 $X2=1.48 $Y2=1.22
cc_106 N_A_c_148_n N_Y_c_194_n 0.00203451f $X=1.325 $Y=1.83 $X2=1.48 $Y2=1.22
cc_107 N_A_M1003_g N_Y_c_195_n 0.00489736f $X=1.265 $Y=4.195 $X2=1.48 $Y2=2.33
cc_108 N_A_c_146_n N_Y_c_195_n 0.00138163f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
cc_109 N_A_c_147_n N_Y_c_195_n 0.00656407f $X=1.14 $Y=3.07 $X2=1.48 $Y2=2.33
cc_110 N_A_c_148_n N_Y_c_195_n 0.00227834f $X=1.325 $Y=1.83 $X2=1.48 $Y2=2.33
