* File: sky130_osu_sc_18T_hs__or2_1.pex.spice
* Created: Thu Oct 29 17:09:35 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__OR2_1%GND 1 2 15 19 23 31 32 34 37
r37 34 37 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r38 31 32 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r39 21 32 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r40 21 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r41 17 19 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r42 15 31 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r43 15 27 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r44 15 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r45 15 17 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r46 15 27 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r47 2 23 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r48 1 19 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_1%VDD 1 10 14 20 21 23 26
r23 30 33 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r24 26 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r25 23 26 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r26 20 33 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r27 20 21 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r28 14 17 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=5.835
r29 12 21 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r30 12 17 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r31 10 33 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r32 10 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r33 1 17 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r34 1 14 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_1%B 3 7 10 15 18
r28 16 18 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.675
+ $X2=0.475 $Y2=2.675
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.675 $X2=0.27 $Y2=2.675
r30 12 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.96
+ $X2=0.27 $Y2=2.675
r31 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.96
+ $X2=0.27 $Y2=2.96
r32 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.84
+ $X2=0.475 $Y2=2.675
r33 5 7 894.777 $w=1.5e-07 $l=1.745e-06 $layer=POLY_cond $X=0.475 $Y=2.84
+ $X2=0.475 $Y2=4.585
r34 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.51
+ $X2=0.475 $Y2=2.675
r35 1 3 735.819 $w=1.5e-07 $l=1.435e-06 $layer=POLY_cond $X=0.475 $Y=2.51
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_1%A 3 7 10 15 16
r44 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=2.55
r45 16 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.385
+ $X2=0.95 $Y2=2.22
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.385 $X2=0.95 $Y2=2.385
r47 12 15 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.95 $Y2=2.385
r48 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=3.33
+ $X2=0.95 $Y2=3.33
r49 7 18 1043.48 $w=1.5e-07 $l=2.035e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.55
r50 3 17 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.22
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_1%A_27_617# 1 2 9 13 14 16 17 20 24 25 27
+ 30 34 37
r70 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r71 32 37 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.935
+ $X2=0.65 $Y2=1.935
r72 32 34 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.935
+ $X2=1.43 $Y2=1.935
r73 28 37 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.65 $Y2=1.935
r74 28 30 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=0.825
r75 26 37 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.65 $Y2=1.935
r76 26 27 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r77 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.63
+ $X2=0.61 $Y2=3.545
r78 24 25 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.63
+ $X2=0.345 $Y2=3.63
r79 20 22 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.26 $Y=3.795
+ $X2=0.26 $Y2=5.835
r80 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.715
+ $X2=0.345 $Y2=3.63
r81 18 20 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=3.715 $X2=0.26
+ $Y2=3.795
r82 16 17 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.81
+ $X2=1.352 $Y2=2.96
r83 14 35 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.412 $Y2=1.935
r84 14 16 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1 $X2=1.37
+ $Y2=2.81
r85 13 17 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.96
r86 7 35 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.412 $Y2=1.935
r87 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r88 2 22 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r89 2 20 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.795
r90 1 30 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OR2_1%Y 1 2 10 13 17 18 21
r35 28 30 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r36 18 28 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r37 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r38 14 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r39 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r40 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r41 8 10 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r42 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r43 7 10 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r44 2 30 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r45 2 28 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r46 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

