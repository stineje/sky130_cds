* File: sky130_osu_sc_18T_ls__oai21_l.pxi.spice
* Created: Fri Nov 12 14:18:52 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%GND N_GND_M1005_d N_GND_M1005_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_LS__OAI21_L%GND
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%VDD N_VDD_M1003_d N_VDD_M1004_b N_VDD_c_39_p
+ N_VDD_c_45_p N_VDD_c_51_p VDD N_VDD_c_40_p
+ PM_SKY130_OSU_SC_18T_LS__OAI21_L%VDD
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%A0 N_A0_c_64_n N_A0_M1005_g N_A0_M1004_g
+ N_A0_c_68_n N_A0_c_69_n N_A0_c_70_n N_A0_c_71_n A0
+ PM_SKY130_OSU_SC_18T_LS__OAI21_L%A0
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%A1 N_A1_M1003_g N_A1_M1001_g N_A1_c_105_n
+ N_A1_c_106_n N_A1_c_107_n A1 PM_SKY130_OSU_SC_18T_LS__OAI21_L%A1
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%B0 N_B0_c_156_n N_B0_M1000_g N_B0_M1002_g
+ N_B0_c_160_n N_B0_c_161_n N_B0_c_162_n B0 PM_SKY130_OSU_SC_18T_LS__OAI21_L%B0
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%Y N_Y_M1002_d N_Y_M1004_s N_Y_M1000_d
+ N_Y_c_214_n N_Y_c_217_n N_Y_c_230_n N_Y_c_208_n N_Y_c_221_n N_Y_c_209_n
+ N_Y_c_224_n Y N_Y_c_212_n N_Y_c_213_n PM_SKY130_OSU_SC_18T_LS__OAI21_L%Y
x_PM_SKY130_OSU_SC_18T_LS__OAI21_L%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1001_d N_A_27_115#_c_267_n N_A_27_115#_c_270_n
+ N_A_27_115#_c_275_n N_A_27_115#_c_272_n
+ PM_SKY130_OSU_SC_18T_LS__OAI21_L%A_27_115#
cc_1 N_GND_M1005_b N_A0_c_64_n 0.0246907f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.7
cc_2 N_GND_c_2_p N_A0_c_64_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.7
cc_3 N_GND_c_3_p N_A0_c_64_n 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.7
cc_4 N_GND_c_4_p N_A0_c_64_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.7
cc_5 N_GND_M1005_b N_A0_c_68_n 0.0245405f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.775
cc_6 N_GND_M1005_b N_A0_c_69_n 0.0342885f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.76
cc_7 N_GND_M1005_b N_A0_c_70_n 0.0620905f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.595
cc_8 N_GND_M1005_b N_A0_c_71_n 0.0028102f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.76
cc_9 N_GND_M1005_b N_A1_M1003_g 0.0270518f $X=-0.045 $Y=0 $X2=0.835 $Y2=4.585
cc_10 N_GND_M1005_b N_A1_M1001_g 0.0452495f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.075
cc_11 N_GND_c_3_p N_A1_M1001_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905 $Y2=1.075
cc_12 N_GND_c_4_p N_A1_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=1.075
cc_13 N_GND_M1005_b N_A1_c_105_n 0.0317916f $X=-0.045 $Y=0 $X2=0.845 $Y2=2.22
cc_14 N_GND_M1005_b N_A1_c_106_n 0.00507239f $X=-0.045 $Y=0 $X2=0.845 $Y2=2.22
cc_15 N_GND_M1005_b N_A1_c_107_n 8.57225e-19 $X=-0.045 $Y=0 $X2=0.895 $Y2=2.96
cc_16 N_GND_M1005_b A1 0.00292188f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.96
cc_17 N_GND_M1005_b N_B0_c_156_n 0.0335277f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.045
cc_18 N_GND_M1005_b N_B0_M1000_g 0.0488857f $X=-0.045 $Y=0 $X2=1.325 $Y2=5.085
cc_19 N_GND_M1005_b N_B0_M1002_g 0.0300879f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.075
cc_20 N_GND_c_4_p N_B0_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335 $Y2=1.075
cc_21 N_GND_M1005_b N_B0_c_160_n 0.00586489f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.59
cc_22 N_GND_M1005_b N_B0_c_161_n 0.00505195f $X=-0.045 $Y=0 $X2=1.285 $Y2=1.88
cc_23 N_GND_M1005_b N_B0_c_162_n 0.00240282f $X=-0.045 $Y=0 $X2=1.395 $Y2=1.88
cc_24 N_GND_M1005_b B0 0.0119375f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.59
cc_25 N_GND_M1005_b N_Y_c_208_n 0.0317947f $X=-0.045 $Y=0 $X2=1.54 $Y2=2.22
cc_26 N_GND_M1005_b N_Y_c_209_n 0.00913846f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.82
cc_27 N_GND_c_4_p N_Y_c_209_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.82
cc_28 N_GND_M1005_b Y 0.0139051f $X=-0.045 $Y=0 $X2=1.54 $Y2=2.22
cc_29 N_GND_M1005_b N_Y_c_212_n 0.0205847f $X=-0.045 $Y=0 $X2=1.54 $Y2=2.105
cc_30 N_GND_M1005_b N_Y_c_213_n 0.0105874f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.48
cc_31 N_GND_M1005_b N_A_27_115#_c_267_n 0.00156053f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_32 N_GND_c_2_p N_A_27_115#_c_267_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_33 N_GND_c_4_p N_A_27_115#_c_267_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_34 N_GND_M1005_d N_A_27_115#_c_270_n 0.00645469f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.42
cc_35 N_GND_c_3_p N_A_27_115#_c_270_n 0.00986105f $X=0.69 $Y=0.825 $X2=1.035
+ $Y2=1.42
cc_36 N_GND_M1005_b N_A_27_115#_c_272_n 0.00889125f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.825
cc_37 N_GND_c_4_p N_A_27_115#_c_272_n 0.00475776f $X=1.02 $Y=0.19 $X2=1.12
+ $Y2=0.825
cc_38 N_VDD_M1004_b N_A0_M1004_g 0.0238089f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_39 N_VDD_c_39_p N_A0_M1004_g 0.00606474f $X=0.965 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_40 N_VDD_c_40_p N_A0_M1004_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=4.585
cc_41 N_VDD_M1004_b N_A0_c_69_n 0.00574563f $X=-0.045 $Y=2.905 $X2=0.415
+ $Y2=2.76
cc_42 N_VDD_M1004_b N_A0_c_71_n 0.00549657f $X=-0.045 $Y=2.905 $X2=0.415
+ $Y2=2.76
cc_43 N_VDD_M1004_b N_A1_M1003_g 0.0185298f $X=-0.045 $Y=2.905 $X2=0.835
+ $Y2=4.585
cc_44 N_VDD_c_39_p N_A1_M1003_g 0.00606474f $X=0.965 $Y=6.507 $X2=0.835
+ $Y2=4.585
cc_45 N_VDD_c_45_p N_A1_M1003_g 0.00373151f $X=1.05 $Y=4.475 $X2=0.835 $Y2=4.585
cc_46 N_VDD_c_40_p N_A1_M1003_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.835 $Y2=4.585
cc_47 N_VDD_M1004_b N_A1_c_107_n 0.00163533f $X=-0.045 $Y=2.905 $X2=0.895
+ $Y2=2.96
cc_48 N_VDD_M1004_b A1 0.00594612f $X=-0.045 $Y=2.905 $X2=0.895 $Y2=2.96
cc_49 N_VDD_M1004_b N_B0_M1000_g 0.0840802f $X=-0.045 $Y=2.905 $X2=1.325
+ $Y2=5.085
cc_50 N_VDD_c_45_p N_B0_M1000_g 0.0192185f $X=1.05 $Y=4.475 $X2=1.325 $Y2=5.085
cc_51 N_VDD_c_51_p N_B0_M1000_g 0.00606474f $X=1.02 $Y=6.47 $X2=1.325 $Y2=5.085
cc_52 N_VDD_c_40_p N_B0_M1000_g 0.00468827f $X=1.02 $Y=6.47 $X2=1.325 $Y2=5.085
cc_53 N_VDD_M1004_b N_Y_c_214_n 0.00156053f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.135
cc_54 N_VDD_c_39_p N_Y_c_214_n 0.00736239f $X=0.965 $Y=6.507 $X2=0.26 $Y2=4.135
cc_55 N_VDD_c_40_p N_Y_c_214_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26 $Y2=4.135
cc_56 N_VDD_M1003_d N_Y_c_217_n 0.00888984f $X=0.91 $Y=3.085 $X2=1.455 $Y2=3.67
cc_57 N_VDD_M1004_b N_Y_c_217_n 0.00886322f $X=-0.045 $Y=2.905 $X2=1.455
+ $Y2=3.67
cc_58 N_VDD_c_45_p N_Y_c_217_n 0.00639099f $X=1.05 $Y=4.475 $X2=1.455 $Y2=3.67
cc_59 N_VDD_M1004_b N_Y_c_208_n 0.032421f $X=-0.045 $Y=2.905 $X2=1.54 $Y2=2.22
cc_60 N_VDD_M1004_b N_Y_c_221_n 0.0170696f $X=-0.045 $Y=2.905 $X2=1.54 $Y2=4.475
cc_61 N_VDD_c_51_p N_Y_c_221_n 0.00757793f $X=1.02 $Y=6.47 $X2=1.54 $Y2=4.475
cc_62 N_VDD_c_40_p N_Y_c_221_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.54 $Y2=4.475
cc_63 N_VDD_M1004_b N_Y_c_224_n 0.00720662f $X=-0.045 $Y=2.905 $X2=1.54 $Y2=3.67
cc_64 N_A0_c_69_n N_A1_M1003_g 0.21737f $X=0.415 $Y=2.76 $X2=0.835 $Y2=4.585
cc_65 N_A0_c_70_n N_A1_M1003_g 0.00894734f $X=0.415 $Y=2.595 $X2=0.835 $Y2=4.585
cc_66 N_A0_c_71_n N_A1_M1003_g 0.00413298f $X=0.415 $Y=2.76 $X2=0.835 $Y2=4.585
cc_67 A0 N_A1_M1003_g 0.00376364f $X=0.415 $Y=3.33 $X2=0.835 $Y2=4.585
cc_68 N_A0_c_64_n N_A1_M1001_g 0.0445799f $X=0.475 $Y=1.7 $X2=0.905 $Y2=1.075
cc_69 N_A0_c_70_n N_A1_M1001_g 0.00745632f $X=0.415 $Y=2.595 $X2=0.905 $Y2=1.075
cc_70 N_A0_c_70_n N_A1_c_105_n 0.014675f $X=0.415 $Y=2.595 $X2=0.845 $Y2=2.22
cc_71 N_A0_c_69_n N_A1_c_106_n 8.44103e-19 $X=0.415 $Y=2.76 $X2=0.845 $Y2=2.22
cc_72 N_A0_c_70_n N_A1_c_106_n 0.00346793f $X=0.415 $Y=2.595 $X2=0.845 $Y2=2.22
cc_73 N_A0_c_71_n N_A1_c_106_n 0.0189532f $X=0.415 $Y=2.76 $X2=0.845 $Y2=2.22
cc_74 N_A0_M1004_g N_A1_c_107_n 8.44103e-19 $X=0.475 $Y=4.585 $X2=0.895 $Y2=2.96
cc_75 N_A0_c_69_n A1 0.00357623f $X=0.415 $Y=2.76 $X2=0.895 $Y2=2.96
cc_76 N_A0_c_71_n A1 0.00685942f $X=0.415 $Y=2.76 $X2=0.895 $Y2=2.96
cc_77 N_A0_c_71_n N_Y_M1004_s 0.00842425f $X=0.415 $Y=2.76 $X2=0.135 $Y2=3.085
cc_78 A0 N_Y_M1004_s 0.0119025f $X=0.415 $Y=3.33 $X2=0.135 $Y2=3.085
cc_79 N_A0_M1004_g N_Y_c_217_n 0.0157489f $X=0.475 $Y=4.585 $X2=1.455 $Y2=3.67
cc_80 N_A0_c_71_n N_Y_c_217_n 0.0069936f $X=0.415 $Y=2.76 $X2=1.455 $Y2=3.67
cc_81 A0 N_Y_c_217_n 0.0116431f $X=0.415 $Y=3.33 $X2=1.455 $Y2=3.67
cc_82 N_A0_c_69_n N_Y_c_230_n 0.00152768f $X=0.415 $Y=2.76 $X2=0.345 $Y2=3.67
cc_83 N_A0_c_71_n N_Y_c_230_n 9.01113e-19 $X=0.415 $Y=2.76 $X2=0.345 $Y2=3.67
cc_84 A0 N_Y_c_230_n 0.00385855f $X=0.415 $Y=3.33 $X2=0.345 $Y2=3.67
cc_85 A0 A_110_617# 0.0100173f $X=0.415 $Y=3.33 $X2=0.55 $Y2=3.085
cc_86 N_A0_c_64_n N_A_27_115#_c_270_n 0.0198204f $X=0.475 $Y=1.7 $X2=1.035
+ $Y2=1.42
cc_87 N_A0_c_68_n N_A_27_115#_c_275_n 0.0030143f $X=0.475 $Y=1.775 $X2=0.345
+ $Y2=1.42
cc_88 N_A1_M1001_g N_B0_c_156_n 0.00505587f $X=0.905 $Y=1.075 $X2=1.325
+ $Y2=2.045
cc_89 N_A1_M1003_g N_B0_M1000_g 0.0969479f $X=0.835 $Y=4.585 $X2=1.325 $Y2=5.085
cc_90 N_A1_c_105_n N_B0_M1000_g 0.014032f $X=0.845 $Y=2.22 $X2=1.325 $Y2=5.085
cc_91 N_A1_c_106_n N_B0_M1000_g 0.00248808f $X=0.845 $Y=2.22 $X2=1.325 $Y2=5.085
cc_92 N_A1_c_107_n N_B0_M1000_g 0.00113925f $X=0.895 $Y=2.96 $X2=1.325 $Y2=5.085
cc_93 A1 N_B0_M1000_g 0.00395308f $X=0.895 $Y=2.96 $X2=1.325 $Y2=5.085
cc_94 N_A1_M1001_g N_B0_M1002_g 0.0348492f $X=0.905 $Y=1.075 $X2=1.335 $Y2=1.075
cc_95 N_A1_M1003_g N_B0_c_160_n 9.28322e-19 $X=0.835 $Y=4.585 $X2=1.2 $Y2=2.59
cc_96 N_A1_M1001_g N_B0_c_160_n 0.00209141f $X=0.905 $Y=1.075 $X2=1.2 $Y2=2.59
cc_97 N_A1_c_105_n N_B0_c_160_n 0.00180004f $X=0.845 $Y=2.22 $X2=1.2 $Y2=2.59
cc_98 N_A1_c_106_n N_B0_c_160_n 0.0395776f $X=0.845 $Y=2.22 $X2=1.2 $Y2=2.59
cc_99 A1 N_B0_c_160_n 2.28089e-19 $X=0.895 $Y=2.96 $X2=1.2 $Y2=2.59
cc_100 N_A1_M1001_g N_B0_c_161_n 0.00444244f $X=0.905 $Y=1.075 $X2=1.285
+ $Y2=1.88
cc_101 N_A1_c_105_n B0 0.00173697f $X=0.845 $Y=2.22 $X2=1.2 $Y2=2.59
cc_102 N_A1_c_106_n B0 0.00816163f $X=0.845 $Y=2.22 $X2=1.2 $Y2=2.59
cc_103 N_A1_c_107_n B0 2.4196e-19 $X=0.895 $Y=2.96 $X2=1.2 $Y2=2.59
cc_104 A1 B0 0.0191116f $X=0.895 $Y=2.96 $X2=1.2 $Y2=2.59
cc_105 N_A1_M1003_g N_Y_c_217_n 0.0165071f $X=0.835 $Y=4.585 $X2=1.455 $Y2=3.67
cc_106 N_A1_c_107_n N_Y_c_217_n 0.00294448f $X=0.895 $Y=2.96 $X2=1.455 $Y2=3.67
cc_107 A1 N_Y_c_217_n 0.0102328f $X=0.895 $Y=2.96 $X2=1.455 $Y2=3.67
cc_108 N_A1_c_106_n N_Y_c_208_n 0.00577978f $X=0.845 $Y=2.22 $X2=1.54 $Y2=2.22
cc_109 N_A1_c_107_n N_Y_c_208_n 0.00365175f $X=0.895 $Y=2.96 $X2=1.54 $Y2=2.22
cc_110 A1 N_Y_c_208_n 0.00695805f $X=0.895 $Y=2.96 $X2=1.54 $Y2=2.22
cc_111 N_A1_M1001_g N_Y_c_212_n 3.31726e-19 $X=0.905 $Y=1.075 $X2=1.54 $Y2=2.105
cc_112 N_A1_M1001_g N_Y_c_213_n 4.01461e-19 $X=0.905 $Y=1.075 $X2=1.55 $Y2=1.48
cc_113 N_A1_M1001_g N_A_27_115#_c_270_n 0.0170616f $X=0.905 $Y=1.075 $X2=1.035
+ $Y2=1.42
cc_114 N_A1_c_105_n N_A_27_115#_c_270_n 0.00211261f $X=0.845 $Y=2.22 $X2=1.035
+ $Y2=1.42
cc_115 N_A1_c_106_n N_A_27_115#_c_270_n 0.00447151f $X=0.845 $Y=2.22 $X2=1.035
+ $Y2=1.42
cc_116 N_B0_M1000_g N_Y_c_217_n 0.0210988f $X=1.325 $Y=5.085 $X2=1.455 $Y2=3.67
cc_117 N_B0_c_156_n N_Y_c_208_n 0.00149952f $X=1.325 $Y=2.045 $X2=1.54 $Y2=2.22
cc_118 N_B0_M1000_g N_Y_c_208_n 0.0418701f $X=1.325 $Y=5.085 $X2=1.54 $Y2=2.22
cc_119 N_B0_c_160_n N_Y_c_208_n 0.0348659f $X=1.2 $Y=2.59 $X2=1.54 $Y2=2.22
cc_120 N_B0_c_162_n N_Y_c_208_n 0.00728781f $X=1.395 $Y=1.88 $X2=1.54 $Y2=2.22
cc_121 B0 N_Y_c_208_n 0.00659213f $X=1.2 $Y=2.59 $X2=1.54 $Y2=2.22
cc_122 N_B0_M1000_g N_Y_c_221_n 0.0175573f $X=1.325 $Y=5.085 $X2=1.54 $Y2=4.475
cc_123 N_B0_c_156_n N_Y_c_209_n 0.00116804f $X=1.325 $Y=2.045 $X2=1.55 $Y2=0.82
cc_124 N_B0_M1002_g N_Y_c_209_n 0.00518773f $X=1.335 $Y=1.075 $X2=1.55 $Y2=0.82
cc_125 N_B0_c_162_n N_Y_c_209_n 0.00472322f $X=1.395 $Y=1.88 $X2=1.55 $Y2=0.82
cc_126 N_B0_c_156_n Y 0.00133576f $X=1.325 $Y=2.045 $X2=1.54 $Y2=2.22
cc_127 N_B0_M1000_g Y 0.00488821f $X=1.325 $Y=5.085 $X2=1.54 $Y2=2.22
cc_128 N_B0_c_160_n Y 0.00656407f $X=1.2 $Y=2.59 $X2=1.54 $Y2=2.22
cc_129 N_B0_c_162_n Y 0.00199558f $X=1.395 $Y=1.88 $X2=1.54 $Y2=2.22
cc_130 N_B0_c_156_n N_Y_c_212_n 0.00526688f $X=1.325 $Y=2.045 $X2=1.54 $Y2=2.105
cc_131 N_B0_M1000_g N_Y_c_212_n 0.00137073f $X=1.325 $Y=5.085 $X2=1.54 $Y2=2.105
cc_132 N_B0_M1002_g N_Y_c_212_n 0.00278116f $X=1.335 $Y=1.075 $X2=1.54 $Y2=2.105
cc_133 N_B0_c_160_n N_Y_c_212_n 0.00553065f $X=1.2 $Y=2.59 $X2=1.54 $Y2=2.105
cc_134 N_B0_c_162_n N_Y_c_212_n 0.0118918f $X=1.395 $Y=1.88 $X2=1.54 $Y2=2.105
cc_135 N_B0_c_156_n N_Y_c_213_n 0.00101197f $X=1.325 $Y=2.045 $X2=1.55 $Y2=1.48
cc_136 N_B0_M1002_g N_Y_c_213_n 0.00586282f $X=1.335 $Y=1.075 $X2=1.55 $Y2=1.48
cc_137 N_B0_c_162_n N_Y_c_213_n 0.00157776f $X=1.395 $Y=1.88 $X2=1.55 $Y2=1.48
cc_138 N_B0_c_161_n N_A_27_115#_c_270_n 0.00556868f $X=1.285 $Y=1.88 $X2=1.035
+ $Y2=1.42
cc_139 N_Y_c_217_n A_110_617# 0.00573878f $X=1.455 $Y=3.67 $X2=0.55 $Y2=3.085
cc_140 N_Y_c_213_n N_A_27_115#_c_270_n 0.00369865f $X=1.55 $Y=1.48 $X2=1.035
+ $Y2=1.42
