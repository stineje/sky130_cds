* File: sky130_osu_sc_18T_ls__pcgate_1.pxi.spice
* Created: Thu Mar 10 13:46:56 2022
* 
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%GND N_GND_M1010_s N_GND_M1018_d
+ N_GND_M1024_d N_GND_M1001_d N_GND_M1017_d N_GND_M1012_d N_GND_M1010_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_14_p N_GND_c_22_p N_GND_c_19_p N_GND_c_33_p
+ N_GND_c_56_p N_GND_c_57_p N_GND_c_112_p N_GND_c_61_p N_GND_c_62_p GND GND GND
+ GND GND GND GND GND GND GND PM_SKY130_OSU_SC_18T_LS__PCGATE_1%GND
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%VDD N_VDD_M1007_d N_VDD_M1022_d
+ N_VDD_M1014_d N_VDD_M1020_d N_VDD_M1021_s N_VDD_M1005_d N_VDD_M1025_b
+ N_VDD_c_182_p N_VDD_c_188_p N_VDD_c_198_p N_VDD_c_199_p N_VDD_c_205_p
+ N_VDD_c_218_p N_VDD_c_219_p N_VDD_c_230_p N_VDD_c_259_p N_VDD_c_260_p
+ N_VDD_c_222_p N_VDD_c_223_p N_VDD_c_284_p VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD PM_SKY130_OSU_SC_18T_LS__PCGATE_1%VDD
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%SE N_SE_M1010_g N_SE_M1025_g N_SE_c_305_n
+ N_SE_c_307_n N_SE_c_309_n SE N_SE_X27_noxref_CONDUCTOR
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%SE
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%E N_E_M1007_g N_E_M1018_g N_E_c_355_n
+ N_E_c_356_n E PM_SKY130_OSU_SC_18T_LS__PCGATE_1%E
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_86_337# N_A_86_337#_M1019_d
+ N_A_86_337#_M1004_d N_A_86_337#_M1024_g N_A_86_337#_M1022_g
+ N_A_86_337#_c_398_n N_A_86_337#_c_400_n N_A_86_337#_c_405_n
+ N_A_86_337#_c_406_n N_A_86_337#_c_407_n N_A_86_337#_c_408_n
+ N_A_86_337#_c_409_n N_A_86_337#_c_421_n N_A_86_337#_c_472_p
+ N_A_86_337#_c_411_n N_A_86_337#_c_454_p N_A_86_337#_c_434_p
+ N_A_86_337#_c_412_n N_A_86_337#_c_423_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_86_337#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_N233_617# N_A_N233_617#_M1010_d
+ N_A_N233_617#_M1025_s N_A_N233_617#_M1023_g N_A_N233_617#_M1002_g
+ N_A_N233_617#_c_489_n N_A_N233_617#_c_490_n N_A_N233_617#_c_491_n
+ N_A_N233_617#_c_494_n N_A_N233_617#_c_495_n N_A_N233_617#_c_496_n
+ N_A_N233_617#_c_497_n N_A_N233_617#_c_498_n N_A_N233_617#_c_501_n
+ N_A_N233_617#_c_502_n N_A_N233_617#_c_503_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_N233_617#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%CK N_CK_M1004_g N_CK_M1011_g N_CK_c_595_n
+ N_CK_M1003_g N_CK_M1000_g N_CK_c_599_n N_CK_M1012_g N_CK_M1005_g N_CK_c_605_n
+ N_CK_c_606_n N_CK_c_607_n N_CK_c_610_n N_CK_c_611_n N_CK_c_612_n N_CK_c_613_n
+ N_CK_c_614_n N_CK_c_616_n N_CK_c_617_n N_CK_c_618_n N_CK_c_619_n N_CK_c_620_n
+ N_CK_c_621_n CK N_CK_c_623_n PM_SKY130_OSU_SC_18T_LS__PCGATE_1%CK
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_254_89# N_A_254_89#_M1003_d
+ N_A_254_89#_M1000_d N_A_254_89#_M1019_g N_A_254_89#_c_792_n
+ N_A_254_89#_c_793_n N_A_254_89#_M1013_g N_A_254_89#_c_794_n
+ N_A_254_89#_c_795_n N_A_254_89#_c_796_n N_A_254_89#_c_797_n
+ N_A_254_89#_c_800_n N_A_254_89#_c_801_n N_A_254_89#_c_802_n
+ N_A_254_89#_c_803_n N_A_254_89#_c_804_n N_A_254_89#_c_805_n
+ N_A_254_89#_c_806_n PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_254_89#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_43_115# N_A_43_115#_M1024_s
+ N_A_43_115#_M1022_s N_A_43_115#_M1001_g N_A_43_115#_M1014_g
+ N_A_43_115#_M1017_g N_A_43_115#_M1020_g N_A_43_115#_c_927_n
+ N_A_43_115#_c_928_n N_A_43_115#_c_929_n N_A_43_115#_c_930_n
+ N_A_43_115#_c_934_n N_A_43_115#_c_935_n N_A_43_115#_c_936_n
+ N_A_43_115#_c_937_n N_A_43_115#_c_938_n N_A_43_115#_c_960_n
+ N_A_43_115#_c_942_n N_A_43_115#_c_943_n N_A_43_115#_c_944_n
+ N_A_43_115#_c_964_n N_A_43_115#_c_946_n N_A_43_115#_c_947_n
+ N_A_43_115#_c_948_n N_A_43_115#_c_949_n N_A_43_115#_c_950_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_43_115#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_687_115# N_A_687_115#_M1017_s
+ N_A_687_115#_M1020_s N_A_687_115#_M1006_g N_A_687_115#_M1009_g
+ N_A_687_115#_M1015_g N_A_687_115#_M1021_g N_A_687_115#_c_1111_n
+ N_A_687_115#_c_1112_n N_A_687_115#_c_1113_n N_A_687_115#_c_1116_n
+ N_A_687_115#_c_1117_n N_A_687_115#_c_1119_n N_A_687_115#_c_1120_n
+ N_A_687_115#_c_1121_n N_A_687_115#_c_1122_n N_A_687_115#_c_1123_n
+ N_A_687_115#_c_1142_n N_A_687_115#_c_1147_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_687_115#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_963_115# N_A_963_115#_M1015_s
+ N_A_963_115#_M1021_d N_A_963_115#_M1008_g N_A_963_115#_M1016_g
+ N_A_963_115#_c_1234_n N_A_963_115#_c_1235_n N_A_963_115#_c_1236_n
+ N_A_963_115#_c_1237_n N_A_963_115#_c_1240_n N_A_963_115#_c_1241_n
+ N_A_963_115#_c_1251_n N_A_963_115#_c_1242_n N_A_963_115#_c_1244_n
+ N_A_963_115#_c_1245_n N_A_963_115#_c_1271_n N_A_963_115#_c_1246_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_963_115#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_856_115# N_A_856_115#_M1006_d
+ N_A_856_115#_M1009_d N_A_856_115#_c_1309_n N_A_856_115#_c_1314_n
+ N_A_856_115#_c_1312_n N_A_856_115#_c_1313_n N_A_856_115#_c_1319_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_856_115#
x_PM_SKY130_OSU_SC_18T_LS__PCGATE_1%ECK N_ECK_M1008_d N_ECK_M1016_d
+ N_ECK_c_1343_n N_ECK_c_1346_n ECK N_ECK_c_1348_n N_ECK_c_1350_n
+ PM_SKY130_OSU_SC_18T_LS__PCGATE_1%ECK
cc_1 N_GND_M1010_b N_SE_M1010_g 0.0397546f $X=-1.345 $Y=0 $X2=-0.825 $Y2=1.075
cc_2 N_GND_c_2_p N_SE_M1010_g 0.00713292f $X=-1.039 $Y=0.825 $X2=-0.825
+ $Y2=1.075
cc_3 N_GND_c_3_p N_SE_M1010_g 0.00606474f $X=-0.265 $Y=0.152 $X2=-0.825
+ $Y2=1.075
cc_4 GND N_SE_M1010_g 0.00468827f $X=5.7 $Y=0.2 $X2=-0.825 $Y2=1.075
cc_5 N_GND_M1010_b N_SE_M1025_g 0.0432223f $X=-1.345 $Y=0 $X2=-0.825 $Y2=4.585
cc_6 N_GND_M1010_b N_SE_c_305_n 0.0362021f $X=-1.345 $Y=0 $X2=-0.884 $Y2=2.09
cc_7 N_GND_c_2_p N_SE_c_305_n 0.00122211f $X=-1.039 $Y=0.825 $X2=-0.884 $Y2=2.09
cc_8 N_GND_M1010_b N_SE_c_307_n 0.0115466f $X=-1.345 $Y=0 $X2=-0.735 $Y2=2.09
cc_9 N_GND_c_2_p N_SE_c_307_n 0.00289632f $X=-1.039 $Y=0.825 $X2=-0.735 $Y2=2.09
cc_10 N_GND_M1010_b N_SE_c_309_n 0.0148494f $X=-1.345 $Y=0 $X2=-0.649 $Y2=2.96
cc_11 N_GND_M1010_b N_SE_X27_noxref_CONDUCTOR 5.7362e-19 $X=-1.345 $Y=0
+ $X2=-0.654 $Y2=2.96
cc_12 N_GND_M1010_b N_E_M1018_g 0.0744003f $X=-1.345 $Y=0 $X2=-0.395 $Y2=1.075
cc_13 N_GND_c_3_p N_E_M1018_g 0.00606474f $X=-0.265 $Y=0.152 $X2=-0.395
+ $Y2=1.075
cc_14 N_GND_c_14_p N_E_M1018_g 0.00713292f $X=-0.179 $Y=0.825 $X2=-0.395
+ $Y2=1.075
cc_15 GND N_E_M1018_g 0.00468827f $X=5.7 $Y=0.2 $X2=-0.395 $Y2=1.075
cc_16 N_GND_M1010_b N_E_c_355_n 0.0320151f $X=-1.345 $Y=0 $X2=-0.309 $Y2=2.755
cc_17 N_GND_M1010_b N_E_c_356_n 0.00121702f $X=-1.345 $Y=0 $X2=-0.309 $Y2=2.755
cc_18 N_GND_M1010_b N_A_86_337#_c_398_n 0.030793f $X=-1.345 $Y=0 $X2=0.565
+ $Y2=1.85
cc_19 N_GND_c_19_p N_A_86_337#_c_398_n 3.17551e-19 $X=0.77 $Y=0.825 $X2=0.565
+ $Y2=1.85
cc_20 N_GND_M1010_b N_A_86_337#_c_400_n 0.0184872f $X=-1.345 $Y=0 $X2=0.565
+ $Y2=1.685
cc_21 N_GND_c_14_p N_A_86_337#_c_400_n 0.00458302f $X=-0.179 $Y=0.825 $X2=0.565
+ $Y2=1.685
cc_22 N_GND_c_22_p N_A_86_337#_c_400_n 0.00606474f $X=0.685 $Y=0.152 $X2=0.565
+ $Y2=1.685
cc_23 N_GND_c_19_p N_A_86_337#_c_400_n 0.00354579f $X=0.77 $Y=0.825 $X2=0.565
+ $Y2=1.685
cc_24 GND N_A_86_337#_c_400_n 0.00468827f $X=5.7 $Y=0.2 $X2=0.565 $Y2=1.685
cc_25 N_GND_M1010_b N_A_86_337#_c_405_n 0.0436413f $X=-1.345 $Y=0 $X2=0.53
+ $Y2=2.805
cc_26 N_GND_M1010_b N_A_86_337#_c_406_n 0.00768983f $X=-1.345 $Y=0 $X2=0.53
+ $Y2=2.975
cc_27 N_GND_M1010_b N_A_86_337#_c_407_n 8.14549e-19 $X=-1.345 $Y=0 $X2=0.565
+ $Y2=1.935
cc_28 N_GND_M1010_b N_A_86_337#_c_408_n 0.00684609f $X=-1.345 $Y=0 $X2=0.565
+ $Y2=3.1
cc_29 N_GND_M1010_b N_A_86_337#_c_409_n 0.00828074f $X=-1.345 $Y=0 $X2=1.025
+ $Y2=1.85
cc_30 N_GND_c_19_p N_A_86_337#_c_409_n 0.00816426f $X=0.77 $Y=0.825 $X2=1.025
+ $Y2=1.85
cc_31 N_GND_M1010_b N_A_86_337#_c_411_n 0.00172671f $X=-1.345 $Y=0 $X2=1.11
+ $Y2=1.765
cc_32 N_GND_M1010_b N_A_86_337#_c_412_n 0.00313975f $X=-1.345 $Y=0 $X2=1.645
+ $Y2=0.825
cc_33 N_GND_c_33_p N_A_86_337#_c_412_n 0.0151591f $X=2.435 $Y=0.152 $X2=1.645
+ $Y2=0.825
cc_34 GND N_A_86_337#_c_412_n 0.00958198f $X=5.7 $Y=0.2 $X2=1.645 $Y2=0.825
cc_35 N_GND_M1010_b N_A_N233_617#_M1023_g 0.040459f $X=-1.345 $Y=0 $X2=0.985
+ $Y2=1.075
cc_36 N_GND_c_19_p N_A_N233_617#_M1023_g 0.00354579f $X=0.77 $Y=0.825 $X2=0.985
+ $Y2=1.075
cc_37 N_GND_c_33_p N_A_N233_617#_M1023_g 0.00606474f $X=2.435 $Y=0.152 $X2=0.985
+ $Y2=1.075
cc_38 GND N_A_N233_617#_M1023_g 0.00468827f $X=5.7 $Y=0.2 $X2=0.985 $Y2=1.075
cc_39 N_GND_M1010_b N_A_N233_617#_M1002_g 0.0152797f $X=-1.345 $Y=0 $X2=0.985
+ $Y2=4.585
cc_40 N_GND_M1010_b N_A_N233_617#_c_489_n 0.0294636f $X=-1.345 $Y=0 $X2=0.925
+ $Y2=2.425
cc_41 N_GND_M1010_b N_A_N233_617#_c_490_n 0.0154673f $X=-1.345 $Y=0 $X2=-1.039
+ $Y2=2.59
cc_42 N_GND_M1010_b N_A_N233_617#_c_491_n 0.00155118f $X=-1.345 $Y=0 $X2=-0.609
+ $Y2=0.825
cc_43 N_GND_c_3_p N_A_N233_617#_c_491_n 0.0075556f $X=-0.265 $Y=0.152 $X2=-0.609
+ $Y2=0.825
cc_44 GND N_A_N233_617#_c_491_n 0.00475776f $X=5.7 $Y=0.2 $X2=-0.609 $Y2=0.825
cc_45 N_GND_M1010_b N_A_N233_617#_c_494_n 0.00123417f $X=-1.345 $Y=0 $X2=0.925
+ $Y2=2.425
cc_46 N_GND_M1010_b N_A_N233_617#_c_495_n 2.54997e-19 $X=-1.345 $Y=0 $X2=-0.71
+ $Y2=2.59
cc_47 N_GND_M1010_b N_A_N233_617#_c_496_n 0.019675f $X=-1.345 $Y=0 $X2=-0.895
+ $Y2=2.59
cc_48 N_GND_M1010_b N_A_N233_617#_c_497_n 0.0195542f $X=-1.345 $Y=0 $X2=-0.61
+ $Y2=2.505
cc_49 N_GND_M1010_b N_A_N233_617#_c_498_n 0.00257875f $X=-1.345 $Y=0 $X2=-0.609
+ $Y2=1.48
cc_50 N_GND_c_2_p N_A_N233_617#_c_498_n 0.00125659f $X=-1.039 $Y=0.825
+ $X2=-0.609 $Y2=1.48
cc_51 N_GND_c_14_p N_A_N233_617#_c_498_n 0.00125659f $X=-0.179 $Y=0.825
+ $X2=-0.609 $Y2=1.48
cc_52 N_GND_M1010_b N_A_N233_617#_c_501_n 2.05597e-19 $X=-1.345 $Y=0 $X2=-0.617
+ $Y2=2.592
cc_53 N_GND_M1010_b N_A_N233_617#_c_502_n 0.00372686f $X=-1.345 $Y=0 $X2=0.925
+ $Y2=2.595
cc_54 N_GND_M1010_b N_A_N233_617#_c_503_n 0.0361375f $X=-1.345 $Y=0 $X2=0.78
+ $Y2=2.595
cc_55 N_GND_M1010_b N_CK_c_595_n 0.0198314f $X=-1.345 $Y=0 $X2=2.735 $Y2=1.665
cc_56 N_GND_c_56_p N_CK_c_595_n 0.00354579f $X=2.52 $Y=0.825 $X2=2.735 $Y2=1.665
cc_57 N_GND_c_57_p N_CK_c_595_n 0.00606474f $X=3.905 $Y=0.152 $X2=2.735
+ $Y2=1.665
cc_58 GND N_CK_c_595_n 0.00468827f $X=5.7 $Y=0.2 $X2=2.735 $Y2=1.665
cc_59 N_GND_M1010_b N_CK_c_599_n 0.0384772f $X=-1.345 $Y=0 $X2=2.79 $Y2=2.015
cc_60 N_GND_M1010_b N_CK_M1012_g 0.0460454f $X=-1.345 $Y=0 $X2=5.515 $Y2=1.075
cc_61 N_GND_c_61_p N_CK_M1012_g 0.00606474f $X=5.645 $Y=0.152 $X2=5.515
+ $Y2=1.075
cc_62 N_GND_c_62_p N_CK_M1012_g 0.00376152f $X=5.73 $Y=0.825 $X2=5.515 $Y2=1.075
cc_63 GND N_CK_M1012_g 0.00468827f $X=5.7 $Y=0.2 $X2=5.515 $Y2=1.075
cc_64 N_GND_M1010_b N_CK_M1005_g 0.0151186f $X=-1.345 $Y=0 $X2=5.585 $Y2=4.585
cc_65 N_GND_M1010_b N_CK_c_605_n 0.019325f $X=-1.345 $Y=0 $X2=1.405 $Y2=2.765
cc_66 N_GND_M1010_b N_CK_c_606_n 0.030276f $X=-1.345 $Y=0 $X2=1.885 $Y2=1.85
cc_67 N_GND_M1010_b N_CK_c_607_n 0.0175443f $X=-1.345 $Y=0 $X2=1.885 $Y2=1.685
cc_68 N_GND_c_33_p N_CK_c_607_n 0.00606474f $X=2.435 $Y=0.152 $X2=1.885
+ $Y2=1.685
cc_69 GND N_CK_c_607_n 0.00468827f $X=5.7 $Y=0.2 $X2=1.885 $Y2=1.685
cc_70 N_GND_M1010_b N_CK_c_610_n 0.0457025f $X=-1.345 $Y=0 $X2=2.762 $Y2=2.78
cc_71 N_GND_M1010_b N_CK_c_611_n 0.0101975f $X=-1.345 $Y=0 $X2=2.762 $Y2=2.935
cc_72 N_GND_M1010_b N_CK_c_612_n 0.0333619f $X=-1.345 $Y=0 $X2=5.63 $Y2=2.425
cc_73 N_GND_M1010_b N_CK_c_613_n 0.0071862f $X=-1.345 $Y=0 $X2=1.485 $Y2=2.68
cc_74 N_GND_M1010_b N_CK_c_614_n 0.0197856f $X=-1.345 $Y=0 $X2=2.785 $Y2=1.85
cc_75 N_GND_c_56_p N_CK_c_614_n 0.00821845f $X=2.52 $Y=0.825 $X2=2.785 $Y2=1.85
cc_76 N_GND_M1010_b N_CK_c_616_n 0.00162414f $X=-1.345 $Y=0 $X2=1.57 $Y2=1.85
cc_77 N_GND_M1010_b N_CK_c_617_n 0.00382966f $X=-1.345 $Y=0 $X2=5.63 $Y2=2.425
cc_78 N_GND_M1010_b N_CK_c_618_n 0.00355685f $X=-1.345 $Y=0 $X2=1.485 $Y2=2.765
cc_79 N_GND_M1010_b N_CK_c_619_n 6.52287e-19 $X=-1.345 $Y=0 $X2=2.87 $Y2=1.85
cc_80 N_GND_M1010_b N_CK_c_620_n 0.0335219f $X=-1.345 $Y=0 $X2=5.485 $Y2=2.96
cc_81 N_GND_M1010_b N_CK_c_621_n 9.0161e-19 $X=-1.345 $Y=0 $X2=1.405 $Y2=2.765
cc_82 N_GND_M1010_b CK 0.00516995f $X=-1.345 $Y=0 $X2=2.87 $Y2=1.85
cc_83 N_GND_M1010_b N_CK_c_623_n 0.00229761f $X=-1.345 $Y=0 $X2=5.63 $Y2=2.96
cc_84 N_GND_M1010_b N_A_254_89#_M1019_g 0.0458897f $X=-1.345 $Y=0 $X2=1.345
+ $Y2=1.075
cc_85 N_GND_c_33_p N_A_254_89#_M1019_g 0.00606474f $X=2.435 $Y=0.152 $X2=1.345
+ $Y2=1.075
cc_86 GND N_A_254_89#_M1019_g 0.00468827f $X=5.7 $Y=0.2 $X2=1.345 $Y2=1.075
cc_87 N_GND_M1010_b N_A_254_89#_c_792_n 0.030995f $X=-1.345 $Y=0 $X2=1.75
+ $Y2=2.3
cc_88 N_GND_M1010_b N_A_254_89#_c_793_n 0.00717301f $X=-1.345 $Y=0 $X2=1.42
+ $Y2=2.3
cc_89 N_GND_M1010_b N_A_254_89#_c_794_n 0.0199715f $X=-1.345 $Y=0 $X2=1.885
+ $Y2=2.765
cc_90 N_GND_M1010_b N_A_254_89#_c_795_n 0.0135787f $X=-1.345 $Y=0 $X2=1.885
+ $Y2=2.6
cc_91 N_GND_M1010_b N_A_254_89#_c_796_n 0.00180771f $X=-1.345 $Y=0 $X2=1.885
+ $Y2=2.59
cc_92 N_GND_M1010_b N_A_254_89#_c_797_n 0.00156053f $X=-1.345 $Y=0 $X2=2.95
+ $Y2=0.825
cc_93 N_GND_c_57_p N_A_254_89#_c_797_n 0.00754714f $X=3.905 $Y=0.152 $X2=2.95
+ $Y2=0.825
cc_94 GND N_A_254_89#_c_797_n 0.00476261f $X=5.7 $Y=0.2 $X2=2.95 $Y2=0.825
cc_95 N_GND_M1010_b N_A_254_89#_c_800_n 0.0161589f $X=-1.345 $Y=0 $X2=2.95
+ $Y2=2.59
cc_96 N_GND_M1010_b N_A_254_89#_c_801_n 0.0147893f $X=-1.345 $Y=0 $X2=3.22
+ $Y2=2.185
cc_97 N_GND_M1010_b N_A_254_89#_c_802_n 0.0118737f $X=-1.345 $Y=0 $X2=3.22
+ $Y2=1.43
cc_98 N_GND_M1010_b N_A_254_89#_c_803_n 0.00984894f $X=-1.345 $Y=0 $X2=3.22
+ $Y2=2.27
cc_99 N_GND_M1010_b N_A_254_89#_c_804_n 0.00651068f $X=-1.345 $Y=0 $X2=2.805
+ $Y2=2.59
cc_100 N_GND_M1010_b N_A_254_89#_c_805_n 0.00333963f $X=-1.345 $Y=0 $X2=2.03
+ $Y2=2.59
cc_101 N_GND_M1010_b N_A_254_89#_c_806_n 0.00457565f $X=-1.345 $Y=0 $X2=2.95
+ $Y2=2.59
cc_102 N_GND_M1010_b N_A_43_115#_M1001_g 0.0341452f $X=-1.345 $Y=0 $X2=2.305
+ $Y2=1.075
cc_103 N_GND_c_33_p N_A_43_115#_M1001_g 0.00606474f $X=2.435 $Y=0.152 $X2=2.305
+ $Y2=1.075
cc_104 N_GND_c_56_p N_A_43_115#_M1001_g 0.00354579f $X=2.52 $Y=0.825 $X2=2.305
+ $Y2=1.075
cc_105 GND N_A_43_115#_M1001_g 0.00468827f $X=5.7 $Y=0.2 $X2=2.305 $Y2=1.075
cc_106 N_GND_M1010_b N_A_43_115#_M1014_g 0.026298f $X=-1.345 $Y=0 $X2=2.305
+ $Y2=4.585
cc_107 N_GND_M1010_b N_A_43_115#_c_927_n 0.0287062f $X=-1.345 $Y=0 $X2=2.365
+ $Y2=2.22
cc_108 N_GND_M1010_b N_A_43_115#_c_928_n 0.0282666f $X=-1.345 $Y=0 $X2=3.66
+ $Y2=2.22
cc_109 N_GND_M1010_b N_A_43_115#_c_929_n 0.0149535f $X=-1.345 $Y=0 $X2=3.662
+ $Y2=2.055
cc_110 N_GND_M1010_b N_A_43_115#_c_930_n 0.0186694f $X=-1.345 $Y=0 $X2=3.75
+ $Y2=1.65
cc_111 N_GND_c_57_p N_A_43_115#_c_930_n 0.00606474f $X=3.905 $Y=0.152 $X2=3.75
+ $Y2=1.65
cc_112 N_GND_c_112_p N_A_43_115#_c_930_n 0.00354579f $X=3.99 $Y=0.825 $X2=3.75
+ $Y2=1.65
cc_113 GND N_A_43_115#_c_930_n 0.00468827f $X=5.7 $Y=0.2 $X2=3.75 $Y2=1.65
cc_114 N_GND_M1010_b N_A_43_115#_c_934_n 0.014038f $X=-1.345 $Y=0 $X2=3.75
+ $Y2=1.8
cc_115 N_GND_M1010_b N_A_43_115#_c_935_n 0.0300269f $X=-1.345 $Y=0 $X2=3.75
+ $Y2=2.855
cc_116 N_GND_M1010_b N_A_43_115#_c_936_n 0.00455351f $X=-1.345 $Y=0 $X2=3.75
+ $Y2=3.005
cc_117 N_GND_M1010_b N_A_43_115#_c_937_n 0.0315483f $X=-1.345 $Y=0 $X2=0.225
+ $Y2=2.22
cc_118 N_GND_M1010_b N_A_43_115#_c_938_n 0.00156053f $X=-1.345 $Y=0 $X2=0.34
+ $Y2=0.825
cc_119 N_GND_c_14_p N_A_43_115#_c_938_n 0.031398f $X=-0.179 $Y=0.825 $X2=0.34
+ $Y2=0.825
cc_120 N_GND_c_22_p N_A_43_115#_c_938_n 0.00757793f $X=0.685 $Y=0.152 $X2=0.34
+ $Y2=0.825
cc_121 GND N_A_43_115#_c_938_n 0.00476261f $X=5.7 $Y=0.2 $X2=0.34 $Y2=0.825
cc_122 N_GND_M1010_b N_A_43_115#_c_942_n 0.00378615f $X=-1.345 $Y=0 $X2=2.365
+ $Y2=2.22
cc_123 N_GND_M1010_b N_A_43_115#_c_943_n 0.00278582f $X=-1.345 $Y=0 $X2=3.66
+ $Y2=2.22
cc_124 N_GND_M1010_b N_A_43_115#_c_944_n 0.00474188f $X=-1.345 $Y=0 $X2=0.34
+ $Y2=1.395
cc_125 N_GND_c_14_p N_A_43_115#_c_944_n 0.00619665f $X=-0.179 $Y=0.825 $X2=0.34
+ $Y2=1.395
cc_126 N_GND_M1010_b N_A_43_115#_c_946_n 0.0198973f $X=-1.345 $Y=0 $X2=3.515
+ $Y2=2.22
cc_127 N_GND_M1010_b N_A_43_115#_c_947_n 0.00257231f $X=-1.345 $Y=0 $X2=2.515
+ $Y2=2.22
cc_128 N_GND_M1010_b N_A_43_115#_c_948_n 0.0101652f $X=-1.345 $Y=0 $X2=0.37
+ $Y2=2.22
cc_129 N_GND_M1010_b N_A_43_115#_c_949_n 0.0205759f $X=-1.345 $Y=0 $X2=2.22
+ $Y2=2.22
cc_130 N_GND_M1010_b N_A_43_115#_c_950_n 0.00118383f $X=-1.345 $Y=0 $X2=3.66
+ $Y2=2.22
cc_131 N_GND_M1010_b N_A_687_115#_M1006_g 0.0404979f $X=-1.345 $Y=0 $X2=4.205
+ $Y2=1.075
cc_132 N_GND_c_112_p N_A_687_115#_M1006_g 0.00354579f $X=3.99 $Y=0.825 $X2=4.205
+ $Y2=1.075
cc_133 N_GND_c_61_p N_A_687_115#_M1006_g 0.00606474f $X=5.645 $Y=0.152 $X2=4.205
+ $Y2=1.075
cc_134 GND N_A_687_115#_M1006_g 0.00468827f $X=5.7 $Y=0.2 $X2=4.205 $Y2=1.075
cc_135 N_GND_M1010_b N_A_687_115#_M1009_g 0.0285024f $X=-1.345 $Y=0 $X2=4.205
+ $Y2=4.585
cc_136 N_GND_M1010_b N_A_687_115#_M1015_g 0.0697889f $X=-1.345 $Y=0 $X2=5.155
+ $Y2=1.075
cc_137 N_GND_c_61_p N_A_687_115#_M1015_g 0.00606474f $X=5.645 $Y=0.152 $X2=5.155
+ $Y2=1.075
cc_138 GND N_A_687_115#_M1015_g 0.00468827f $X=5.7 $Y=0.2 $X2=5.155 $Y2=1.075
cc_139 N_GND_M1010_b N_A_687_115#_c_1111_n 0.0289774f $X=-1.345 $Y=0 $X2=4.145
+ $Y2=2.22
cc_140 N_GND_M1010_b N_A_687_115#_c_1112_n 0.0338801f $X=-1.345 $Y=0 $X2=5.155
+ $Y2=2.765
cc_141 N_GND_M1010_b N_A_687_115#_c_1113_n 0.00470373f $X=-1.345 $Y=0 $X2=3.56
+ $Y2=0.825
cc_142 N_GND_c_57_p N_A_687_115#_c_1113_n 0.00745733f $X=3.905 $Y=0.152 $X2=3.56
+ $Y2=0.825
cc_143 GND N_A_687_115#_c_1113_n 0.00476261f $X=5.7 $Y=0.2 $X2=3.56 $Y2=0.825
cc_144 N_GND_M1010_b N_A_687_115#_c_1116_n 0.0010765f $X=-1.345 $Y=0 $X2=3.56
+ $Y2=3.33
cc_145 N_GND_M1010_b N_A_687_115#_c_1117_n 0.0132938f $X=-1.345 $Y=0 $X2=4.06
+ $Y2=1.85
cc_146 N_GND_c_112_p N_A_687_115#_c_1117_n 0.00827205f $X=3.99 $Y=0.825 $X2=4.06
+ $Y2=1.85
cc_147 N_GND_M1010_b N_A_687_115#_c_1119_n 0.0022559f $X=-1.345 $Y=0 $X2=3.645
+ $Y2=1.85
cc_148 N_GND_M1010_b N_A_687_115#_c_1120_n 0.0100696f $X=-1.345 $Y=0 $X2=4.06
+ $Y2=2.765
cc_149 N_GND_M1010_b N_A_687_115#_c_1121_n 0.00339088f $X=-1.345 $Y=0 $X2=3.645
+ $Y2=2.765
cc_150 N_GND_M1010_b N_A_687_115#_c_1122_n 0.00425131f $X=-1.345 $Y=0 $X2=4.145
+ $Y2=2.22
cc_151 N_GND_M1010_b N_A_687_115#_c_1123_n 0.00270174f $X=-1.345 $Y=0 $X2=4.95
+ $Y2=2.765
cc_152 N_GND_M1010_b N_A_963_115#_M1008_g 0.0346079f $X=-1.345 $Y=0 $X2=6.015
+ $Y2=1.075
cc_153 N_GND_c_62_p N_A_963_115#_M1008_g 0.0103278f $X=5.73 $Y=0.825 $X2=6.015
+ $Y2=1.075
cc_154 GND N_A_963_115#_M1008_g 0.00468827f $X=5.7 $Y=0.2 $X2=6.015 $Y2=1.075
cc_155 N_GND_M1010_b N_A_963_115#_c_1234_n 0.0369919f $X=-1.345 $Y=0 $X2=6.05
+ $Y2=2.1
cc_156 N_GND_M1010_b N_A_963_115#_c_1235_n 0.0470206f $X=-1.345 $Y=0 $X2=6.032
+ $Y2=2.81
cc_157 N_GND_M1010_b N_A_963_115#_c_1236_n 0.0076653f $X=-1.345 $Y=0 $X2=6.032
+ $Y2=2.96
cc_158 N_GND_M1010_b N_A_963_115#_c_1237_n 0.00711704f $X=-1.345 $Y=0 $X2=4.94
+ $Y2=0.825
cc_159 N_GND_c_61_p N_A_963_115#_c_1237_n 0.00736239f $X=5.645 $Y=0.152 $X2=4.94
+ $Y2=0.825
cc_160 GND N_A_963_115#_c_1237_n 0.00476261f $X=5.7 $Y=0.2 $X2=4.94 $Y2=0.825
cc_161 N_GND_M1010_b N_A_963_115#_c_1240_n 0.00258316f $X=-1.345 $Y=0 $X2=5.205
+ $Y2=1.935
cc_162 N_GND_M1010_b N_A_963_115#_c_1241_n 0.0037072f $X=-1.345 $Y=0 $X2=5.025
+ $Y2=1.935
cc_163 N_GND_M1010_b N_A_963_115#_c_1242_n 0.0215129f $X=-1.345 $Y=0 $X2=6.025
+ $Y2=1.935
cc_164 N_GND_c_62_p N_A_963_115#_c_1242_n 0.00704977f $X=5.73 $Y=0.825 $X2=6.025
+ $Y2=1.935
cc_165 N_GND_M1010_b N_A_963_115#_c_1244_n 0.00590548f $X=-1.345 $Y=0 $X2=5.29
+ $Y2=1.935
cc_166 N_GND_M1010_b N_A_963_115#_c_1245_n 0.00579444f $X=-1.345 $Y=0 $X2=5.33
+ $Y2=3.545
cc_167 N_GND_M1010_b N_A_963_115#_c_1246_n 0.00148267f $X=-1.345 $Y=0 $X2=6.11
+ $Y2=1.935
cc_168 N_GND_M1010_b N_A_856_115#_c_1309_n 0.00156053f $X=-1.345 $Y=0 $X2=4.42
+ $Y2=0.825
cc_169 N_GND_c_61_p N_A_856_115#_c_1309_n 0.00757793f $X=5.645 $Y=0.152 $X2=4.42
+ $Y2=0.825
cc_170 GND N_A_856_115#_c_1309_n 0.00476261f $X=5.7 $Y=0.2 $X2=4.42 $Y2=0.825
cc_171 N_GND_M1010_b N_A_856_115#_c_1312_n 0.045388f $X=-1.345 $Y=0 $X2=4.485
+ $Y2=1.85
cc_172 N_GND_M1010_b N_A_856_115#_c_1313_n 0.00370735f $X=-1.345 $Y=0 $X2=4.452
+ $Y2=1.595
cc_173 N_GND_M1010_b N_ECK_c_1343_n 0.00913846f $X=-1.345 $Y=0 $X2=6.23
+ $Y2=0.825
cc_174 N_GND_c_62_p N_ECK_c_1343_n 0.0187614f $X=5.73 $Y=0.825 $X2=6.23
+ $Y2=0.825
cc_175 GND N_ECK_c_1343_n 0.00476261f $X=5.7 $Y=0.2 $X2=6.23 $Y2=0.825
cc_176 N_GND_M1010_b N_ECK_c_1346_n 0.0167615f $X=-1.345 $Y=0 $X2=6.23 $Y2=2.59
cc_177 N_GND_M1010_b ECK 0.0396909f $X=-1.345 $Y=0 $X2=6.225 $Y2=2.215
cc_178 N_GND_M1010_b N_ECK_c_1348_n 0.0121289f $X=-1.345 $Y=0 $X2=6.23 $Y2=1.48
cc_179 N_GND_c_62_p N_ECK_c_1348_n 0.00119317f $X=5.73 $Y=0.825 $X2=6.23
+ $Y2=1.48
cc_180 N_GND_M1010_b N_ECK_c_1350_n 0.0141494f $X=-1.345 $Y=0 $X2=6.23 $Y2=2.59
cc_181 N_VDD_M1025_b N_SE_M1025_g 0.0246289f $X=-1.345 $Y=2.905 $X2=-0.825
+ $Y2=4.585
cc_182 N_VDD_c_182_p N_SE_M1025_g 0.00606474f $X=-0.335 $Y=6.507 $X2=-0.825
+ $Y2=4.585
cc_183 VDD N_SE_M1025_g 0.00468827f $X=5.705 $Y=6.465 $X2=-0.825 $Y2=4.585
cc_184 N_VDD_M1025_b N_SE_c_309_n 0.00408216f $X=-1.345 $Y=2.905 $X2=-0.649
+ $Y2=2.96
cc_185 N_VDD_M1025_b N_SE_X27_noxref_CONDUCTOR 0.00838127f $X=-1.345 $Y=2.905
+ $X2=-0.654 $Y2=2.96
cc_186 N_VDD_M1025_b N_E_M1007_g 0.0199366f $X=-1.345 $Y=2.905 $X2=-0.465
+ $Y2=4.585
cc_187 N_VDD_c_182_p N_E_M1007_g 0.00606474f $X=-0.335 $Y=6.507 $X2=-0.465
+ $Y2=4.585
cc_188 N_VDD_c_188_p N_E_M1007_g 0.00713292f $X=-0.249 $Y=4.135 $X2=-0.465
+ $Y2=4.585
cc_189 VDD N_E_M1007_g 0.00468827f $X=5.705 $Y=6.465 $X2=-0.465 $Y2=4.585
cc_190 N_VDD_M1025_b N_E_c_355_n 0.007742f $X=-1.345 $Y=2.905 $X2=-0.309
+ $Y2=2.755
cc_191 N_VDD_M1007_d N_E_c_356_n 0.00499194f $X=-0.39 $Y=3.085 $X2=-0.309
+ $Y2=2.755
cc_192 N_VDD_M1025_b N_E_c_356_n 0.00192816f $X=-1.345 $Y=2.905 $X2=-0.309
+ $Y2=2.755
cc_193 N_VDD_c_188_p N_E_c_356_n 0.00252874f $X=-0.249 $Y=4.135 $X2=-0.309
+ $Y2=2.755
cc_194 N_VDD_M1007_d E 0.00722851f $X=-0.39 $Y=3.085 $X2=-0.31 $Y2=3.335
cc_195 N_VDD_c_188_p E 0.00522047f $X=-0.249 $Y=4.135 $X2=-0.31 $Y2=3.335
cc_196 N_VDD_M1025_b N_A_86_337#_c_406_n 0.02482f $X=-1.345 $Y=2.905 $X2=0.53
+ $Y2=2.975
cc_197 N_VDD_c_188_p N_A_86_337#_c_406_n 0.00742312f $X=-0.249 $Y=4.135 $X2=0.53
+ $Y2=2.975
cc_198 N_VDD_c_198_p N_A_86_337#_c_406_n 0.00606474f $X=0.685 $Y=6.507 $X2=0.53
+ $Y2=2.975
cc_199 N_VDD_c_199_p N_A_86_337#_c_406_n 0.00354579f $X=0.77 $Y=3.795 $X2=0.53
+ $Y2=2.975
cc_200 VDD N_A_86_337#_c_406_n 0.00468827f $X=5.705 $Y=6.465 $X2=0.53 $Y2=2.975
cc_201 N_VDD_M1025_b N_A_86_337#_c_408_n 0.00184258f $X=-1.345 $Y=2.905
+ $X2=0.565 $Y2=3.1
cc_202 N_VDD_M1022_d N_A_86_337#_c_421_n 0.00444289f $X=0.63 $Y=3.085 $X2=1.475
+ $Y2=3.185
cc_203 N_VDD_c_199_p N_A_86_337#_c_421_n 0.00946335f $X=0.77 $Y=3.795 $X2=1.475
+ $Y2=3.185
cc_204 N_VDD_M1025_b N_A_86_337#_c_423_n 0.00313975f $X=-1.345 $Y=2.905
+ $X2=1.645 $Y2=3.455
cc_205 N_VDD_c_205_p N_A_86_337#_c_423_n 0.0151591f $X=2.435 $Y=6.507 $X2=1.645
+ $Y2=3.455
cc_206 VDD N_A_86_337#_c_423_n 0.00958198f $X=5.705 $Y=6.465 $X2=1.645 $Y2=3.455
cc_207 N_VDD_M1025_b N_A_N233_617#_M1002_g 0.019736f $X=-1.345 $Y=2.905
+ $X2=0.985 $Y2=4.585
cc_208 N_VDD_c_199_p N_A_N233_617#_M1002_g 0.00354579f $X=0.77 $Y=3.795
+ $X2=0.985 $Y2=4.585
cc_209 N_VDD_c_205_p N_A_N233_617#_M1002_g 0.00606474f $X=2.435 $Y=6.507
+ $X2=0.985 $Y2=4.585
cc_210 VDD N_A_N233_617#_M1002_g 0.00468827f $X=5.705 $Y=6.465 $X2=0.985
+ $Y2=4.585
cc_211 N_VDD_M1025_b N_A_N233_617#_c_490_n 0.00981538f $X=-1.345 $Y=2.905
+ $X2=-1.039 $Y2=2.59
cc_212 N_VDD_c_182_p N_A_N233_617#_c_490_n 0.00736239f $X=-0.335 $Y=6.507
+ $X2=-1.039 $Y2=2.59
cc_213 VDD N_A_N233_617#_c_490_n 0.00476261f $X=5.705 $Y=6.465 $X2=-1.039
+ $Y2=2.59
cc_214 N_VDD_M1025_b N_CK_M1004_g 0.0195114f $X=-1.345 $Y=2.905 $X2=1.345
+ $Y2=4.585
cc_215 N_VDD_c_205_p N_CK_M1004_g 0.00606474f $X=2.435 $Y=6.507 $X2=1.345
+ $Y2=4.585
cc_216 VDD N_CK_M1004_g 0.00468827f $X=5.705 $Y=6.465 $X2=1.345 $Y2=4.585
cc_217 N_VDD_M1025_b N_CK_M1000_g 0.0236813f $X=-1.345 $Y=2.905 $X2=2.735
+ $Y2=4.585
cc_218 N_VDD_c_218_p N_CK_M1000_g 0.00354579f $X=2.52 $Y=3.455 $X2=2.735
+ $Y2=4.585
cc_219 N_VDD_c_219_p N_CK_M1000_g 0.00606474f $X=3.905 $Y=6.507 $X2=2.735
+ $Y2=4.585
cc_220 VDD N_CK_M1000_g 0.00468827f $X=5.705 $Y=6.465 $X2=2.735 $Y2=4.585
cc_221 N_VDD_M1025_b N_CK_M1005_g 0.0187476f $X=-1.345 $Y=2.905 $X2=5.585
+ $Y2=4.585
cc_222 N_VDD_c_222_p N_CK_M1005_g 0.00606474f $X=5.715 $Y=6.507 $X2=5.585
+ $Y2=4.585
cc_223 N_VDD_c_223_p N_CK_M1005_g 0.00354579f $X=5.8 $Y=3.795 $X2=5.585
+ $Y2=4.585
cc_224 VDD N_CK_M1005_g 0.00468827f $X=5.705 $Y=6.465 $X2=5.585 $Y2=4.585
cc_225 N_VDD_M1025_b N_CK_c_605_n 0.00547126f $X=-1.345 $Y=2.905 $X2=1.405
+ $Y2=2.765
cc_226 N_VDD_M1025_b N_CK_c_611_n 0.00395347f $X=-1.345 $Y=2.905 $X2=2.762
+ $Y2=2.935
cc_227 N_VDD_M1025_b N_CK_c_617_n 0.00170274f $X=-1.345 $Y=2.905 $X2=5.63
+ $Y2=2.425
cc_228 N_VDD_M1025_b N_CK_c_620_n 0.0415575f $X=-1.345 $Y=2.905 $X2=5.485
+ $Y2=2.96
cc_229 N_VDD_c_218_p N_CK_c_620_n 0.0090257f $X=2.52 $Y=3.455 $X2=5.485 $Y2=2.96
cc_230 N_VDD_c_230_p N_CK_c_620_n 0.00183313f $X=3.99 $Y=3.455 $X2=5.485
+ $Y2=2.96
cc_231 N_VDD_M1025_b N_CK_c_621_n 9.01251e-19 $X=-1.345 $Y=2.905 $X2=1.405
+ $Y2=2.765
cc_232 N_VDD_M1025_b N_CK_c_623_n 0.0055239f $X=-1.345 $Y=2.905 $X2=5.63
+ $Y2=2.96
cc_233 N_VDD_c_223_p N_CK_c_623_n 0.00240671f $X=5.8 $Y=3.795 $X2=5.63 $Y2=2.96
cc_234 N_VDD_M1025_b N_A_254_89#_M1013_g 0.0188823f $X=-1.345 $Y=2.905 $X2=1.945
+ $Y2=4.585
cc_235 N_VDD_c_205_p N_A_254_89#_M1013_g 0.00606474f $X=2.435 $Y=6.507 $X2=1.945
+ $Y2=4.585
cc_236 VDD N_A_254_89#_M1013_g 0.00468827f $X=5.705 $Y=6.465 $X2=1.945 $Y2=4.585
cc_237 N_VDD_M1025_b N_A_254_89#_c_794_n 0.00496173f $X=-1.345 $Y=2.905
+ $X2=1.885 $Y2=2.765
cc_238 N_VDD_M1025_b N_A_254_89#_c_796_n 7.56914e-19 $X=-1.345 $Y=2.905
+ $X2=1.885 $Y2=2.59
cc_239 N_VDD_M1025_b N_A_254_89#_c_800_n 0.00628451f $X=-1.345 $Y=2.905 $X2=2.95
+ $Y2=2.59
cc_240 N_VDD_c_219_p N_A_254_89#_c_800_n 0.00754714f $X=3.905 $Y=6.507 $X2=2.95
+ $Y2=2.59
cc_241 VDD N_A_254_89#_c_800_n 0.00476261f $X=5.705 $Y=6.465 $X2=2.95 $Y2=2.59
cc_242 N_VDD_M1025_b N_A_43_115#_M1014_g 0.0182457f $X=-1.345 $Y=2.905 $X2=2.305
+ $Y2=4.585
cc_243 N_VDD_c_205_p N_A_43_115#_M1014_g 0.00606474f $X=2.435 $Y=6.507 $X2=2.305
+ $Y2=4.585
cc_244 N_VDD_c_218_p N_A_43_115#_M1014_g 0.00354579f $X=2.52 $Y=3.455 $X2=2.305
+ $Y2=4.585
cc_245 VDD N_A_43_115#_M1014_g 0.00468827f $X=5.705 $Y=6.465 $X2=2.305 $Y2=4.585
cc_246 N_VDD_M1025_b N_A_43_115#_c_936_n 0.0278214f $X=-1.345 $Y=2.905 $X2=3.75
+ $Y2=3.005
cc_247 N_VDD_c_219_p N_A_43_115#_c_936_n 0.00606474f $X=3.905 $Y=6.507 $X2=3.75
+ $Y2=3.005
cc_248 N_VDD_c_230_p N_A_43_115#_c_936_n 0.00383121f $X=3.99 $Y=3.455 $X2=3.75
+ $Y2=3.005
cc_249 VDD N_A_43_115#_c_936_n 0.00468827f $X=5.705 $Y=6.465 $X2=3.75 $Y2=3.005
cc_250 N_VDD_M1025_b N_A_43_115#_c_937_n 0.00930728f $X=-1.345 $Y=2.905
+ $X2=0.225 $Y2=2.22
cc_251 N_VDD_M1025_b N_A_43_115#_c_960_n 0.00156053f $X=-1.345 $Y=2.905 $X2=0.34
+ $Y2=4.135
cc_252 N_VDD_c_188_p N_A_43_115#_c_960_n 0.0794385f $X=-0.249 $Y=4.135 $X2=0.34
+ $Y2=4.135
cc_253 N_VDD_c_198_p N_A_43_115#_c_960_n 0.00757793f $X=0.685 $Y=6.507 $X2=0.34
+ $Y2=4.135
cc_254 VDD N_A_43_115#_c_960_n 0.00476261f $X=5.705 $Y=6.465 $X2=0.34 $Y2=4.135
cc_255 N_VDD_M1025_b N_A_43_115#_c_964_n 0.00962373f $X=-1.345 $Y=2.905 $X2=0.34
+ $Y2=3.795
cc_256 N_VDD_c_188_p N_A_43_115#_c_964_n 0.00355502f $X=-0.249 $Y=4.135 $X2=0.34
+ $Y2=3.795
cc_257 N_VDD_M1025_b N_A_687_115#_M1009_g 0.0231061f $X=-1.345 $Y=2.905
+ $X2=4.205 $Y2=4.585
cc_258 N_VDD_c_230_p N_A_687_115#_M1009_g 0.00383121f $X=3.99 $Y=3.455 $X2=4.205
+ $Y2=4.585
cc_259 N_VDD_c_259_p N_A_687_115#_M1009_g 0.00606474f $X=4.855 $Y=6.507
+ $X2=4.205 $Y2=4.585
cc_260 N_VDD_c_260_p N_A_687_115#_M1009_g 0.00742269f $X=4.94 $Y=4.135 $X2=4.205
+ $Y2=4.585
cc_261 VDD N_A_687_115#_M1009_g 0.00468827f $X=5.705 $Y=6.465 $X2=4.205
+ $Y2=4.585
cc_262 N_VDD_M1025_b N_A_687_115#_M1021_g 0.0203786f $X=-1.345 $Y=2.905
+ $X2=5.155 $Y2=4.585
cc_263 N_VDD_c_260_p N_A_687_115#_M1021_g 0.00713292f $X=4.94 $Y=4.135 $X2=5.155
+ $Y2=4.585
cc_264 N_VDD_c_222_p N_A_687_115#_M1021_g 0.00606474f $X=5.715 $Y=6.507
+ $X2=5.155 $Y2=4.585
cc_265 VDD N_A_687_115#_M1021_g 0.00468827f $X=5.705 $Y=6.465 $X2=5.155
+ $Y2=4.585
cc_266 N_VDD_M1025_b N_A_687_115#_c_1112_n 0.0100684f $X=-1.345 $Y=2.905
+ $X2=5.155 $Y2=2.765
cc_267 N_VDD_M1025_b N_A_687_115#_c_1116_n 0.00551401f $X=-1.345 $Y=2.905
+ $X2=3.56 $Y2=3.33
cc_268 N_VDD_c_219_p N_A_687_115#_c_1116_n 0.00745733f $X=3.905 $Y=6.507
+ $X2=3.56 $Y2=3.33
cc_269 N_VDD_c_230_p N_A_687_115#_c_1116_n 0.00465312f $X=3.99 $Y=3.455 $X2=3.56
+ $Y2=3.33
cc_270 VDD N_A_687_115#_c_1116_n 0.00476261f $X=5.705 $Y=6.465 $X2=3.56 $Y2=3.33
cc_271 N_VDD_c_230_p N_A_687_115#_c_1120_n 0.00435485f $X=3.99 $Y=3.455 $X2=4.06
+ $Y2=2.765
cc_272 N_VDD_M1021_s N_A_687_115#_c_1123_n 0.00763092f $X=4.815 $Y=3.085
+ $X2=4.95 $Y2=2.765
cc_273 N_VDD_M1025_b N_A_687_115#_c_1123_n 0.00159171f $X=-1.345 $Y=2.905
+ $X2=4.95 $Y2=2.765
cc_274 N_VDD_c_260_p N_A_687_115#_c_1123_n 0.00370742f $X=4.94 $Y=4.135 $X2=4.95
+ $Y2=2.765
cc_275 N_VDD_M1020_d N_A_687_115#_c_1142_n 0.00474309f $X=3.85 $Y=3.085
+ $X2=4.805 $Y2=3.33
cc_276 N_VDD_M1021_s N_A_687_115#_c_1142_n 0.00648605f $X=4.815 $Y=3.085
+ $X2=4.805 $Y2=3.33
cc_277 N_VDD_M1025_b N_A_687_115#_c_1142_n 0.012701f $X=-1.345 $Y=2.905
+ $X2=4.805 $Y2=3.33
cc_278 N_VDD_c_230_p N_A_687_115#_c_1142_n 0.0183176f $X=3.99 $Y=3.455 $X2=4.805
+ $Y2=3.33
cc_279 N_VDD_c_260_p N_A_687_115#_c_1142_n 0.00434783f $X=4.94 $Y=4.135
+ $X2=4.805 $Y2=3.33
cc_280 N_VDD_M1025_b N_A_687_115#_c_1147_n 0.00341488f $X=-1.345 $Y=2.905
+ $X2=3.7 $Y2=3.33
cc_281 N_VDD_c_230_p N_A_687_115#_c_1147_n 0.00161445f $X=3.99 $Y=3.455 $X2=3.7
+ $Y2=3.33
cc_282 N_VDD_M1025_b N_A_963_115#_c_1236_n 0.0267233f $X=-1.345 $Y=2.905
+ $X2=6.032 $Y2=2.96
cc_283 N_VDD_c_223_p N_A_963_115#_c_1236_n 0.00354579f $X=5.8 $Y=3.795 $X2=6.032
+ $Y2=2.96
cc_284 N_VDD_c_284_p N_A_963_115#_c_1236_n 0.00606474f $X=5.8 $Y=6.507 $X2=6.032
+ $Y2=2.96
cc_285 VDD N_A_963_115#_c_1236_n 0.00468827f $X=5.705 $Y=6.465 $X2=6.032
+ $Y2=2.96
cc_286 N_VDD_M1025_b N_A_963_115#_c_1251_n 0.00155118f $X=-1.345 $Y=2.905
+ $X2=5.37 $Y2=3.795
cc_287 N_VDD_c_222_p N_A_963_115#_c_1251_n 0.0075556f $X=5.715 $Y=6.507 $X2=5.37
+ $Y2=3.795
cc_288 VDD N_A_963_115#_c_1251_n 0.00475776f $X=5.705 $Y=6.465 $X2=5.37
+ $Y2=3.795
cc_289 N_VDD_M1025_b N_A_963_115#_c_1245_n 6.57756e-19 $X=-1.345 $Y=2.905
+ $X2=5.33 $Y2=3.545
cc_290 N_VDD_M1025_b N_A_856_115#_c_1314_n 0.00156053f $X=-1.345 $Y=2.905
+ $X2=4.42 $Y2=3.455
cc_291 N_VDD_c_259_p N_A_856_115#_c_1314_n 0.00757793f $X=4.855 $Y=6.507
+ $X2=4.42 $Y2=3.455
cc_292 N_VDD_c_260_p N_A_856_115#_c_1314_n 0.0939805f $X=4.94 $Y=4.135 $X2=4.42
+ $Y2=3.455
cc_293 VDD N_A_856_115#_c_1314_n 0.00476261f $X=5.705 $Y=6.465 $X2=4.42
+ $Y2=3.455
cc_294 N_VDD_M1025_b N_A_856_115#_c_1312_n 0.00506395f $X=-1.345 $Y=2.905
+ $X2=4.485 $Y2=1.85
cc_295 N_VDD_M1025_b N_A_856_115#_c_1319_n 0.00162237f $X=-1.345 $Y=2.905
+ $X2=4.452 $Y2=3.33
cc_296 N_VDD_c_230_p N_A_856_115#_c_1319_n 0.00395367f $X=3.99 $Y=3.455
+ $X2=4.452 $Y2=3.33
cc_297 N_VDD_M1025_b N_ECK_c_1346_n 0.0100094f $X=-1.345 $Y=2.905 $X2=6.23
+ $Y2=2.59
cc_298 N_VDD_c_284_p N_ECK_c_1346_n 0.00757793f $X=5.8 $Y=6.507 $X2=6.23
+ $Y2=2.59
cc_299 VDD N_ECK_c_1346_n 0.00476261f $X=5.705 $Y=6.465 $X2=6.23 $Y2=2.59
cc_300 N_SE_X27_noxref_CONDUCTOR N_E_M1007_g 0.00231474f $X=-0.654 $Y=2.96
+ $X2=-0.465 $Y2=4.585
cc_301 N_SE_M1010_g N_E_M1018_g 0.060867f $X=-0.825 $Y=1.075 $X2=-0.395
+ $Y2=1.075
cc_302 N_SE_c_307_n N_E_M1018_g 0.00368334f $X=-0.735 $Y=2.09 $X2=-0.395
+ $Y2=1.075
cc_303 N_SE_c_309_n N_E_M1018_g 0.00800257f $X=-0.649 $Y=2.96 $X2=-0.395
+ $Y2=1.075
cc_304 N_SE_M1025_g N_E_c_355_n 0.217221f $X=-0.825 $Y=4.585 $X2=-0.309
+ $Y2=2.755
cc_305 N_SE_c_309_n N_E_c_355_n 0.00287105f $X=-0.649 $Y=2.96 $X2=-0.309
+ $Y2=2.755
cc_306 N_SE_X27_noxref_CONDUCTOR N_E_c_355_n 0.00130895f $X=-0.654 $Y=2.96
+ $X2=-0.309 $Y2=2.755
cc_307 N_SE_M1025_g N_E_c_356_n 0.00140248f $X=-0.825 $Y=4.585 $X2=-0.309
+ $Y2=2.755
cc_308 N_SE_c_309_n N_E_c_356_n 0.0302217f $X=-0.649 $Y=2.96 $X2=-0.309
+ $Y2=2.755
cc_309 N_SE_X27_noxref_CONDUCTOR N_E_c_356_n 0.00643447f $X=-0.654 $Y=2.96
+ $X2=-0.309 $Y2=2.755
cc_310 N_SE_M1025_g E 0.00297933f $X=-0.825 $Y=4.585 $X2=-0.31 $Y2=3.335
cc_311 N_SE_X27_noxref_CONDUCTOR E 0.0050603f $X=-0.654 $Y=2.96 $X2=-0.31
+ $Y2=3.335
cc_312 N_SE_M1025_g N_A_N233_617#_c_490_n 0.016616f $X=-0.825 $Y=4.585
+ $X2=-1.039 $Y2=2.59
cc_313 N_SE_c_305_n N_A_N233_617#_c_490_n 0.00138434f $X=-0.884 $Y=2.09
+ $X2=-1.039 $Y2=2.59
cc_314 N_SE_c_307_n N_A_N233_617#_c_490_n 0.00308264f $X=-0.735 $Y=2.09
+ $X2=-1.039 $Y2=2.59
cc_315 N_SE_c_309_n N_A_N233_617#_c_490_n 0.0294278f $X=-0.649 $Y=2.96
+ $X2=-1.039 $Y2=2.59
cc_316 N_SE_X27_noxref_CONDUCTOR N_A_N233_617#_c_490_n 0.00774605f $X=-0.654
+ $Y=2.96 $X2=-1.039 $Y2=2.59
cc_317 N_SE_M1010_g N_A_N233_617#_c_491_n 0.00231637f $X=-0.825 $Y=1.075
+ $X2=-0.609 $Y2=0.825
cc_318 N_SE_c_307_n N_A_N233_617#_c_491_n 0.00336259f $X=-0.735 $Y=2.09
+ $X2=-0.609 $Y2=0.825
cc_319 N_SE_M1025_g N_A_N233_617#_c_495_n 0.00412998f $X=-0.825 $Y=4.585
+ $X2=-0.71 $Y2=2.59
cc_320 N_SE_c_307_n N_A_N233_617#_c_495_n 0.00523952f $X=-0.735 $Y=2.09
+ $X2=-0.71 $Y2=2.59
cc_321 N_SE_c_309_n N_A_N233_617#_c_495_n 0.0040117f $X=-0.649 $Y=2.96 $X2=-0.71
+ $Y2=2.59
cc_322 N_SE_X27_noxref_CONDUCTOR N_A_N233_617#_c_495_n 0.0158416f $X=-0.654
+ $Y=2.96 $X2=-0.71 $Y2=2.59
cc_323 N_SE_M1025_g N_A_N233_617#_c_496_n 0.00325397f $X=-0.825 $Y=4.585
+ $X2=-0.895 $Y2=2.59
cc_324 N_SE_c_305_n N_A_N233_617#_c_496_n 0.00301446f $X=-0.884 $Y=2.09
+ $X2=-0.895 $Y2=2.59
cc_325 N_SE_c_307_n N_A_N233_617#_c_496_n 0.00469337f $X=-0.735 $Y=2.09
+ $X2=-0.895 $Y2=2.59
cc_326 N_SE_c_309_n N_A_N233_617#_c_496_n 0.00147755f $X=-0.649 $Y=2.96
+ $X2=-0.895 $Y2=2.59
cc_327 N_SE_X27_noxref_CONDUCTOR N_A_N233_617#_c_496_n 9.25684e-19 $X=-0.654
+ $Y=2.96 $X2=-0.895 $Y2=2.59
cc_328 N_SE_M1010_g N_A_N233_617#_c_497_n 0.00594872f $X=-0.825 $Y=1.075
+ $X2=-0.61 $Y2=2.505
cc_329 N_SE_c_307_n N_A_N233_617#_c_497_n 0.0124433f $X=-0.735 $Y=2.09 $X2=-0.61
+ $Y2=2.505
cc_330 N_SE_c_309_n N_A_N233_617#_c_497_n 0.0178687f $X=-0.649 $Y=2.96 $X2=-0.61
+ $Y2=2.505
cc_331 N_SE_M1010_g N_A_N233_617#_c_498_n 0.0089989f $X=-0.825 $Y=1.075
+ $X2=-0.609 $Y2=1.48
cc_332 N_SE_c_307_n N_A_N233_617#_c_498_n 0.00244196f $X=-0.735 $Y=2.09
+ $X2=-0.609 $Y2=1.48
cc_333 N_SE_c_309_n N_A_N233_617#_c_501_n 0.00954344f $X=-0.649 $Y=2.96
+ $X2=-0.617 $Y2=2.592
cc_334 N_SE_X27_noxref_CONDUCTOR N_A_N233_617#_c_501_n 0.0189236f $X=-0.654
+ $Y=2.96 $X2=-0.617 $Y2=2.592
cc_335 N_E_c_355_n N_A_86_337#_c_405_n 0.00469974f $X=-0.309 $Y=2.755 $X2=0.53
+ $Y2=2.805
cc_336 N_E_c_356_n N_A_N233_617#_c_490_n 0.00350166f $X=-0.309 $Y=2.755
+ $X2=-1.039 $Y2=2.59
cc_337 E N_A_N233_617#_c_490_n 0.00623956f $X=-0.31 $Y=3.335 $X2=-1.039 $Y2=2.59
cc_338 N_E_M1018_g N_A_N233_617#_c_491_n 0.00162674f $X=-0.395 $Y=1.075
+ $X2=-0.609 $Y2=0.825
cc_339 N_E_M1018_g N_A_N233_617#_c_497_n 0.013109f $X=-0.395 $Y=1.075 $X2=-0.61
+ $Y2=2.505
cc_340 N_E_M1018_g N_A_N233_617#_c_498_n 0.00476605f $X=-0.395 $Y=1.075
+ $X2=-0.609 $Y2=1.48
cc_341 N_E_c_355_n N_A_N233_617#_c_501_n 8.20266e-19 $X=-0.309 $Y=2.755
+ $X2=-0.617 $Y2=2.592
cc_342 N_E_M1018_g N_A_N233_617#_c_503_n 0.0081763f $X=-0.395 $Y=1.075 $X2=0.78
+ $Y2=2.595
cc_343 N_E_c_355_n N_A_N233_617#_c_503_n 0.00674587f $X=-0.309 $Y=2.755 $X2=0.78
+ $Y2=2.595
cc_344 N_E_c_356_n N_A_N233_617#_c_503_n 0.0112856f $X=-0.309 $Y=2.755 $X2=0.78
+ $Y2=2.595
cc_345 E N_A_N233_617#_c_503_n 0.012686f $X=-0.31 $Y=3.335 $X2=0.78 $Y2=2.595
cc_346 N_E_M1007_g N_A_43_115#_c_937_n 0.0137937f $X=-0.465 $Y=4.585 $X2=0.225
+ $Y2=2.22
cc_347 N_E_M1018_g N_A_43_115#_c_937_n 0.0254566f $X=-0.395 $Y=1.075 $X2=0.225
+ $Y2=2.22
cc_348 N_E_c_355_n N_A_43_115#_c_937_n 0.00281578f $X=-0.309 $Y=2.755 $X2=0.225
+ $Y2=2.22
cc_349 N_E_c_356_n N_A_43_115#_c_937_n 0.0309935f $X=-0.309 $Y=2.755 $X2=0.225
+ $Y2=2.22
cc_350 E N_A_43_115#_c_937_n 0.00692722f $X=-0.31 $Y=3.335 $X2=0.225 $Y2=2.22
cc_351 N_E_M1018_g N_A_43_115#_c_944_n 0.00130963f $X=-0.395 $Y=1.075 $X2=0.34
+ $Y2=1.395
cc_352 N_E_M1018_g N_A_43_115#_c_948_n 0.00532884f $X=-0.395 $Y=1.075 $X2=0.37
+ $Y2=2.22
cc_353 E A_N150_617# 0.00289505f $X=-0.31 $Y=3.335 $X2=-0.75 $Y2=3.085
cc_354 N_A_86_337#_c_398_n N_A_N233_617#_M1023_g 0.0207333f $X=0.565 $Y=1.85
+ $X2=0.985 $Y2=1.075
cc_355 N_A_86_337#_c_400_n N_A_N233_617#_M1023_g 0.0196577f $X=0.565 $Y=1.685
+ $X2=0.985 $Y2=1.075
cc_356 N_A_86_337#_c_405_n N_A_N233_617#_M1023_g 0.00885564f $X=0.53 $Y=2.805
+ $X2=0.985 $Y2=1.075
cc_357 N_A_86_337#_c_407_n N_A_N233_617#_M1023_g 2.45848e-19 $X=0.565 $Y=1.935
+ $X2=0.985 $Y2=1.075
cc_358 N_A_86_337#_c_408_n N_A_N233_617#_M1023_g 0.00448652f $X=0.565 $Y=3.1
+ $X2=0.985 $Y2=1.075
cc_359 N_A_86_337#_c_409_n N_A_N233_617#_M1023_g 0.0125105f $X=1.025 $Y=1.85
+ $X2=0.985 $Y2=1.075
cc_360 N_A_86_337#_c_411_n N_A_N233_617#_M1023_g 0.00552645f $X=1.11 $Y=1.765
+ $X2=0.985 $Y2=1.075
cc_361 N_A_86_337#_c_434_p N_A_N233_617#_M1023_g 0.00605553f $X=1.195 $Y=1.43
+ $X2=0.985 $Y2=1.075
cc_362 N_A_86_337#_c_405_n N_A_N233_617#_M1002_g 0.00755439f $X=0.53 $Y=2.805
+ $X2=0.985 $Y2=4.585
cc_363 N_A_86_337#_c_406_n N_A_N233_617#_M1002_g 0.0412319f $X=0.53 $Y=2.975
+ $X2=0.985 $Y2=4.585
cc_364 N_A_86_337#_c_408_n N_A_N233_617#_M1002_g 0.00605506f $X=0.565 $Y=3.1
+ $X2=0.985 $Y2=4.585
cc_365 N_A_86_337#_c_421_n N_A_N233_617#_M1002_g 0.0156361f $X=1.475 $Y=3.185
+ $X2=0.985 $Y2=4.585
cc_366 N_A_86_337#_c_405_n N_A_N233_617#_c_489_n 0.0209207f $X=0.53 $Y=2.805
+ $X2=0.925 $Y2=2.425
cc_367 N_A_86_337#_c_408_n N_A_N233_617#_c_489_n 0.00174544f $X=0.565 $Y=3.1
+ $X2=0.925 $Y2=2.425
cc_368 N_A_86_337#_c_409_n N_A_N233_617#_c_489_n 0.00174867f $X=1.025 $Y=1.85
+ $X2=0.925 $Y2=2.425
cc_369 N_A_86_337#_c_421_n N_A_N233_617#_c_489_n 0.00122128f $X=1.475 $Y=3.185
+ $X2=0.925 $Y2=2.425
cc_370 N_A_86_337#_c_405_n N_A_N233_617#_c_494_n 6.09588e-19 $X=0.53 $Y=2.805
+ $X2=0.925 $Y2=2.425
cc_371 N_A_86_337#_c_408_n N_A_N233_617#_c_494_n 0.026399f $X=0.565 $Y=3.1
+ $X2=0.925 $Y2=2.425
cc_372 N_A_86_337#_c_409_n N_A_N233_617#_c_494_n 0.00476537f $X=1.025 $Y=1.85
+ $X2=0.925 $Y2=2.425
cc_373 N_A_86_337#_c_421_n N_A_N233_617#_c_494_n 0.00315222f $X=1.475 $Y=3.185
+ $X2=0.925 $Y2=2.425
cc_374 N_A_86_337#_c_408_n N_A_N233_617#_c_502_n 0.00185593f $X=0.565 $Y=3.1
+ $X2=0.925 $Y2=2.595
cc_375 N_A_86_337#_c_421_n N_A_N233_617#_c_502_n 0.00814733f $X=1.475 $Y=3.185
+ $X2=0.925 $Y2=2.595
cc_376 N_A_86_337#_c_405_n N_A_N233_617#_c_503_n 0.00475993f $X=0.53 $Y=2.805
+ $X2=0.78 $Y2=2.595
cc_377 N_A_86_337#_c_408_n N_A_N233_617#_c_503_n 0.0174958f $X=0.565 $Y=3.1
+ $X2=0.78 $Y2=2.595
cc_378 N_A_86_337#_c_421_n N_A_N233_617#_c_503_n 0.00469772f $X=1.475 $Y=3.185
+ $X2=0.78 $Y2=2.595
cc_379 N_A_86_337#_c_421_n N_CK_M1004_g 0.0154244f $X=1.475 $Y=3.185 $X2=1.345
+ $Y2=4.585
cc_380 N_A_86_337#_c_421_n N_CK_c_605_n 0.00123862f $X=1.475 $Y=3.185 $X2=1.405
+ $Y2=2.765
cc_381 N_A_86_337#_c_454_p N_CK_c_606_n 0.00158944f $X=1.475 $Y=1.43 $X2=1.885
+ $Y2=1.85
cc_382 N_A_86_337#_c_454_p N_CK_c_614_n 0.0139878f $X=1.475 $Y=1.43 $X2=2.785
+ $Y2=1.85
cc_383 N_A_86_337#_c_409_n N_CK_c_616_n 0.0132034f $X=1.025 $Y=1.85 $X2=1.57
+ $Y2=1.85
cc_384 N_A_86_337#_c_454_p N_CK_c_616_n 0.00917449f $X=1.475 $Y=1.43 $X2=1.57
+ $Y2=1.85
cc_385 N_A_86_337#_c_408_n N_CK_c_618_n 0.00406731f $X=0.565 $Y=3.1 $X2=1.485
+ $Y2=2.765
cc_386 N_A_86_337#_c_421_n N_CK_c_618_n 0.0116127f $X=1.475 $Y=3.185 $X2=1.485
+ $Y2=2.765
cc_387 N_A_86_337#_c_408_n N_CK_c_621_n 0.00186527f $X=0.565 $Y=3.1 $X2=1.405
+ $Y2=2.765
cc_388 N_A_86_337#_c_421_n N_CK_c_621_n 0.0242675f $X=1.475 $Y=3.185 $X2=1.405
+ $Y2=2.765
cc_389 N_A_86_337#_c_409_n N_A_254_89#_M1019_g 0.00127357f $X=1.025 $Y=1.85
+ $X2=1.345 $Y2=1.075
cc_390 N_A_86_337#_c_411_n N_A_254_89#_M1019_g 0.00554866f $X=1.11 $Y=1.765
+ $X2=1.345 $Y2=1.075
cc_391 N_A_86_337#_c_454_p N_A_254_89#_M1019_g 0.0165456f $X=1.475 $Y=1.43
+ $X2=1.345 $Y2=1.075
cc_392 N_A_86_337#_c_421_n N_A_254_89#_c_794_n 0.00216878f $X=1.475 $Y=3.185
+ $X2=1.885 $Y2=2.765
cc_393 N_A_86_337#_c_421_n N_A_254_89#_c_796_n 8.86954e-19 $X=1.475 $Y=3.185
+ $X2=1.885 $Y2=2.59
cc_394 N_A_86_337#_c_398_n N_A_43_115#_c_937_n 0.0225097f $X=0.565 $Y=1.85
+ $X2=0.225 $Y2=2.22
cc_395 N_A_86_337#_c_400_n N_A_43_115#_c_937_n 0.00700162f $X=0.565 $Y=1.685
+ $X2=0.225 $Y2=2.22
cc_396 N_A_86_337#_c_406_n N_A_43_115#_c_937_n 0.0128109f $X=0.53 $Y=2.975
+ $X2=0.225 $Y2=2.22
cc_397 N_A_86_337#_c_407_n N_A_43_115#_c_937_n 0.0193917f $X=0.565 $Y=1.935
+ $X2=0.225 $Y2=2.22
cc_398 N_A_86_337#_c_408_n N_A_43_115#_c_937_n 0.0809207f $X=0.565 $Y=3.1
+ $X2=0.225 $Y2=2.22
cc_399 N_A_86_337#_c_472_p N_A_43_115#_c_937_n 0.0133619f $X=0.65 $Y=3.185
+ $X2=0.225 $Y2=2.22
cc_400 N_A_86_337#_c_405_n N_A_43_115#_c_948_n 0.0022955f $X=0.53 $Y=2.805
+ $X2=0.37 $Y2=2.22
cc_401 N_A_86_337#_c_408_n N_A_43_115#_c_948_n 0.00271681f $X=0.565 $Y=3.1
+ $X2=0.37 $Y2=2.22
cc_402 N_A_86_337#_c_398_n N_A_43_115#_c_949_n 0.00127165f $X=0.565 $Y=1.85
+ $X2=2.22 $Y2=2.22
cc_403 N_A_86_337#_c_405_n N_A_43_115#_c_949_n 0.00421591f $X=0.53 $Y=2.805
+ $X2=2.22 $Y2=2.22
cc_404 N_A_86_337#_c_408_n N_A_43_115#_c_949_n 0.0177917f $X=0.565 $Y=3.1
+ $X2=2.22 $Y2=2.22
cc_405 N_A_86_337#_c_409_n N_A_43_115#_c_949_n 0.021201f $X=1.025 $Y=1.85
+ $X2=2.22 $Y2=2.22
cc_406 N_A_86_337#_c_454_p N_A_43_115#_c_949_n 0.00659867f $X=1.475 $Y=1.43
+ $X2=2.22 $Y2=2.22
cc_407 N_A_86_337#_c_421_n A_212_617# 0.00732587f $X=1.475 $Y=3.185 $X2=1.06
+ $Y2=3.085
cc_408 N_A_86_337#_c_411_n A_212_115# 6.51949e-19 $X=1.11 $Y=1.765 $X2=1.06
+ $Y2=0.575
cc_409 N_A_86_337#_c_454_p A_212_115# 9.96211e-19 $X=1.475 $Y=1.43 $X2=1.06
+ $Y2=0.575
cc_410 N_A_86_337#_c_434_p A_212_115# 0.0034593f $X=1.195 $Y=1.43 $X2=1.06
+ $Y2=0.575
cc_411 N_A_N233_617#_M1002_g N_CK_c_605_n 0.215528f $X=0.985 $Y=4.585 $X2=1.405
+ $Y2=2.765
cc_412 N_A_N233_617#_c_494_n N_CK_c_605_n 3.28181e-19 $X=0.925 $Y=2.425
+ $X2=1.405 $Y2=2.765
cc_413 N_A_N233_617#_c_502_n N_CK_c_605_n 0.00103767f $X=0.925 $Y=2.595
+ $X2=1.405 $Y2=2.765
cc_414 N_A_N233_617#_M1023_g N_CK_c_613_n 0.00234107f $X=0.985 $Y=1.075
+ $X2=1.485 $Y2=2.68
cc_415 N_A_N233_617#_c_489_n N_CK_c_613_n 0.00185841f $X=0.925 $Y=2.425
+ $X2=1.485 $Y2=2.68
cc_416 N_A_N233_617#_c_494_n N_CK_c_613_n 0.012661f $X=0.925 $Y=2.425 $X2=1.485
+ $Y2=2.68
cc_417 N_A_N233_617#_c_502_n N_CK_c_613_n 0.00523973f $X=0.925 $Y=2.595
+ $X2=1.485 $Y2=2.68
cc_418 N_A_N233_617#_M1002_g N_CK_c_618_n 0.00165169f $X=0.985 $Y=4.585
+ $X2=1.485 $Y2=2.765
cc_419 N_A_N233_617#_c_502_n N_CK_c_618_n 3.8955e-19 $X=0.925 $Y=2.595 $X2=1.485
+ $Y2=2.765
cc_420 N_A_N233_617#_M1002_g N_CK_c_621_n 0.00138271f $X=0.985 $Y=4.585
+ $X2=1.405 $Y2=2.765
cc_421 N_A_N233_617#_c_502_n N_CK_c_621_n 0.00563153f $X=0.925 $Y=2.595
+ $X2=1.405 $Y2=2.765
cc_422 N_A_N233_617#_M1023_g N_A_254_89#_M1019_g 0.0581908f $X=0.985 $Y=1.075
+ $X2=1.345 $Y2=1.075
cc_423 N_A_N233_617#_c_489_n N_A_254_89#_c_793_n 0.0581908f $X=0.925 $Y=2.425
+ $X2=1.42 $Y2=2.3
cc_424 N_A_N233_617#_c_494_n N_A_254_89#_c_793_n 4.5169e-19 $X=0.925 $Y=2.425
+ $X2=1.42 $Y2=2.3
cc_425 N_A_N233_617#_c_489_n N_A_254_89#_c_795_n 0.00287606f $X=0.925 $Y=2.425
+ $X2=1.885 $Y2=2.6
cc_426 N_A_N233_617#_c_491_n N_A_43_115#_c_937_n 9.77657e-19 $X=-0.609 $Y=0.825
+ $X2=0.225 $Y2=2.22
cc_427 N_A_N233_617#_c_498_n N_A_43_115#_c_937_n 0.00241421f $X=-0.609 $Y=1.48
+ $X2=0.225 $Y2=2.22
cc_428 N_A_N233_617#_c_503_n N_A_43_115#_c_937_n 0.0211452f $X=0.78 $Y=2.595
+ $X2=0.225 $Y2=2.22
cc_429 N_A_N233_617#_c_491_n N_A_43_115#_c_944_n 7.79024e-19 $X=-0.609 $Y=0.825
+ $X2=0.34 $Y2=1.395
cc_430 N_A_N233_617#_c_498_n N_A_43_115#_c_944_n 0.00130395f $X=-0.609 $Y=1.48
+ $X2=0.34 $Y2=1.395
cc_431 N_A_N233_617#_c_503_n N_A_43_115#_c_948_n 0.0259649f $X=0.78 $Y=2.595
+ $X2=0.37 $Y2=2.22
cc_432 N_A_N233_617#_M1023_g N_A_43_115#_c_949_n 0.00314369f $X=0.985 $Y=1.075
+ $X2=2.22 $Y2=2.22
cc_433 N_A_N233_617#_c_489_n N_A_43_115#_c_949_n 0.00237496f $X=0.925 $Y=2.425
+ $X2=2.22 $Y2=2.22
cc_434 N_A_N233_617#_c_494_n N_A_43_115#_c_949_n 0.00482511f $X=0.925 $Y=2.425
+ $X2=2.22 $Y2=2.22
cc_435 N_A_N233_617#_c_502_n N_A_43_115#_c_949_n 0.0229251f $X=0.925 $Y=2.595
+ $X2=2.22 $Y2=2.22
cc_436 N_A_N233_617#_c_503_n N_A_43_115#_c_949_n 0.030411f $X=0.78 $Y=2.595
+ $X2=2.22 $Y2=2.22
cc_437 N_CK_c_606_n N_A_254_89#_M1019_g 0.0122005f $X=1.885 $Y=1.85 $X2=1.345
+ $Y2=1.075
cc_438 N_CK_c_607_n N_A_254_89#_M1019_g 0.0256778f $X=1.885 $Y=1.685 $X2=1.345
+ $Y2=1.075
cc_439 N_CK_c_613_n N_A_254_89#_M1019_g 0.00936286f $X=1.485 $Y=2.68 $X2=1.345
+ $Y2=1.075
cc_440 N_CK_c_616_n N_A_254_89#_M1019_g 0.00439496f $X=1.57 $Y=1.85 $X2=1.345
+ $Y2=1.075
cc_441 N_CK_c_606_n N_A_254_89#_c_792_n 0.0107061f $X=1.885 $Y=1.85 $X2=1.75
+ $Y2=2.3
cc_442 N_CK_c_613_n N_A_254_89#_c_792_n 0.00994433f $X=1.485 $Y=2.68 $X2=1.75
+ $Y2=2.3
cc_443 N_CK_c_614_n N_A_254_89#_c_792_n 0.00524719f $X=2.785 $Y=1.85 $X2=1.75
+ $Y2=2.3
cc_444 N_CK_c_620_n N_A_254_89#_c_792_n 0.00307624f $X=5.485 $Y=2.96 $X2=1.75
+ $Y2=2.3
cc_445 N_CK_c_605_n N_A_254_89#_c_793_n 0.0174061f $X=1.405 $Y=2.765 $X2=1.42
+ $Y2=2.3
cc_446 N_CK_c_613_n N_A_254_89#_c_793_n 0.00254254f $X=1.485 $Y=2.68 $X2=1.42
+ $Y2=2.3
cc_447 N_CK_c_618_n N_A_254_89#_c_793_n 0.00139326f $X=1.485 $Y=2.765 $X2=1.42
+ $Y2=2.3
cc_448 N_CK_c_621_n N_A_254_89#_c_793_n 4.25865e-19 $X=1.405 $Y=2.765 $X2=1.42
+ $Y2=2.3
cc_449 N_CK_M1004_g N_A_254_89#_M1013_g 0.060737f $X=1.345 $Y=4.585 $X2=1.945
+ $Y2=4.585
cc_450 N_CK_c_620_n N_A_254_89#_M1013_g 0.00796817f $X=5.485 $Y=2.96 $X2=1.945
+ $Y2=4.585
cc_451 N_CK_c_605_n N_A_254_89#_c_794_n 0.0216681f $X=1.405 $Y=2.765 $X2=1.885
+ $Y2=2.765
cc_452 N_CK_c_606_n N_A_254_89#_c_794_n 0.00224211f $X=1.885 $Y=1.85 $X2=1.885
+ $Y2=2.765
cc_453 N_CK_c_614_n N_A_254_89#_c_794_n 2.46382e-19 $X=2.785 $Y=1.85 $X2=1.885
+ $Y2=2.765
cc_454 N_CK_c_618_n N_A_254_89#_c_794_n 0.00102234f $X=1.485 $Y=2.765 $X2=1.885
+ $Y2=2.765
cc_455 N_CK_c_620_n N_A_254_89#_c_794_n 0.00270602f $X=5.485 $Y=2.96 $X2=1.885
+ $Y2=2.765
cc_456 N_CK_c_621_n N_A_254_89#_c_794_n 3.83845e-19 $X=1.405 $Y=2.765 $X2=1.885
+ $Y2=2.765
cc_457 N_CK_c_613_n N_A_254_89#_c_795_n 0.00426729f $X=1.485 $Y=2.68 $X2=1.885
+ $Y2=2.6
cc_458 N_CK_c_605_n N_A_254_89#_c_796_n 0.00100395f $X=1.405 $Y=2.765 $X2=1.885
+ $Y2=2.59
cc_459 N_CK_c_606_n N_A_254_89#_c_796_n 8.65047e-19 $X=1.885 $Y=1.85 $X2=1.885
+ $Y2=2.59
cc_460 N_CK_c_613_n N_A_254_89#_c_796_n 0.00783596f $X=1.485 $Y=2.68 $X2=1.885
+ $Y2=2.59
cc_461 N_CK_c_614_n N_A_254_89#_c_796_n 0.00210861f $X=2.785 $Y=1.85 $X2=1.885
+ $Y2=2.59
cc_462 N_CK_c_618_n N_A_254_89#_c_796_n 0.00887913f $X=1.485 $Y=2.765 $X2=1.885
+ $Y2=2.59
cc_463 N_CK_c_620_n N_A_254_89#_c_796_n 0.00873145f $X=5.485 $Y=2.96 $X2=1.885
+ $Y2=2.59
cc_464 N_CK_c_621_n N_A_254_89#_c_796_n 0.00210487f $X=1.405 $Y=2.765 $X2=1.885
+ $Y2=2.59
cc_465 N_CK_M1000_g N_A_254_89#_c_800_n 0.00957264f $X=2.735 $Y=4.585 $X2=2.95
+ $Y2=2.59
cc_466 N_CK_c_610_n N_A_254_89#_c_800_n 0.0224019f $X=2.762 $Y=2.78 $X2=2.95
+ $Y2=2.59
cc_467 N_CK_c_620_n N_A_254_89#_c_800_n 0.0239275f $X=5.485 $Y=2.96 $X2=2.95
+ $Y2=2.59
cc_468 N_CK_c_595_n N_A_254_89#_c_801_n 0.00433902f $X=2.735 $Y=1.665 $X2=3.22
+ $Y2=2.185
cc_469 N_CK_c_599_n N_A_254_89#_c_801_n 0.0037106f $X=2.79 $Y=2.015 $X2=3.22
+ $Y2=2.185
cc_470 N_CK_c_610_n N_A_254_89#_c_801_n 0.00338699f $X=2.762 $Y=2.78 $X2=3.22
+ $Y2=2.185
cc_471 N_CK_c_619_n N_A_254_89#_c_801_n 0.0202967f $X=2.87 $Y=1.85 $X2=3.22
+ $Y2=2.185
cc_472 CK N_A_254_89#_c_801_n 0.00733025f $X=2.87 $Y=1.85 $X2=3.22 $Y2=2.185
cc_473 N_CK_c_599_n N_A_254_89#_c_802_n 0.00350695f $X=2.79 $Y=2.015 $X2=3.22
+ $Y2=1.43
cc_474 N_CK_c_619_n N_A_254_89#_c_802_n 0.00599875f $X=2.87 $Y=1.85 $X2=3.22
+ $Y2=1.43
cc_475 CK N_A_254_89#_c_802_n 0.0023488f $X=2.87 $Y=1.85 $X2=3.22 $Y2=1.43
cc_476 N_CK_c_599_n N_A_254_89#_c_803_n 0.00191656f $X=2.79 $Y=2.015 $X2=3.22
+ $Y2=2.27
cc_477 N_CK_c_610_n N_A_254_89#_c_803_n 0.00357453f $X=2.762 $Y=2.78 $X2=3.22
+ $Y2=2.27
cc_478 N_CK_c_619_n N_A_254_89#_c_803_n 0.00584453f $X=2.87 $Y=1.85 $X2=3.22
+ $Y2=2.27
cc_479 N_CK_c_620_n N_A_254_89#_c_803_n 0.00705533f $X=5.485 $Y=2.96 $X2=3.22
+ $Y2=2.27
cc_480 CK N_A_254_89#_c_803_n 3.48296e-19 $X=2.87 $Y=1.85 $X2=3.22 $Y2=2.27
cc_481 N_CK_c_610_n N_A_254_89#_c_804_n 0.00324642f $X=2.762 $Y=2.78 $X2=2.805
+ $Y2=2.59
cc_482 N_CK_c_611_n N_A_254_89#_c_804_n 0.00109164f $X=2.762 $Y=2.935 $X2=2.805
+ $Y2=2.59
cc_483 N_CK_c_620_n N_A_254_89#_c_804_n 0.0656508f $X=5.485 $Y=2.96 $X2=2.805
+ $Y2=2.59
cc_484 N_CK_c_613_n N_A_254_89#_c_805_n 0.00665965f $X=1.485 $Y=2.68 $X2=2.03
+ $Y2=2.59
cc_485 N_CK_c_620_n N_A_254_89#_c_805_n 0.0251714f $X=5.485 $Y=2.96 $X2=2.03
+ $Y2=2.59
cc_486 N_CK_c_621_n N_A_254_89#_c_805_n 0.00488293f $X=1.405 $Y=2.765 $X2=2.03
+ $Y2=2.59
cc_487 N_CK_c_610_n N_A_254_89#_c_806_n 0.00474676f $X=2.762 $Y=2.78 $X2=2.95
+ $Y2=2.59
cc_488 N_CK_c_620_n N_A_254_89#_c_806_n 0.025192f $X=5.485 $Y=2.96 $X2=2.95
+ $Y2=2.59
cc_489 N_CK_c_595_n N_A_43_115#_M1001_g 0.0278936f $X=2.735 $Y=1.665 $X2=2.305
+ $Y2=1.075
cc_490 N_CK_c_599_n N_A_43_115#_M1001_g 0.00907125f $X=2.79 $Y=2.015 $X2=2.305
+ $Y2=1.075
cc_491 N_CK_c_607_n N_A_43_115#_M1001_g 0.0962296f $X=1.885 $Y=1.685 $X2=2.305
+ $Y2=1.075
cc_492 N_CK_c_613_n N_A_43_115#_M1001_g 0.00249296f $X=1.485 $Y=2.68 $X2=2.305
+ $Y2=1.075
cc_493 N_CK_c_614_n N_A_43_115#_M1001_g 0.0148268f $X=2.785 $Y=1.85 $X2=2.305
+ $Y2=1.075
cc_494 N_CK_c_619_n N_A_43_115#_M1001_g 0.00110864f $X=2.87 $Y=1.85 $X2=2.305
+ $Y2=1.075
cc_495 CK N_A_43_115#_M1001_g 3.04379e-19 $X=2.87 $Y=1.85 $X2=2.305 $Y2=1.075
cc_496 N_CK_c_610_n N_A_43_115#_M1014_g 0.015555f $X=2.762 $Y=2.78 $X2=2.305
+ $Y2=4.585
cc_497 N_CK_c_611_n N_A_43_115#_M1014_g 0.0285866f $X=2.762 $Y=2.935 $X2=2.305
+ $Y2=4.585
cc_498 N_CK_c_620_n N_A_43_115#_M1014_g 0.010536f $X=5.485 $Y=2.96 $X2=2.305
+ $Y2=4.585
cc_499 N_CK_c_610_n N_A_43_115#_c_927_n 0.0211647f $X=2.762 $Y=2.78 $X2=2.365
+ $Y2=2.22
cc_500 N_CK_c_613_n N_A_43_115#_c_927_n 6.23191e-19 $X=1.485 $Y=2.68 $X2=2.365
+ $Y2=2.22
cc_501 N_CK_c_614_n N_A_43_115#_c_927_n 0.00290043f $X=2.785 $Y=1.85 $X2=2.365
+ $Y2=2.22
cc_502 N_CK_c_610_n N_A_43_115#_c_928_n 0.00388214f $X=2.762 $Y=2.78 $X2=3.66
+ $Y2=2.22
cc_503 N_CK_c_599_n N_A_43_115#_c_934_n 0.00457353f $X=2.79 $Y=2.015 $X2=3.75
+ $Y2=1.8
cc_504 N_CK_c_620_n N_A_43_115#_c_936_n 0.00817637f $X=5.485 $Y=2.96 $X2=3.75
+ $Y2=3.005
cc_505 N_CK_c_610_n N_A_43_115#_c_942_n 0.0010711f $X=2.762 $Y=2.78 $X2=2.365
+ $Y2=2.22
cc_506 N_CK_c_613_n N_A_43_115#_c_942_n 0.00297176f $X=1.485 $Y=2.68 $X2=2.365
+ $Y2=2.22
cc_507 N_CK_c_614_n N_A_43_115#_c_942_n 0.0171514f $X=2.785 $Y=1.85 $X2=2.365
+ $Y2=2.22
cc_508 N_CK_c_620_n N_A_43_115#_c_943_n 5.60079e-19 $X=5.485 $Y=2.96 $X2=3.66
+ $Y2=2.22
cc_509 N_CK_c_599_n N_A_43_115#_c_946_n 8.00474e-19 $X=2.79 $Y=2.015 $X2=3.515
+ $Y2=2.22
cc_510 N_CK_c_610_n N_A_43_115#_c_946_n 0.00380983f $X=2.762 $Y=2.78 $X2=3.515
+ $Y2=2.22
cc_511 N_CK_c_614_n N_A_43_115#_c_946_n 0.00511933f $X=2.785 $Y=1.85 $X2=3.515
+ $Y2=2.22
cc_512 N_CK_c_619_n N_A_43_115#_c_946_n 0.00262273f $X=2.87 $Y=1.85 $X2=3.515
+ $Y2=2.22
cc_513 CK N_A_43_115#_c_946_n 0.0344805f $X=2.87 $Y=1.85 $X2=3.515 $Y2=2.22
cc_514 N_CK_c_610_n N_A_43_115#_c_947_n 9.27087e-19 $X=2.762 $Y=2.78 $X2=2.515
+ $Y2=2.22
cc_515 N_CK_c_614_n N_A_43_115#_c_947_n 0.00713297f $X=2.785 $Y=1.85 $X2=2.515
+ $Y2=2.22
cc_516 N_CK_c_605_n N_A_43_115#_c_949_n 3.87465e-19 $X=1.405 $Y=2.765 $X2=2.22
+ $Y2=2.22
cc_517 N_CK_c_606_n N_A_43_115#_c_949_n 0.00411095f $X=1.885 $Y=1.85 $X2=2.22
+ $Y2=2.22
cc_518 N_CK_c_613_n N_A_43_115#_c_949_n 0.0164585f $X=1.485 $Y=2.68 $X2=2.22
+ $Y2=2.22
cc_519 N_CK_c_614_n N_A_43_115#_c_949_n 0.0253127f $X=2.785 $Y=1.85 $X2=2.22
+ $Y2=2.22
cc_520 N_CK_c_618_n N_A_43_115#_c_949_n 0.00245762f $X=1.485 $Y=2.765 $X2=2.22
+ $Y2=2.22
cc_521 N_CK_c_621_n N_A_43_115#_c_949_n 0.0166169f $X=1.405 $Y=2.765 $X2=2.22
+ $Y2=2.22
cc_522 N_CK_c_620_n N_A_43_115#_c_950_n 0.0132278f $X=5.485 $Y=2.96 $X2=3.66
+ $Y2=2.22
cc_523 N_CK_c_620_n N_A_687_115#_M1009_g 0.00905521f $X=5.485 $Y=2.96 $X2=4.205
+ $Y2=4.585
cc_524 N_CK_M1012_g N_A_687_115#_M1015_g 0.129148f $X=5.515 $Y=1.075 $X2=5.155
+ $Y2=1.075
cc_525 N_CK_M1005_g N_A_687_115#_M1015_g 0.0498038f $X=5.585 $Y=4.585 $X2=5.155
+ $Y2=1.075
cc_526 N_CK_c_617_n N_A_687_115#_M1015_g 7.8234e-19 $X=5.63 $Y=2.425 $X2=5.155
+ $Y2=1.075
cc_527 N_CK_c_620_n N_A_687_115#_M1021_g 0.00308514f $X=5.485 $Y=2.96 $X2=5.155
+ $Y2=4.585
cc_528 N_CK_c_620_n N_A_687_115#_c_1112_n 0.0103899f $X=5.485 $Y=2.96 $X2=5.155
+ $Y2=2.765
cc_529 N_CK_c_595_n N_A_687_115#_c_1113_n 0.00199257f $X=2.735 $Y=1.665 $X2=3.56
+ $Y2=0.825
cc_530 N_CK_c_620_n N_A_687_115#_c_1116_n 0.0186937f $X=5.485 $Y=2.96 $X2=3.56
+ $Y2=3.33
cc_531 N_CK_c_620_n N_A_687_115#_c_1120_n 0.0250747f $X=5.485 $Y=2.96 $X2=4.06
+ $Y2=2.765
cc_532 N_CK_c_620_n N_A_687_115#_c_1123_n 0.0178125f $X=5.485 $Y=2.96 $X2=4.95
+ $Y2=2.765
cc_533 N_CK_c_620_n N_A_687_115#_c_1142_n 0.124925f $X=5.485 $Y=2.96 $X2=4.805
+ $Y2=3.33
cc_534 N_CK_c_620_n N_A_687_115#_c_1147_n 0.0252959f $X=5.485 $Y=2.96 $X2=3.7
+ $Y2=3.33
cc_535 N_CK_M1012_g N_A_963_115#_M1008_g 0.0344598f $X=5.515 $Y=1.075 $X2=6.015
+ $Y2=1.075
cc_536 N_CK_M1012_g N_A_963_115#_c_1234_n 0.0102133f $X=5.515 $Y=1.075 $X2=6.05
+ $Y2=2.1
cc_537 N_CK_M1005_g N_A_963_115#_c_1235_n 0.00773101f $X=5.585 $Y=4.585
+ $X2=6.032 $Y2=2.81
cc_538 N_CK_c_612_n N_A_963_115#_c_1235_n 0.0206104f $X=5.63 $Y=2.425 $X2=6.032
+ $Y2=2.81
cc_539 N_CK_c_617_n N_A_963_115#_c_1235_n 0.0033451f $X=5.63 $Y=2.425 $X2=6.032
+ $Y2=2.81
cc_540 N_CK_M1005_g N_A_963_115#_c_1236_n 0.0395234f $X=5.585 $Y=4.585 $X2=6.032
+ $Y2=2.96
cc_541 N_CK_c_617_n N_A_963_115#_c_1236_n 0.00156524f $X=5.63 $Y=2.425 $X2=6.032
+ $Y2=2.96
cc_542 N_CK_c_623_n N_A_963_115#_c_1236_n 0.00425751f $X=5.63 $Y=2.96 $X2=6.032
+ $Y2=2.96
cc_543 N_CK_M1012_g N_A_963_115#_c_1242_n 0.0182215f $X=5.515 $Y=1.075 $X2=6.025
+ $Y2=1.935
cc_544 N_CK_c_612_n N_A_963_115#_c_1242_n 0.00258465f $X=5.63 $Y=2.425 $X2=6.025
+ $Y2=1.935
cc_545 N_CK_c_617_n N_A_963_115#_c_1242_n 0.0101796f $X=5.63 $Y=2.425 $X2=6.025
+ $Y2=1.935
cc_546 N_CK_M1012_g N_A_963_115#_c_1245_n 0.00669183f $X=5.515 $Y=1.075 $X2=5.33
+ $Y2=3.545
cc_547 N_CK_M1005_g N_A_963_115#_c_1245_n 0.013242f $X=5.585 $Y=4.585 $X2=5.33
+ $Y2=3.545
cc_548 N_CK_c_617_n N_A_963_115#_c_1245_n 0.0551821f $X=5.63 $Y=2.425 $X2=5.33
+ $Y2=3.545
cc_549 N_CK_c_620_n N_A_963_115#_c_1245_n 0.0247063f $X=5.485 $Y=2.96 $X2=5.33
+ $Y2=3.545
cc_550 N_CK_c_623_n N_A_963_115#_c_1245_n 0.00247429f $X=5.63 $Y=2.96 $X2=5.33
+ $Y2=3.545
cc_551 N_CK_c_620_n N_A_963_115#_c_1271_n 0.00306237f $X=5.485 $Y=2.96 $X2=5.33
+ $Y2=3.715
cc_552 N_CK_M1012_g N_A_963_115#_c_1246_n 7.99074e-19 $X=5.515 $Y=1.075 $X2=6.11
+ $Y2=1.935
cc_553 N_CK_c_620_n N_A_856_115#_c_1312_n 0.0234059f $X=5.485 $Y=2.96 $X2=4.485
+ $Y2=1.85
cc_554 N_CK_c_620_n N_A_856_115#_c_1319_n 0.00226318f $X=5.485 $Y=2.96 $X2=4.452
+ $Y2=3.33
cc_555 N_CK_c_617_n N_ECK_c_1346_n 0.0153635f $X=5.63 $Y=2.425 $X2=6.23 $Y2=2.59
cc_556 N_CK_c_623_n N_ECK_c_1346_n 0.00701975f $X=5.63 $Y=2.96 $X2=6.23 $Y2=2.59
cc_557 N_CK_c_617_n ECK 0.00695761f $X=5.63 $Y=2.425 $X2=6.225 $Y2=2.215
cc_558 N_CK_M1012_g N_ECK_c_1348_n 7.96664e-19 $X=5.515 $Y=1.075 $X2=6.23
+ $Y2=1.48
cc_559 N_CK_c_612_n N_ECK_c_1350_n 5.70769e-19 $X=5.63 $Y=2.425 $X2=6.23
+ $Y2=2.59
cc_560 N_CK_c_617_n N_ECK_c_1350_n 0.00532157f $X=5.63 $Y=2.425 $X2=6.23
+ $Y2=2.59
cc_561 N_A_254_89#_c_794_n N_A_43_115#_M1014_g 0.215582f $X=1.885 $Y=2.765
+ $X2=2.305 $Y2=4.585
cc_562 N_A_254_89#_c_795_n N_A_43_115#_M1014_g 0.00761683f $X=1.885 $Y=2.6
+ $X2=2.305 $Y2=4.585
cc_563 N_A_254_89#_c_796_n N_A_43_115#_M1014_g 0.00386252f $X=1.885 $Y=2.59
+ $X2=2.305 $Y2=4.585
cc_564 N_A_254_89#_c_804_n N_A_43_115#_M1014_g 0.00582207f $X=2.805 $Y=2.59
+ $X2=2.305 $Y2=4.585
cc_565 N_A_254_89#_c_805_n N_A_43_115#_M1014_g 8.90723e-19 $X=2.03 $Y=2.59
+ $X2=2.305 $Y2=4.585
cc_566 N_A_254_89#_c_806_n N_A_43_115#_M1014_g 2.82435e-19 $X=2.95 $Y=2.59
+ $X2=2.305 $Y2=4.585
cc_567 N_A_254_89#_c_792_n N_A_43_115#_c_927_n 0.00761683f $X=1.75 $Y=2.3
+ $X2=2.365 $Y2=2.22
cc_568 N_A_254_89#_c_803_n N_A_43_115#_c_927_n 4.25625e-19 $X=3.22 $Y=2.27
+ $X2=2.365 $Y2=2.22
cc_569 N_A_254_89#_c_804_n N_A_43_115#_c_927_n 0.00186852f $X=2.805 $Y=2.59
+ $X2=2.365 $Y2=2.22
cc_570 N_A_254_89#_c_800_n N_A_43_115#_c_928_n 5.07664e-19 $X=2.95 $Y=2.59
+ $X2=3.66 $Y2=2.22
cc_571 N_A_254_89#_c_801_n N_A_43_115#_c_928_n 0.00201953f $X=3.22 $Y=2.185
+ $X2=3.66 $Y2=2.22
cc_572 N_A_254_89#_c_803_n N_A_43_115#_c_928_n 0.00174839f $X=3.22 $Y=2.27
+ $X2=3.66 $Y2=2.22
cc_573 N_A_254_89#_c_801_n N_A_43_115#_c_929_n 0.00267523f $X=3.22 $Y=2.185
+ $X2=3.662 $Y2=2.055
cc_574 N_A_254_89#_c_801_n N_A_43_115#_c_934_n 6.33282e-19 $X=3.22 $Y=2.185
+ $X2=3.75 $Y2=1.8
cc_575 N_A_254_89#_c_800_n N_A_43_115#_c_935_n 0.00634397f $X=2.95 $Y=2.59
+ $X2=3.75 $Y2=2.855
cc_576 N_A_254_89#_c_806_n N_A_43_115#_c_935_n 0.00448469f $X=2.95 $Y=2.59
+ $X2=3.75 $Y2=2.855
cc_577 N_A_254_89#_c_792_n N_A_43_115#_c_942_n 6.64388e-19 $X=1.75 $Y=2.3
+ $X2=2.365 $Y2=2.22
cc_578 N_A_254_89#_c_801_n N_A_43_115#_c_942_n 0.00105677f $X=3.22 $Y=2.185
+ $X2=2.365 $Y2=2.22
cc_579 N_A_254_89#_c_803_n N_A_43_115#_c_942_n 0.0040427f $X=3.22 $Y=2.27
+ $X2=2.365 $Y2=2.22
cc_580 N_A_254_89#_c_804_n N_A_43_115#_c_942_n 0.00487271f $X=2.805 $Y=2.59
+ $X2=2.365 $Y2=2.22
cc_581 N_A_254_89#_c_801_n N_A_43_115#_c_943_n 0.00317568f $X=3.22 $Y=2.185
+ $X2=3.66 $Y2=2.22
cc_582 N_A_254_89#_c_803_n N_A_43_115#_c_943_n 0.00780498f $X=3.22 $Y=2.27
+ $X2=3.66 $Y2=2.22
cc_583 N_A_254_89#_c_800_n N_A_43_115#_c_946_n 2.32884e-19 $X=2.95 $Y=2.59
+ $X2=3.515 $Y2=2.22
cc_584 N_A_254_89#_c_801_n N_A_43_115#_c_946_n 0.0108765f $X=3.22 $Y=2.185
+ $X2=3.515 $Y2=2.22
cc_585 N_A_254_89#_c_803_n N_A_43_115#_c_946_n 0.021195f $X=3.22 $Y=2.27
+ $X2=3.515 $Y2=2.22
cc_586 N_A_254_89#_c_804_n N_A_43_115#_c_946_n 0.0233812f $X=2.805 $Y=2.59
+ $X2=3.515 $Y2=2.22
cc_587 N_A_254_89#_c_806_n N_A_43_115#_c_946_n 0.0236535f $X=2.95 $Y=2.59
+ $X2=3.515 $Y2=2.22
cc_588 N_A_254_89#_c_792_n N_A_43_115#_c_947_n 4.70316e-19 $X=1.75 $Y=2.3
+ $X2=2.515 $Y2=2.22
cc_589 N_A_254_89#_c_803_n N_A_43_115#_c_947_n 0.00136849f $X=3.22 $Y=2.27
+ $X2=2.515 $Y2=2.22
cc_590 N_A_254_89#_c_804_n N_A_43_115#_c_947_n 0.0270759f $X=2.805 $Y=2.59
+ $X2=2.515 $Y2=2.22
cc_591 N_A_254_89#_M1019_g N_A_43_115#_c_949_n 0.00255623f $X=1.345 $Y=1.075
+ $X2=2.22 $Y2=2.22
cc_592 N_A_254_89#_c_792_n N_A_43_115#_c_949_n 0.00985983f $X=1.75 $Y=2.3
+ $X2=2.22 $Y2=2.22
cc_593 N_A_254_89#_c_793_n N_A_43_115#_c_949_n 0.00102805f $X=1.42 $Y=2.3
+ $X2=2.22 $Y2=2.22
cc_594 N_A_254_89#_c_796_n N_A_43_115#_c_949_n 9.69764e-19 $X=1.885 $Y=2.59
+ $X2=2.22 $Y2=2.22
cc_595 N_A_254_89#_c_804_n N_A_43_115#_c_949_n 0.0147541f $X=2.805 $Y=2.59
+ $X2=2.22 $Y2=2.22
cc_596 N_A_254_89#_c_805_n N_A_43_115#_c_949_n 0.0242903f $X=2.03 $Y=2.59
+ $X2=2.22 $Y2=2.22
cc_597 N_A_254_89#_c_801_n N_A_43_115#_c_950_n 0.00155231f $X=3.22 $Y=2.185
+ $X2=3.66 $Y2=2.22
cc_598 N_A_254_89#_c_803_n N_A_43_115#_c_950_n 0.00170428f $X=3.22 $Y=2.27
+ $X2=3.66 $Y2=2.22
cc_599 N_A_254_89#_c_797_n N_A_687_115#_c_1113_n 0.0277349f $X=2.95 $Y=0.825
+ $X2=3.56 $Y2=0.825
cc_600 N_A_254_89#_c_801_n N_A_687_115#_c_1113_n 0.0186176f $X=3.22 $Y=2.185
+ $X2=3.56 $Y2=0.825
cc_601 N_A_254_89#_c_802_n N_A_687_115#_c_1113_n 0.0134687f $X=3.22 $Y=1.43
+ $X2=3.56 $Y2=0.825
cc_602 N_A_254_89#_c_800_n N_A_687_115#_c_1116_n 0.111887f $X=2.95 $Y=2.59
+ $X2=3.56 $Y2=3.33
cc_603 N_A_254_89#_c_801_n N_A_687_115#_c_1119_n 0.0137171f $X=3.22 $Y=2.185
+ $X2=3.645 $Y2=1.85
cc_604 N_A_254_89#_c_800_n N_A_687_115#_c_1121_n 0.00701167f $X=2.95 $Y=2.59
+ $X2=3.645 $Y2=2.765
cc_605 N_A_254_89#_c_806_n N_A_687_115#_c_1121_n 6.78681e-19 $X=2.95 $Y=2.59
+ $X2=3.645 $Y2=2.765
cc_606 N_A_254_89#_c_800_n N_A_687_115#_c_1147_n 0.00657714f $X=2.95 $Y=2.59
+ $X2=3.7 $Y2=3.33
cc_607 N_A_43_115#_c_929_n N_A_687_115#_M1006_g 0.00883234f $X=3.662 $Y=2.055
+ $X2=4.205 $Y2=1.075
cc_608 N_A_43_115#_c_930_n N_A_687_115#_M1006_g 0.0248201f $X=3.75 $Y=1.65
+ $X2=4.205 $Y2=1.075
cc_609 N_A_43_115#_c_935_n N_A_687_115#_M1009_g 0.0160728f $X=3.75 $Y=2.855
+ $X2=4.205 $Y2=4.585
cc_610 N_A_43_115#_c_936_n N_A_687_115#_M1009_g 0.0248168f $X=3.75 $Y=3.005
+ $X2=4.205 $Y2=4.585
cc_611 N_A_43_115#_c_928_n N_A_687_115#_c_1111_n 0.0213149f $X=3.66 $Y=2.22
+ $X2=4.145 $Y2=2.22
cc_612 N_A_43_115#_c_943_n N_A_687_115#_c_1111_n 0.00104076f $X=3.66 $Y=2.22
+ $X2=4.145 $Y2=2.22
cc_613 N_A_43_115#_c_950_n N_A_687_115#_c_1111_n 9.12123e-19 $X=3.66 $Y=2.22
+ $X2=4.145 $Y2=2.22
cc_614 N_A_43_115#_c_930_n N_A_687_115#_c_1113_n 0.00804393f $X=3.75 $Y=1.65
+ $X2=3.56 $Y2=0.825
cc_615 N_A_43_115#_c_934_n N_A_687_115#_c_1113_n 0.00367332f $X=3.75 $Y=1.8
+ $X2=3.56 $Y2=0.825
cc_616 N_A_43_115#_c_935_n N_A_687_115#_c_1116_n 0.00580778f $X=3.75 $Y=2.855
+ $X2=3.56 $Y2=3.33
cc_617 N_A_43_115#_c_936_n N_A_687_115#_c_1116_n 0.00752714f $X=3.75 $Y=3.005
+ $X2=3.56 $Y2=3.33
cc_618 N_A_43_115#_c_929_n N_A_687_115#_c_1117_n 0.00765395f $X=3.662 $Y=2.055
+ $X2=4.06 $Y2=1.85
cc_619 N_A_43_115#_c_934_n N_A_687_115#_c_1117_n 0.0108995f $X=3.75 $Y=1.8
+ $X2=4.06 $Y2=1.85
cc_620 N_A_43_115#_c_943_n N_A_687_115#_c_1117_n 0.0093039f $X=3.66 $Y=2.22
+ $X2=4.06 $Y2=1.85
cc_621 N_A_43_115#_c_950_n N_A_687_115#_c_1117_n 0.0037949f $X=3.66 $Y=2.22
+ $X2=4.06 $Y2=1.85
cc_622 N_A_43_115#_c_928_n N_A_687_115#_c_1119_n 0.00303508f $X=3.66 $Y=2.22
+ $X2=3.645 $Y2=1.85
cc_623 N_A_43_115#_c_943_n N_A_687_115#_c_1119_n 0.00899348f $X=3.66 $Y=2.22
+ $X2=3.645 $Y2=1.85
cc_624 N_A_43_115#_c_946_n N_A_687_115#_c_1119_n 0.0011692f $X=3.515 $Y=2.22
+ $X2=3.645 $Y2=1.85
cc_625 N_A_43_115#_c_950_n N_A_687_115#_c_1119_n 0.00331526f $X=3.66 $Y=2.22
+ $X2=3.645 $Y2=1.85
cc_626 N_A_43_115#_c_935_n N_A_687_115#_c_1120_n 0.0127247f $X=3.75 $Y=2.855
+ $X2=4.06 $Y2=2.765
cc_627 N_A_43_115#_c_936_n N_A_687_115#_c_1120_n 0.00248624f $X=3.75 $Y=3.005
+ $X2=4.06 $Y2=2.765
cc_628 N_A_43_115#_c_943_n N_A_687_115#_c_1120_n 0.00455409f $X=3.66 $Y=2.22
+ $X2=4.06 $Y2=2.765
cc_629 N_A_43_115#_c_950_n N_A_687_115#_c_1120_n 0.00140317f $X=3.66 $Y=2.22
+ $X2=4.06 $Y2=2.765
cc_630 N_A_43_115#_c_928_n N_A_687_115#_c_1121_n 0.00271474f $X=3.66 $Y=2.22
+ $X2=3.645 $Y2=2.765
cc_631 N_A_43_115#_c_943_n N_A_687_115#_c_1121_n 0.00449684f $X=3.66 $Y=2.22
+ $X2=3.645 $Y2=2.765
cc_632 N_A_43_115#_c_946_n N_A_687_115#_c_1121_n 0.00100888f $X=3.515 $Y=2.22
+ $X2=3.645 $Y2=2.765
cc_633 N_A_43_115#_c_950_n N_A_687_115#_c_1121_n 0.00142628f $X=3.66 $Y=2.22
+ $X2=3.645 $Y2=2.765
cc_634 N_A_43_115#_c_928_n N_A_687_115#_c_1122_n 0.00116148f $X=3.66 $Y=2.22
+ $X2=4.145 $Y2=2.22
cc_635 N_A_43_115#_c_929_n N_A_687_115#_c_1122_n 0.0022611f $X=3.662 $Y=2.055
+ $X2=4.145 $Y2=2.22
cc_636 N_A_43_115#_c_935_n N_A_687_115#_c_1122_n 0.00558624f $X=3.75 $Y=2.855
+ $X2=4.145 $Y2=2.22
cc_637 N_A_43_115#_c_943_n N_A_687_115#_c_1122_n 0.00887114f $X=3.66 $Y=2.22
+ $X2=4.145 $Y2=2.22
cc_638 N_A_43_115#_c_950_n N_A_687_115#_c_1122_n 0.0035858f $X=3.66 $Y=2.22
+ $X2=4.145 $Y2=2.22
cc_639 N_A_43_115#_c_936_n N_A_687_115#_c_1142_n 0.00783529f $X=3.75 $Y=3.005
+ $X2=4.805 $Y2=3.33
cc_640 N_A_43_115#_c_936_n N_A_687_115#_c_1147_n 0.00124458f $X=3.75 $Y=3.005
+ $X2=3.7 $Y2=3.33
cc_641 N_A_687_115#_M1015_g N_A_963_115#_c_1237_n 0.0158058f $X=5.155 $Y=1.075
+ $X2=4.94 $Y2=0.825
cc_642 N_A_687_115#_M1015_g N_A_963_115#_c_1240_n 0.0160984f $X=5.155 $Y=1.075
+ $X2=5.205 $Y2=1.935
cc_643 N_A_687_115#_c_1112_n N_A_963_115#_c_1240_n 0.00117122f $X=5.155 $Y=2.765
+ $X2=5.205 $Y2=1.935
cc_644 N_A_687_115#_c_1123_n N_A_963_115#_c_1240_n 2.65873e-19 $X=4.95 $Y=2.765
+ $X2=5.205 $Y2=1.935
cc_645 N_A_687_115#_c_1112_n N_A_963_115#_c_1241_n 0.00133457f $X=5.155 $Y=2.765
+ $X2=5.025 $Y2=1.935
cc_646 N_A_687_115#_c_1123_n N_A_963_115#_c_1241_n 0.0055861f $X=4.95 $Y=2.765
+ $X2=5.025 $Y2=1.935
cc_647 N_A_687_115#_M1015_g N_A_963_115#_c_1244_n 0.00322084f $X=5.155 $Y=1.075
+ $X2=5.29 $Y2=1.935
cc_648 N_A_687_115#_M1015_g N_A_963_115#_c_1245_n 0.0157754f $X=5.155 $Y=1.075
+ $X2=5.33 $Y2=3.545
cc_649 N_A_687_115#_M1021_g N_A_963_115#_c_1245_n 0.0135873f $X=5.155 $Y=4.585
+ $X2=5.33 $Y2=3.545
cc_650 N_A_687_115#_c_1112_n N_A_963_115#_c_1245_n 0.00732579f $X=5.155 $Y=2.765
+ $X2=5.33 $Y2=3.545
cc_651 N_A_687_115#_c_1123_n N_A_963_115#_c_1245_n 0.0458366f $X=4.95 $Y=2.765
+ $X2=5.33 $Y2=3.545
cc_652 N_A_687_115#_c_1142_n N_A_963_115#_c_1245_n 0.00818047f $X=4.805 $Y=3.33
+ $X2=5.33 $Y2=3.545
cc_653 N_A_687_115#_M1021_g N_A_963_115#_c_1271_n 0.00884152f $X=5.155 $Y=4.585
+ $X2=5.33 $Y2=3.715
cc_654 N_A_687_115#_c_1142_n N_A_856_115#_M1009_d 0.00413125f $X=4.805 $Y=3.33
+ $X2=4.28 $Y2=3.085
cc_655 N_A_687_115#_M1021_g N_A_856_115#_c_1314_n 0.0150285f $X=5.155 $Y=4.585
+ $X2=4.42 $Y2=3.455
cc_656 N_A_687_115#_c_1123_n N_A_856_115#_c_1314_n 0.00259908f $X=4.95 $Y=2.765
+ $X2=4.42 $Y2=3.455
cc_657 N_A_687_115#_c_1142_n N_A_856_115#_c_1314_n 0.0146401f $X=4.805 $Y=3.33
+ $X2=4.42 $Y2=3.455
cc_658 N_A_687_115#_M1006_g N_A_856_115#_c_1312_n 0.0419193f $X=4.205 $Y=1.075
+ $X2=4.485 $Y2=1.85
cc_659 N_A_687_115#_M1015_g N_A_856_115#_c_1312_n 0.00968085f $X=5.155 $Y=1.075
+ $X2=4.485 $Y2=1.85
cc_660 N_A_687_115#_c_1112_n N_A_856_115#_c_1312_n 0.00298112f $X=5.155 $Y=2.765
+ $X2=4.485 $Y2=1.85
cc_661 N_A_687_115#_c_1117_n N_A_856_115#_c_1312_n 0.0172537f $X=4.06 $Y=1.85
+ $X2=4.485 $Y2=1.85
cc_662 N_A_687_115#_c_1120_n N_A_856_115#_c_1312_n 0.0135849f $X=4.06 $Y=2.765
+ $X2=4.485 $Y2=1.85
cc_663 N_A_687_115#_c_1122_n N_A_856_115#_c_1312_n 0.0536632f $X=4.145 $Y=2.22
+ $X2=4.485 $Y2=1.85
cc_664 N_A_687_115#_c_1123_n N_A_856_115#_c_1312_n 0.0329503f $X=4.95 $Y=2.765
+ $X2=4.485 $Y2=1.85
cc_665 N_A_687_115#_M1006_g N_A_856_115#_c_1313_n 0.00595737f $X=4.205 $Y=1.075
+ $X2=4.452 $Y2=1.595
cc_666 N_A_687_115#_M1015_g N_A_856_115#_c_1313_n 7.46224e-19 $X=5.155 $Y=1.075
+ $X2=4.452 $Y2=1.595
cc_667 N_A_687_115#_M1009_g N_A_856_115#_c_1319_n 0.00322743f $X=4.205 $Y=4.585
+ $X2=4.452 $Y2=3.33
cc_668 N_A_687_115#_c_1142_n N_A_856_115#_c_1319_n 0.0102888f $X=4.805 $Y=3.33
+ $X2=4.452 $Y2=3.33
cc_669 N_A_963_115#_c_1237_n N_A_856_115#_c_1309_n 0.0362893f $X=4.94 $Y=0.825
+ $X2=4.42 $Y2=0.825
cc_670 N_A_963_115#_c_1237_n N_A_856_115#_c_1312_n 0.00408378f $X=4.94 $Y=0.825
+ $X2=4.485 $Y2=1.85
cc_671 N_A_963_115#_c_1241_n N_A_856_115#_c_1312_n 0.0120678f $X=5.025 $Y=1.935
+ $X2=4.485 $Y2=1.85
cc_672 N_A_963_115#_c_1245_n N_A_856_115#_c_1312_n 0.0152471f $X=5.33 $Y=3.545
+ $X2=4.485 $Y2=1.85
cc_673 N_A_963_115#_c_1237_n N_A_856_115#_c_1313_n 0.0203997f $X=4.94 $Y=0.825
+ $X2=4.452 $Y2=1.595
cc_674 N_A_963_115#_M1008_g N_ECK_c_1343_n 0.00580462f $X=6.015 $Y=1.075
+ $X2=6.23 $Y2=0.825
cc_675 N_A_963_115#_c_1234_n N_ECK_c_1343_n 0.00181201f $X=6.05 $Y=2.1 $X2=6.23
+ $Y2=0.825
cc_676 N_A_963_115#_c_1246_n N_ECK_c_1343_n 0.00269883f $X=6.11 $Y=1.935
+ $X2=6.23 $Y2=0.825
cc_677 N_A_963_115#_c_1234_n N_ECK_c_1346_n 0.00130065f $X=6.05 $Y=2.1 $X2=6.23
+ $Y2=2.59
cc_678 N_A_963_115#_c_1235_n N_ECK_c_1346_n 0.0115869f $X=6.032 $Y=2.81 $X2=6.23
+ $Y2=2.59
cc_679 N_A_963_115#_c_1236_n N_ECK_c_1346_n 0.00807887f $X=6.032 $Y=2.96
+ $X2=6.23 $Y2=2.59
cc_680 N_A_963_115#_c_1246_n N_ECK_c_1346_n 0.00127238f $X=6.11 $Y=1.935
+ $X2=6.23 $Y2=2.59
cc_681 N_A_963_115#_M1008_g ECK 0.00406656f $X=6.015 $Y=1.075 $X2=6.225
+ $Y2=2.215
cc_682 N_A_963_115#_c_1234_n ECK 0.00577838f $X=6.05 $Y=2.1 $X2=6.225 $Y2=2.215
cc_683 N_A_963_115#_c_1235_n ECK 0.00892438f $X=6.032 $Y=2.81 $X2=6.225
+ $Y2=2.215
cc_684 N_A_963_115#_c_1242_n ECK 0.00102878f $X=6.025 $Y=1.935 $X2=6.225
+ $Y2=2.215
cc_685 N_A_963_115#_c_1246_n ECK 0.0140245f $X=6.11 $Y=1.935 $X2=6.225 $Y2=2.215
cc_686 N_A_963_115#_M1008_g N_ECK_c_1348_n 0.00680733f $X=6.015 $Y=1.075
+ $X2=6.23 $Y2=1.48
cc_687 N_A_963_115#_c_1246_n N_ECK_c_1348_n 0.00278861f $X=6.11 $Y=1.935
+ $X2=6.23 $Y2=1.48
cc_688 N_A_963_115#_c_1235_n N_ECK_c_1350_n 0.00716935f $X=6.032 $Y=2.81
+ $X2=6.23 $Y2=2.59
cc_689 N_A_963_115#_c_1246_n N_ECK_c_1350_n 0.00212692f $X=6.11 $Y=1.935
+ $X2=6.23 $Y2=2.59
