magic
tech sky130A
magscale 1 2
timestamp 1606864611
<< checkpaint >>
rect -1209 -1243 2025 2575
<< nwell >>
rect -9 581 837 1341
<< pmos >>
rect 80 617 110 1217
rect 178 617 208 1217
rect 264 617 294 1217
rect 362 617 392 1217
rect 552 617 582 1217
rect 638 617 668 1217
rect 710 617 740 1217
<< nmoslvt >>
rect 80 115 110 315
rect 178 115 208 315
rect 250 115 280 315
rect 442 115 472 315
rect 540 115 570 315
rect 626 115 656 315
rect 712 115 742 315
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 178 315
rect 110 131 133 267
rect 167 131 178 267
rect 110 115 178 131
rect 208 115 250 315
rect 280 267 333 315
rect 280 131 291 267
rect 325 131 333 267
rect 280 115 333 131
rect 389 267 442 315
rect 389 131 397 267
rect 431 131 442 267
rect 389 115 442 131
rect 472 267 540 315
rect 472 131 495 267
rect 529 131 540 267
rect 472 115 540 131
rect 570 267 626 315
rect 570 131 581 267
rect 615 131 626 267
rect 570 115 626 131
rect 656 267 712 315
rect 656 199 667 267
rect 701 199 712 267
rect 656 115 712 199
rect 742 267 795 315
rect 742 131 753 267
rect 787 131 795 267
rect 742 115 795 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 657 35 1201
rect 69 657 80 1201
rect 27 617 80 657
rect 110 1201 178 1217
rect 110 657 133 1201
rect 167 657 178 1201
rect 110 617 178 657
rect 208 1201 264 1217
rect 208 725 219 1201
rect 253 725 264 1201
rect 208 617 264 725
rect 294 1201 362 1217
rect 294 725 305 1201
rect 339 725 362 1201
rect 294 617 362 725
rect 392 1201 445 1217
rect 392 657 403 1201
rect 437 657 445 1201
rect 392 617 445 657
rect 499 1201 552 1217
rect 499 657 507 1201
rect 541 657 552 1201
rect 499 617 552 657
rect 582 1201 638 1217
rect 582 657 593 1201
rect 627 657 638 1201
rect 582 617 638 657
rect 668 617 710 1217
rect 740 1201 796 1217
rect 740 657 751 1201
rect 785 657 796 1201
rect 740 617 796 657
<< ndiffc >>
rect 35 131 69 267
rect 133 131 167 267
rect 291 131 325 267
rect 397 131 431 267
rect 495 131 529 267
rect 581 131 615 267
rect 667 199 701 267
rect 753 131 787 267
<< pdiffc >>
rect 35 657 69 1201
rect 133 657 167 1201
rect 219 725 253 1201
rect 305 725 339 1201
rect 403 657 437 1201
rect 507 657 541 1201
rect 593 657 627 1201
rect 751 657 785 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
rect 707 1271 731 1305
rect 765 1271 789 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
rect 731 1271 765 1305
<< poly >>
rect 80 1217 110 1243
rect 178 1217 208 1243
rect 264 1217 294 1243
rect 362 1217 392 1243
rect 552 1217 582 1243
rect 638 1217 668 1243
rect 710 1217 740 1243
rect 80 403 110 617
rect 178 477 208 617
rect 264 551 294 617
rect 154 461 208 477
rect 154 427 164 461
rect 198 427 208 461
rect 154 411 208 427
rect 43 387 110 403
rect 43 353 53 387
rect 87 353 110 387
rect 43 337 110 353
rect 80 315 110 337
rect 178 315 208 411
rect 250 535 304 551
rect 250 501 260 535
rect 294 501 304 535
rect 250 485 304 501
rect 362 549 392 617
rect 552 549 582 617
rect 362 519 582 549
rect 250 315 280 485
rect 362 424 392 519
rect 638 477 668 617
rect 710 551 740 617
rect 710 535 764 551
rect 710 501 720 535
rect 754 501 764 535
rect 710 485 764 501
rect 338 408 392 424
rect 614 461 668 477
rect 614 427 624 461
rect 658 427 668 461
rect 614 411 668 427
rect 338 374 348 408
rect 382 375 392 408
rect 382 374 570 375
rect 338 345 570 374
rect 442 315 472 345
rect 540 315 570 345
rect 626 315 656 411
rect 712 315 742 485
rect 80 89 110 115
rect 178 89 208 115
rect 250 89 280 115
rect 442 89 472 115
rect 540 89 570 115
rect 626 89 656 115
rect 712 89 742 115
<< polycont >>
rect 164 427 198 461
rect 53 353 87 387
rect 260 501 294 535
rect 720 501 754 535
rect 624 427 658 461
rect 348 374 382 408
<< locali >>
rect 0 1311 836 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 595 1311
rect 629 1271 731 1311
rect 765 1271 836 1311
rect 35 1201 69 1217
rect 35 623 69 649
rect 133 1201 167 1271
rect 133 641 167 657
rect 219 1201 253 1217
rect 219 619 253 725
rect 305 1201 339 1271
rect 305 709 339 725
rect 403 1201 437 1217
rect 219 585 362 619
rect 260 535 294 551
rect 260 485 294 501
rect 148 427 164 461
rect 198 427 214 461
rect 328 424 362 585
rect 403 609 437 657
rect 507 1201 541 1217
rect 403 575 418 609
rect 328 408 382 424
rect 328 392 348 408
rect 37 353 53 387
rect 87 353 110 387
rect 291 374 348 392
rect 291 358 382 374
rect 35 267 69 278
rect 35 115 69 131
rect 133 267 167 283
rect 133 61 167 131
rect 291 267 325 358
rect 418 312 452 575
rect 507 607 541 657
rect 593 1201 627 1271
rect 593 641 627 657
rect 751 1201 785 1217
rect 751 607 785 657
rect 507 573 785 607
rect 507 387 541 573
rect 704 501 720 535
rect 754 501 770 535
rect 608 427 624 461
rect 658 427 674 461
rect 541 353 667 387
rect 291 115 325 131
rect 397 277 452 312
rect 397 267 431 277
rect 397 115 431 131
rect 495 267 529 283
rect 495 61 529 131
rect 581 267 615 283
rect 667 267 701 353
rect 667 183 701 199
rect 753 267 787 283
rect 615 131 753 144
rect 581 110 787 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 836 61
rect 0 0 836 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 595 1305 629 1311
rect 595 1277 629 1305
rect 731 1305 765 1311
rect 731 1277 765 1305
rect 35 657 69 683
rect 35 649 69 657
rect 260 501 294 535
rect 164 427 198 461
rect 418 575 452 609
rect 110 353 144 387
rect 35 278 69 312
rect 720 501 754 535
rect 624 427 658 461
rect 507 353 541 387
rect 667 353 701 387
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
<< metal1 >>
rect 0 1311 836 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 595 1311
rect 629 1277 731 1311
rect 765 1277 836 1311
rect 0 1271 836 1277
rect 23 683 81 689
rect 23 649 35 683
rect 69 649 81 683
rect 23 643 81 649
rect 35 318 69 643
rect 406 609 464 615
rect 406 575 418 609
rect 452 575 486 609
rect 406 569 464 575
rect 248 535 306 541
rect 708 535 766 541
rect 248 501 260 535
rect 294 501 720 535
rect 754 501 766 535
rect 248 500 766 501
rect 248 495 306 500
rect 708 495 766 500
rect 152 462 210 467
rect 612 462 670 467
rect 152 461 670 462
rect 152 427 164 461
rect 198 427 624 461
rect 658 427 670 461
rect 152 421 210 427
rect 612 421 670 427
rect 98 387 156 393
rect 495 387 553 393
rect 655 387 713 393
rect 98 353 110 387
rect 144 353 507 387
rect 541 353 553 387
rect 633 353 667 387
rect 701 353 713 387
rect 98 347 156 353
rect 495 347 553 353
rect 655 347 713 353
rect 23 312 81 318
rect 23 278 35 312
rect 69 278 81 312
rect 23 272 81 278
rect 0 55 836 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 836 55
rect 0 0 836 21
<< labels >>
rlabel metal1 50 477 50 477 1 S
port 1 n
rlabel metal1 737 518 737 518 1 A
port 2 n
rlabel metal1 642 444 642 444 1 B
port 3 n
rlabel metal1 435 592 435 592 1 CO
port 4 n
rlabel metal1 684 370 684 370 1 CON
port 5 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
