magic
tech sky130A
magscale 1 2
timestamp 1612371843
<< nwell >>
rect -9 529 374 1119
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
<< nmoslvt >>
rect 80 115 110 243
rect 152 115 182 243
rect 250 115 280 225
<< ndiff >>
rect 27 228 80 243
rect 27 131 35 228
rect 69 131 80 228
rect 27 115 80 131
rect 110 115 152 243
rect 182 228 235 243
rect 182 131 193 228
rect 227 225 235 228
rect 227 131 250 225
rect 182 115 250 131
rect 280 165 333 225
rect 280 131 291 165
rect 325 131 333 165
rect 280 115 333 131
<< pdiff >>
rect 27 949 80 965
rect 27 745 35 949
rect 69 745 80 949
rect 27 565 80 745
rect 110 949 166 965
rect 110 813 121 949
rect 155 813 166 949
rect 110 565 166 813
rect 196 949 252 965
rect 196 745 207 949
rect 241 745 252 949
rect 196 565 252 745
rect 282 949 335 965
rect 282 677 293 949
rect 327 677 335 949
rect 282 565 335 677
<< ndiffc >>
rect 35 131 69 228
rect 193 131 227 228
rect 291 131 325 165
<< pdiffc >>
rect 35 745 69 949
rect 121 813 155 949
rect 207 745 241 949
rect 293 677 327 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 991
rect 80 528 110 565
rect 44 518 110 528
rect 44 484 60 518
rect 94 484 110 518
rect 44 474 110 484
rect 44 318 74 474
rect 166 432 196 565
rect 252 527 282 565
rect 252 497 309 527
rect 134 416 196 432
rect 134 382 146 416
rect 180 382 196 416
rect 134 366 196 382
rect 44 286 110 318
rect 80 243 110 286
rect 152 243 182 366
rect 279 353 309 497
rect 279 337 333 353
rect 279 319 289 337
rect 250 303 289 319
rect 323 303 333 337
rect 250 287 333 303
rect 250 225 280 287
rect 80 89 110 115
rect 152 89 182 115
rect 250 89 280 115
<< polycont >>
rect 60 484 94 518
rect 146 382 180 416
rect 289 303 323 337
<< locali >>
rect 0 1089 374 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 374 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 797 155 813
rect 207 949 241 965
rect 69 745 207 763
rect 35 729 241 745
rect 293 949 327 965
rect 60 518 94 597
rect 60 468 94 484
rect 128 432 162 523
rect 128 416 180 432
rect 128 382 146 416
rect 128 366 180 382
rect 216 337 250 449
rect 293 409 327 677
rect 216 303 289 337
rect 323 303 339 337
rect 35 228 69 249
rect 35 61 69 131
rect 193 115 227 131
rect 291 165 325 181
rect 291 61 325 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 60 597 94 631
rect 128 523 162 557
rect 216 449 250 483
rect 293 375 327 409
rect 193 228 227 261
rect 193 227 227 228
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 374 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 374 1089
rect 0 1049 374 1055
rect 48 631 106 637
rect 48 597 60 631
rect 94 597 128 631
rect 48 591 106 597
rect 116 557 174 563
rect 116 523 128 557
rect 162 523 196 557
rect 116 517 174 523
rect 204 483 262 489
rect 182 449 216 483
rect 250 449 262 483
rect 204 443 262 449
rect 281 409 339 415
rect 281 375 293 409
rect 327 375 339 409
rect 281 369 339 375
rect 181 261 239 267
rect 293 261 327 369
rect 181 227 193 261
rect 227 227 327 261
rect 181 221 239 227
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel viali 77 614 77 614 1 A0
port 1 n
rlabel viali 233 466 233 466 1 B0
port 2 n
rlabel metal1 310 362 310 362 1 Y
port 3 n
rlabel viali 145 540 145 540 1 A1
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
