* File: sky130_osu_sc_18T_ls__ndlat_l.pxi.spice
* Created: Thu Mar 10 13:45:31 2022
* 
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%GND N_GND_M1001_d N_GND_M1008_d N_GND_M1009_d
+ N_GND_M1001_b N_GND_c_4_p N_GND_c_2_p N_GND_c_15_p N_GND_c_26_p N_GND_c_27_p
+ N_GND_c_70_p GND GND GND GND GND GND PM_SKY130_OSU_SC_18T_LS__NDLAT_L%GND
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%VDD N_VDD_M1005_d N_VDD_M1002_d N_VDD_M1012_d
+ VDD N_VDD_c_107_p N_VDD_c_108_p N_VDD_c_114_p N_VDD_c_124_p N_VDD_c_125_p
+ N_VDD_c_145_p N_VDD_c_154_p VDD VDD VDD VDD
+ PM_SKY130_OSU_SC_18T_LS__NDLAT_L%VDD
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_161_337# N_A_161_337#_M1010_d
+ N_A_161_337#_M1000_d N_A_161_337#_M1001_g N_A_161_337#_M1005_g
+ N_A_161_337#_c_171_n N_A_161_337#_c_173_n N_A_161_337#_c_177_n
+ N_A_161_337#_c_178_n N_A_161_337#_c_179_n N_A_161_337#_c_180_n
+ N_A_161_337#_c_181_n N_A_161_337#_c_192_n N_A_161_337#_c_241_p
+ N_A_161_337#_c_183_n N_A_161_337#_c_221_p N_A_161_337#_c_204_p
+ N_A_161_337#_c_184_n N_A_161_337#_c_194_n
+ PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_161_337#
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%D N_D_M1013_g N_D_M1015_g N_D_c_258_n
+ N_D_c_259_n D PM_SKY130_OSU_SC_18T_LS__NDLAT_L%D
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%CK N_CK_M1000_g N_CK_M1006_g N_CK_c_304_n
+ N_CK_M1003_g N_CK_M1014_g N_CK_c_308_n N_CK_c_309_n N_CK_c_310_n N_CK_c_311_n
+ N_CK_c_314_n N_CK_c_315_n N_CK_c_316_n N_CK_c_317_n N_CK_c_318_n N_CK_c_319_n
+ N_CK_c_320_n N_CK_c_321_n N_CK_c_323_n CK PM_SKY130_OSU_SC_18T_LS__NDLAT_L%CK
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_329_89# N_A_329_89#_M1003_d
+ N_A_329_89#_M1014_d N_A_329_89#_M1010_g N_A_329_89#_c_430_n
+ N_A_329_89#_c_431_n N_A_329_89#_M1004_g N_A_329_89#_c_432_n
+ N_A_329_89#_c_433_n N_A_329_89#_c_434_n N_A_329_89#_c_435_n
+ N_A_329_89#_c_438_n N_A_329_89#_c_439_n N_A_329_89#_c_440_n
+ N_A_329_89#_c_441_n N_A_329_89#_c_442_n N_A_329_89#_c_443_n
+ N_A_329_89#_c_444_n PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_329_89#
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_118_115# N_A_118_115#_M1001_s
+ N_A_118_115#_M1005_s N_A_118_115#_M1008_g N_A_118_115#_M1002_g
+ N_A_118_115#_M1009_g N_A_118_115#_M1012_g N_A_118_115#_c_560_n
+ N_A_118_115#_c_562_n N_A_118_115#_c_563_n N_A_118_115#_c_564_n
+ N_A_118_115#_c_565_n N_A_118_115#_c_583_n N_A_118_115#_c_566_n
+ N_A_118_115#_c_567_n N_A_118_115#_c_588_n N_A_118_115#_c_570_n
+ N_A_118_115#_c_571_n N_A_118_115#_c_572_n N_A_118_115#_c_591_n
+ N_A_118_115#_c_573_n N_A_118_115#_c_574_n N_A_118_115#_c_575_n
+ N_A_118_115#_c_576_n N_A_118_115#_c_577_n
+ PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_118_115#
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%QN N_QN_M1009_s N_QN_M1012_s N_QN_M1011_g
+ N_QN_M1007_g N_QN_c_709_n N_QN_c_710_n N_QN_c_721_n N_QN_c_713_n N_QN_c_715_n
+ N_QN_c_724_n N_QN_c_726_n N_QN_c_716_n QN PM_SKY130_OSU_SC_18T_LS__NDLAT_L%QN
x_PM_SKY130_OSU_SC_18T_LS__NDLAT_L%Q N_Q_M1011_d N_Q_M1007_d N_Q_c_773_n
+ N_Q_c_777_n N_Q_c_778_n N_Q_c_775_n N_Q_c_776_n Q
+ PM_SKY130_OSU_SC_18T_LS__NDLAT_L%Q
cc_1 N_GND_M1001_b N_A_161_337#_c_171_n 0.030793f $X=0.27 $Y=0 $X2=0.94 $Y2=1.85
cc_2 N_GND_c_2_p N_A_161_337#_c_171_n 3.17551e-19 $X=1.145 $Y=0.825 $X2=0.94
+ $Y2=1.85
cc_3 N_GND_M1001_b N_A_161_337#_c_173_n 0.0207466f $X=0.27 $Y=0 $X2=0.94
+ $Y2=1.685
cc_4 N_GND_c_4_p N_A_161_337#_c_173_n 0.00606474f $X=1.06 $Y=0.152 $X2=0.94
+ $Y2=1.685
cc_5 N_GND_c_2_p N_A_161_337#_c_173_n 0.00354579f $X=1.145 $Y=0.825 $X2=0.94
+ $Y2=1.685
cc_6 GND N_A_161_337#_c_173_n 0.00468827f $X=4.43 $Y=0.17 $X2=0.94 $Y2=1.685
cc_7 N_GND_M1001_b N_A_161_337#_c_177_n 0.0417126f $X=0.27 $Y=0 $X2=0.905
+ $Y2=2.805
cc_8 N_GND_M1001_b N_A_161_337#_c_178_n 0.00712311f $X=0.27 $Y=0 $X2=0.905
+ $Y2=2.975
cc_9 N_GND_M1001_b N_A_161_337#_c_179_n 8.14549e-19 $X=0.27 $Y=0 $X2=0.94
+ $Y2=1.935
cc_10 N_GND_M1001_b N_A_161_337#_c_180_n 0.00733729f $X=0.27 $Y=0 $X2=0.94
+ $Y2=3.1
cc_11 N_GND_M1001_b N_A_161_337#_c_181_n 0.00818088f $X=0.27 $Y=0 $X2=1.4
+ $Y2=1.85
cc_12 N_GND_c_2_p N_A_161_337#_c_181_n 0.00816426f $X=1.145 $Y=0.825 $X2=1.4
+ $Y2=1.85
cc_13 N_GND_M1001_b N_A_161_337#_c_183_n 0.00158881f $X=0.27 $Y=0 $X2=1.485
+ $Y2=1.765
cc_14 N_GND_M1001_b N_A_161_337#_c_184_n 0.00313975f $X=0.27 $Y=0 $X2=2.02
+ $Y2=0.825
cc_15 N_GND_c_15_p N_A_161_337#_c_184_n 0.0151591f $X=2.81 $Y=0.152 $X2=2.02
+ $Y2=0.825
cc_16 GND N_A_161_337#_c_184_n 0.00958198f $X=4.43 $Y=0.17 $X2=2.02 $Y2=0.825
cc_17 N_GND_M1001_b N_D_M1013_g 0.040459f $X=0.27 $Y=0 $X2=1.36 $Y2=1.075
cc_18 N_GND_c_2_p N_D_M1013_g 0.00354579f $X=1.145 $Y=0.825 $X2=1.36 $Y2=1.075
cc_19 N_GND_c_15_p N_D_M1013_g 0.00606474f $X=2.81 $Y=0.152 $X2=1.36 $Y2=1.075
cc_20 GND N_D_M1013_g 0.00468827f $X=4.43 $Y=0.17 $X2=1.36 $Y2=1.075
cc_21 N_GND_M1001_b N_D_M1015_g 0.0152798f $X=0.27 $Y=0 $X2=1.36 $Y2=4.585
cc_22 N_GND_M1001_b N_D_c_258_n 0.0294636f $X=0.27 $Y=0 $X2=1.3 $Y2=2.425
cc_23 N_GND_M1001_b N_D_c_259_n 0.00123417f $X=0.27 $Y=0 $X2=1.3 $Y2=2.425
cc_24 N_GND_M1001_b D 0.00683932f $X=0.27 $Y=0 $X2=1.3 $Y2=2.59
cc_25 N_GND_M1001_b N_CK_c_304_n 0.0198314f $X=0.27 $Y=0 $X2=3.11 $Y2=1.665
cc_26 N_GND_c_26_p N_CK_c_304_n 0.00354579f $X=2.895 $Y=0.825 $X2=3.11 $Y2=1.665
cc_27 N_GND_c_27_p N_CK_c_304_n 0.00606474f $X=4.28 $Y=0.152 $X2=3.11 $Y2=1.665
cc_28 GND N_CK_c_304_n 0.00468827f $X=4.43 $Y=0.17 $X2=3.11 $Y2=1.665
cc_29 N_GND_M1001_b N_CK_c_308_n 0.040678f $X=0.27 $Y=0 $X2=3.165 $Y2=2.015
cc_30 N_GND_M1001_b N_CK_c_309_n 0.019996f $X=0.27 $Y=0 $X2=1.78 $Y2=2.765
cc_31 N_GND_M1001_b N_CK_c_310_n 0.0295442f $X=0.27 $Y=0 $X2=2.26 $Y2=1.85
cc_32 N_GND_M1001_b N_CK_c_311_n 0.0175443f $X=0.27 $Y=0 $X2=2.26 $Y2=1.685
cc_33 N_GND_c_15_p N_CK_c_311_n 0.00606474f $X=2.81 $Y=0.152 $X2=2.26 $Y2=1.685
cc_34 GND N_CK_c_311_n 0.00468827f $X=4.43 $Y=0.17 $X2=2.26 $Y2=1.685
cc_35 N_GND_M1001_b N_CK_c_314_n 0.0457025f $X=0.27 $Y=0 $X2=3.137 $Y2=2.78
cc_36 N_GND_M1001_b N_CK_c_315_n 0.0100026f $X=0.27 $Y=0 $X2=3.137 $Y2=2.93
cc_37 N_GND_M1001_b N_CK_c_316_n 0.00696442f $X=0.27 $Y=0 $X2=1.86 $Y2=2.68
cc_38 N_GND_M1001_b N_CK_c_317_n 0.00162414f $X=0.27 $Y=0 $X2=1.945 $Y2=1.85
cc_39 N_GND_M1001_b N_CK_c_318_n 0.00587053f $X=0.27 $Y=0 $X2=2.26 $Y2=1.85
cc_40 N_GND_M1001_b N_CK_c_319_n 6.52287e-19 $X=0.27 $Y=0 $X2=3.245 $Y2=1.85
cc_41 N_GND_M1001_b N_CK_c_320_n 0.00375832f $X=0.27 $Y=0 $X2=1.86 $Y2=2.765
cc_42 N_GND_M1001_b N_CK_c_321_n 0.0180591f $X=0.27 $Y=0 $X2=3.075 $Y2=1.85
cc_43 N_GND_c_26_p N_CK_c_321_n 0.00748954f $X=2.895 $Y=0.825 $X2=3.075 $Y2=1.85
cc_44 N_GND_M1001_b N_CK_c_323_n 0.00401265f $X=0.27 $Y=0 $X2=2.41 $Y2=1.85
cc_45 N_GND_M1001_b N_A_329_89#_M1010_g 0.045859f $X=0.27 $Y=0 $X2=1.72
+ $Y2=1.075
cc_46 N_GND_c_15_p N_A_329_89#_M1010_g 0.00606474f $X=2.81 $Y=0.152 $X2=1.72
+ $Y2=1.075
cc_47 GND N_A_329_89#_M1010_g 0.00468827f $X=4.43 $Y=0.17 $X2=1.72 $Y2=1.075
cc_48 N_GND_M1001_b N_A_329_89#_c_430_n 0.032998f $X=0.27 $Y=0 $X2=2.125 $Y2=2.3
cc_49 N_GND_M1001_b N_A_329_89#_c_431_n 0.00717301f $X=0.27 $Y=0 $X2=1.795
+ $Y2=2.3
cc_50 N_GND_M1001_b N_A_329_89#_c_432_n 0.0203203f $X=0.27 $Y=0 $X2=2.26
+ $Y2=2.765
cc_51 N_GND_M1001_b N_A_329_89#_c_433_n 0.0135787f $X=0.27 $Y=0 $X2=2.26 $Y2=2.6
cc_52 N_GND_M1001_b N_A_329_89#_c_434_n 0.00180771f $X=0.27 $Y=0 $X2=2.26
+ $Y2=2.59
cc_53 N_GND_M1001_b N_A_329_89#_c_435_n 0.00156053f $X=0.27 $Y=0 $X2=3.325
+ $Y2=0.825
cc_54 N_GND_c_27_p N_A_329_89#_c_435_n 0.00754714f $X=4.28 $Y=0.152 $X2=3.325
+ $Y2=0.825
cc_55 GND N_A_329_89#_c_435_n 0.00476261f $X=4.43 $Y=0.17 $X2=3.325 $Y2=0.825
cc_56 N_GND_M1001_b N_A_329_89#_c_438_n 0.0169785f $X=0.27 $Y=0 $X2=3.325
+ $Y2=2.59
cc_57 N_GND_M1001_b N_A_329_89#_c_439_n 0.0150035f $X=0.27 $Y=0 $X2=3.595
+ $Y2=2.185
cc_58 N_GND_M1001_b N_A_329_89#_c_440_n 0.0130615f $X=0.27 $Y=0 $X2=3.595
+ $Y2=1.42
cc_59 N_GND_M1001_b N_A_329_89#_c_441_n 0.0143239f $X=0.27 $Y=0 $X2=3.595
+ $Y2=2.27
cc_60 N_GND_M1001_b N_A_329_89#_c_442_n 0.0175086f $X=0.27 $Y=0 $X2=3.18
+ $Y2=2.59
cc_61 N_GND_M1001_b N_A_329_89#_c_443_n 0.00388969f $X=0.27 $Y=0 $X2=2.405
+ $Y2=2.59
cc_62 N_GND_M1001_b N_A_329_89#_c_444_n 0.00654158f $X=0.27 $Y=0 $X2=3.325
+ $Y2=2.59
cc_63 N_GND_M1001_b N_A_118_115#_M1008_g 0.0343418f $X=0.27 $Y=0 $X2=2.68
+ $Y2=1.075
cc_64 N_GND_c_15_p N_A_118_115#_M1008_g 0.00606474f $X=2.81 $Y=0.152 $X2=2.68
+ $Y2=1.075
cc_65 N_GND_c_26_p N_A_118_115#_M1008_g 0.00354579f $X=2.895 $Y=0.825 $X2=2.68
+ $Y2=1.075
cc_66 GND N_A_118_115#_M1008_g 0.00468827f $X=4.43 $Y=0.17 $X2=2.68 $Y2=1.075
cc_67 N_GND_M1001_b N_A_118_115#_M1002_g 0.0266196f $X=0.27 $Y=0 $X2=2.68
+ $Y2=4.585
cc_68 N_GND_M1001_b N_A_118_115#_M1009_g 0.0332734f $X=0.27 $Y=0 $X2=4.15
+ $Y2=0.945
cc_69 N_GND_c_27_p N_A_118_115#_M1009_g 0.00606474f $X=4.28 $Y=0.152 $X2=4.15
+ $Y2=0.945
cc_70 N_GND_c_70_p N_A_118_115#_M1009_g 0.00388248f $X=4.365 $Y=0.865 $X2=4.15
+ $Y2=0.945
cc_71 GND N_A_118_115#_M1009_g 0.00468827f $X=4.43 $Y=0.17 $X2=4.15 $Y2=0.945
cc_72 N_GND_M1001_b N_A_118_115#_c_560_n 0.030036f $X=0.27 $Y=0 $X2=2.74
+ $Y2=2.22
cc_73 N_GND_c_26_p N_A_118_115#_c_560_n 0.00173465f $X=2.895 $Y=0.825 $X2=2.74
+ $Y2=2.22
cc_74 N_GND_M1001_b N_A_118_115#_c_562_n 0.0313626f $X=0.27 $Y=0 $X2=4.035
+ $Y2=2.22
cc_75 N_GND_M1001_b N_A_118_115#_c_563_n 0.0148769f $X=0.27 $Y=0 $X2=4.037
+ $Y2=2.055
cc_76 N_GND_M1001_b N_A_118_115#_c_564_n 0.0139901f $X=0.27 $Y=0 $X2=4.125
+ $Y2=1.8
cc_77 N_GND_M1001_b N_A_118_115#_c_565_n 0.0348506f $X=0.27 $Y=0 $X2=4.125
+ $Y2=3.855
cc_78 N_GND_M1001_b N_A_118_115#_c_566_n 0.059876f $X=0.27 $Y=0 $X2=0.6 $Y2=2.22
cc_79 N_GND_M1001_b N_A_118_115#_c_567_n 0.00156053f $X=0.27 $Y=0 $X2=0.715
+ $Y2=0.825
cc_80 N_GND_c_4_p N_A_118_115#_c_567_n 0.00757793f $X=1.06 $Y=0.152 $X2=0.715
+ $Y2=0.825
cc_81 GND N_A_118_115#_c_567_n 0.00476261f $X=4.43 $Y=0.17 $X2=0.715 $Y2=0.825
cc_82 N_GND_M1001_b N_A_118_115#_c_570_n 0.00420018f $X=0.27 $Y=0 $X2=2.74
+ $Y2=2.22
cc_83 N_GND_M1001_b N_A_118_115#_c_571_n 0.00383975f $X=0.27 $Y=0 $X2=4.035
+ $Y2=2.22
cc_84 N_GND_M1001_b N_A_118_115#_c_572_n 0.00940876f $X=0.27 $Y=0 $X2=0.715
+ $Y2=1.395
cc_85 N_GND_M1001_b N_A_118_115#_c_573_n 0.0202039f $X=0.27 $Y=0 $X2=3.89
+ $Y2=2.22
cc_86 N_GND_M1001_b N_A_118_115#_c_574_n 0.00259173f $X=0.27 $Y=0 $X2=2.89
+ $Y2=2.22
cc_87 N_GND_M1001_b N_A_118_115#_c_575_n 0.019191f $X=0.27 $Y=0 $X2=0.745
+ $Y2=2.22
cc_88 N_GND_M1001_b N_A_118_115#_c_576_n 0.0218071f $X=0.27 $Y=0 $X2=2.595
+ $Y2=2.22
cc_89 N_GND_M1001_b N_A_118_115#_c_577_n 0.00164722f $X=0.27 $Y=0 $X2=4.035
+ $Y2=2.22
cc_90 N_GND_M1001_b N_QN_M1011_g 0.0613252f $X=0.27 $Y=0 $X2=4.58 $Y2=0.945
cc_91 N_GND_c_70_p N_QN_M1011_g 0.00388248f $X=4.365 $Y=0.865 $X2=4.58 $Y2=0.945
cc_92 GND N_QN_M1011_g 0.00468827f $X=4.43 $Y=0.17 $X2=4.58 $Y2=0.945
cc_93 N_GND_M1001_b N_QN_M1007_g 0.0274779f $X=0.27 $Y=0 $X2=4.58 $Y2=5.085
cc_94 N_GND_M1001_b N_QN_c_709_n 0.0302659f $X=0.27 $Y=0 $X2=4.52 $Y2=2.22
cc_95 N_GND_M1001_b N_QN_c_710_n 0.0107211f $X=0.27 $Y=0 $X2=3.935 $Y2=0.865
cc_96 N_GND_c_27_p N_QN_c_710_n 0.00745733f $X=4.28 $Y=0.152 $X2=3.935 $Y2=0.865
cc_97 GND N_QN_c_710_n 0.00476261f $X=4.43 $Y=0.17 $X2=3.935 $Y2=0.865
cc_98 N_GND_M1001_b N_QN_c_713_n 0.0139291f $X=0.27 $Y=0 $X2=4.435 $Y2=1.85
cc_99 N_GND_c_70_p N_QN_c_713_n 0.00549483f $X=4.365 $Y=0.865 $X2=4.435 $Y2=1.85
cc_100 N_GND_M1001_b N_QN_c_715_n 0.0022353f $X=0.27 $Y=0 $X2=4.02 $Y2=1.85
cc_101 N_GND_M1001_b N_QN_c_716_n 0.00657769f $X=0.27 $Y=0 $X2=4.52 $Y2=2.22
cc_102 N_GND_M1001_b N_Q_c_773_n 0.00913846f $X=0.27 $Y=0 $X2=4.795 $Y2=0.865
cc_103 GND N_Q_c_773_n 0.00476261f $X=4.43 $Y=0.17 $X2=4.795 $Y2=0.865
cc_104 N_GND_M1001_b N_Q_c_775_n 0.0101464f $X=0.27 $Y=0 $X2=4.827 $Y2=1.335
cc_105 N_GND_M1001_b N_Q_c_776_n 0.0738686f $X=0.27 $Y=0 $X2=4.827 $Y2=4.16
cc_106 VDD N_A_161_337#_c_178_n 0.0268222f $X=0.27 $Y=2.905 $X2=0.905 $Y2=2.975
cc_107 N_VDD_c_107_p N_A_161_337#_c_178_n 0.00606474f $X=1.06 $Y=6.507 $X2=0.905
+ $Y2=2.975
cc_108 N_VDD_c_108_p N_A_161_337#_c_178_n 0.00354579f $X=1.145 $Y=3.795
+ $X2=0.905 $Y2=2.975
cc_109 VDD N_A_161_337#_c_178_n 0.00468827f $X=4.425 $Y=6.48 $X2=0.905 $Y2=2.975
cc_110 VDD N_A_161_337#_c_180_n 0.00184258f $X=0.27 $Y=2.905 $X2=0.94 $Y2=3.1
cc_111 N_VDD_M1005_d N_A_161_337#_c_192_n 0.0064093f $X=1.005 $Y=3.085 $X2=1.85
+ $Y2=3.185
cc_112 N_VDD_c_108_p N_A_161_337#_c_192_n 0.00946335f $X=1.145 $Y=3.795 $X2=1.85
+ $Y2=3.185
cc_113 VDD N_A_161_337#_c_194_n 0.00313975f $X=0.27 $Y=2.905 $X2=2.02 $Y2=3.455
cc_114 N_VDD_c_114_p N_A_161_337#_c_194_n 0.0151591f $X=2.81 $Y=6.507 $X2=2.02
+ $Y2=3.455
cc_115 VDD N_A_161_337#_c_194_n 0.00958198f $X=4.425 $Y=6.48 $X2=2.02 $Y2=3.455
cc_116 VDD N_D_M1015_g 0.0197362f $X=0.27 $Y=2.905 $X2=1.36 $Y2=4.585
cc_117 N_VDD_c_108_p N_D_M1015_g 0.00354579f $X=1.145 $Y=3.795 $X2=1.36
+ $Y2=4.585
cc_118 N_VDD_c_114_p N_D_M1015_g 0.00606474f $X=2.81 $Y=6.507 $X2=1.36 $Y2=4.585
cc_119 VDD N_D_M1015_g 0.00468827f $X=4.425 $Y=6.48 $X2=1.36 $Y2=4.585
cc_120 VDD N_CK_M1000_g 0.0201267f $X=0.27 $Y=2.905 $X2=1.72 $Y2=4.585
cc_121 N_VDD_c_114_p N_CK_M1000_g 0.00606474f $X=2.81 $Y=6.507 $X2=1.72
+ $Y2=4.585
cc_122 VDD N_CK_M1000_g 0.00468827f $X=4.425 $Y=6.48 $X2=1.72 $Y2=4.585
cc_123 VDD N_CK_M1014_g 0.0231809f $X=0.27 $Y=2.905 $X2=3.11 $Y2=4.585
cc_124 N_VDD_c_124_p N_CK_M1014_g 0.00354579f $X=2.895 $Y=3.455 $X2=3.11
+ $Y2=4.585
cc_125 N_VDD_c_125_p N_CK_M1014_g 0.00606474f $X=4.28 $Y=6.507 $X2=3.11
+ $Y2=4.585
cc_126 VDD N_CK_M1014_g 0.00468827f $X=4.425 $Y=6.48 $X2=3.11 $Y2=4.585
cc_127 VDD N_CK_c_309_n 0.00444465f $X=0.27 $Y=2.905 $X2=1.78 $Y2=2.765
cc_128 VDD N_CK_c_315_n 0.00461288f $X=0.27 $Y=2.905 $X2=3.137 $Y2=2.93
cc_129 VDD N_A_329_89#_M1004_g 0.020128f $X=0.27 $Y=2.905 $X2=2.32 $Y2=4.585
cc_130 N_VDD_c_114_p N_A_329_89#_M1004_g 0.00606474f $X=2.81 $Y=6.507 $X2=2.32
+ $Y2=4.585
cc_131 VDD N_A_329_89#_M1004_g 0.00468827f $X=4.425 $Y=6.48 $X2=2.32 $Y2=4.585
cc_132 VDD N_A_329_89#_c_432_n 0.00484874f $X=0.27 $Y=2.905 $X2=2.26 $Y2=2.765
cc_133 VDD N_A_329_89#_c_434_n 0.0022456f $X=0.27 $Y=2.905 $X2=2.26 $Y2=2.59
cc_134 VDD N_A_329_89#_c_438_n 0.00685406f $X=0.27 $Y=2.905 $X2=3.325 $Y2=2.59
cc_135 N_VDD_c_125_p N_A_329_89#_c_438_n 0.00754714f $X=4.28 $Y=6.507 $X2=3.325
+ $Y2=2.59
cc_136 VDD N_A_329_89#_c_438_n 0.00476261f $X=4.425 $Y=6.48 $X2=3.325 $Y2=2.59
cc_137 N_VDD_c_124_p N_A_329_89#_c_442_n 0.00634153f $X=2.895 $Y=3.455 $X2=3.18
+ $Y2=2.59
cc_138 VDD N_A_118_115#_M1002_g 0.019758f $X=0.27 $Y=2.905 $X2=2.68 $Y2=4.585
cc_139 N_VDD_c_114_p N_A_118_115#_M1002_g 0.00606474f $X=2.81 $Y=6.507 $X2=2.68
+ $Y2=4.585
cc_140 N_VDD_c_124_p N_A_118_115#_M1002_g 0.00354579f $X=2.895 $Y=3.455 $X2=2.68
+ $Y2=4.585
cc_141 VDD N_A_118_115#_M1002_g 0.00468827f $X=4.425 $Y=6.48 $X2=2.68 $Y2=4.585
cc_142 VDD N_A_118_115#_c_565_n 0.0623258f $X=0.27 $Y=2.905 $X2=4.125 $Y2=3.855
cc_143 VDD N_A_118_115#_c_583_n 0.03391f $X=0.27 $Y=2.905 $X2=4.125 $Y2=4.005
cc_144 N_VDD_c_125_p N_A_118_115#_c_583_n 0.00606474f $X=4.28 $Y=6.507 $X2=4.125
+ $Y2=4.005
cc_145 N_VDD_c_145_p N_A_118_115#_c_583_n 0.00362996f $X=4.365 $Y=4.465
+ $X2=4.125 $Y2=4.005
cc_146 VDD N_A_118_115#_c_583_n 0.00468827f $X=4.425 $Y=6.48 $X2=4.125 $Y2=4.005
cc_147 VDD N_A_118_115#_c_566_n 0.0251549f $X=0.27 $Y=2.905 $X2=0.6 $Y2=2.22
cc_148 VDD N_A_118_115#_c_588_n 0.00156053f $X=0.27 $Y=2.905 $X2=0.715 $Y2=4.135
cc_149 N_VDD_c_107_p N_A_118_115#_c_588_n 0.00757793f $X=1.06 $Y=6.507 $X2=0.715
+ $Y2=4.135
cc_150 VDD N_A_118_115#_c_588_n 0.00476261f $X=4.425 $Y=6.48 $X2=0.715 $Y2=4.135
cc_151 VDD N_A_118_115#_c_591_n 0.0193408f $X=0.27 $Y=2.905 $X2=0.715 $Y2=3.795
cc_152 VDD N_QN_M1007_g 0.07787f $X=0.27 $Y=2.905 $X2=4.58 $Y2=5.085
cc_153 N_VDD_c_145_p N_QN_M1007_g 0.00362996f $X=4.365 $Y=4.465 $X2=4.58
+ $Y2=5.085
cc_154 N_VDD_c_154_p N_QN_M1007_g 0.00606474f $X=4.42 $Y=6.47 $X2=4.58 $Y2=5.085
cc_155 VDD N_QN_M1007_g 0.00468827f $X=4.425 $Y=6.48 $X2=4.58 $Y2=5.085
cc_156 VDD N_QN_c_721_n 0.00659871f $X=0.27 $Y=2.905 $X2=3.935 $Y2=3.96
cc_157 N_VDD_c_125_p N_QN_c_721_n 0.00745733f $X=4.28 $Y=6.507 $X2=3.935
+ $Y2=3.96
cc_158 VDD N_QN_c_721_n 0.00476261f $X=4.425 $Y=6.48 $X2=3.935 $Y2=3.96
cc_159 VDD N_QN_c_724_n 0.0155976f $X=0.27 $Y=2.905 $X2=4.435 $Y2=3.765
cc_160 N_VDD_c_145_p N_QN_c_724_n 0.00816054f $X=4.365 $Y=4.465 $X2=4.435
+ $Y2=3.765
cc_161 VDD N_QN_c_726_n 0.00882478f $X=0.27 $Y=2.905 $X2=4.02 $Y2=3.765
cc_162 VDD N_QN_c_716_n 0.00796734f $X=0.27 $Y=2.905 $X2=4.52 $Y2=2.22
cc_163 VDD QN 0.0168298f $X=0.27 $Y=2.905 $X2=3.94 $Y2=3.96
cc_164 VDD N_Q_c_777_n 0.00648717f $X=0.27 $Y=2.905 $X2=4.795 $Y2=4.33
cc_165 VDD N_Q_c_778_n 0.00156053f $X=0.27 $Y=2.905 $X2=4.795 $Y2=4.465
cc_166 N_VDD_c_154_p N_Q_c_778_n 0.00757793f $X=4.42 $Y=6.47 $X2=4.795 $Y2=4.465
cc_167 VDD N_Q_c_778_n 0.00476261f $X=4.425 $Y=6.48 $X2=4.795 $Y2=4.465
cc_168 VDD N_Q_c_776_n 0.057865f $X=0.27 $Y=2.905 $X2=4.827 $Y2=4.16
cc_169 VDD Q 0.00522778f $X=0.27 $Y=2.905 $X2=4.795 $Y2=4.33
cc_170 N_VDD_c_145_p Q 0.00677841f $X=4.365 $Y=4.465 $X2=4.795 $Y2=4.33
cc_171 N_A_161_337#_c_171_n N_D_M1013_g 0.0207333f $X=0.94 $Y=1.85 $X2=1.36
+ $Y2=1.075
cc_172 N_A_161_337#_c_173_n N_D_M1013_g 0.0196577f $X=0.94 $Y=1.685 $X2=1.36
+ $Y2=1.075
cc_173 N_A_161_337#_c_177_n N_D_M1013_g 0.00885564f $X=0.905 $Y=2.805 $X2=1.36
+ $Y2=1.075
cc_174 N_A_161_337#_c_179_n N_D_M1013_g 2.45848e-19 $X=0.94 $Y=1.935 $X2=1.36
+ $Y2=1.075
cc_175 N_A_161_337#_c_180_n N_D_M1013_g 0.00448652f $X=0.94 $Y=3.1 $X2=1.36
+ $Y2=1.075
cc_176 N_A_161_337#_c_181_n N_D_M1013_g 0.0125105f $X=1.4 $Y=1.85 $X2=1.36
+ $Y2=1.075
cc_177 N_A_161_337#_c_183_n N_D_M1013_g 0.00552645f $X=1.485 $Y=1.765 $X2=1.36
+ $Y2=1.075
cc_178 N_A_161_337#_c_204_p N_D_M1013_g 0.00605553f $X=1.57 $Y=1.43 $X2=1.36
+ $Y2=1.075
cc_179 N_A_161_337#_c_177_n N_D_M1015_g 0.00755439f $X=0.905 $Y=2.805 $X2=1.36
+ $Y2=4.585
cc_180 N_A_161_337#_c_178_n N_D_M1015_g 0.0412319f $X=0.905 $Y=2.975 $X2=1.36
+ $Y2=4.585
cc_181 N_A_161_337#_c_180_n N_D_M1015_g 0.00610289f $X=0.94 $Y=3.1 $X2=1.36
+ $Y2=4.585
cc_182 N_A_161_337#_c_192_n N_D_M1015_g 0.0156361f $X=1.85 $Y=3.185 $X2=1.36
+ $Y2=4.585
cc_183 N_A_161_337#_c_177_n N_D_c_258_n 0.0209207f $X=0.905 $Y=2.805 $X2=1.3
+ $Y2=2.425
cc_184 N_A_161_337#_c_180_n N_D_c_258_n 0.00178864f $X=0.94 $Y=3.1 $X2=1.3
+ $Y2=2.425
cc_185 N_A_161_337#_c_181_n N_D_c_258_n 0.00174867f $X=1.4 $Y=1.85 $X2=1.3
+ $Y2=2.425
cc_186 N_A_161_337#_c_192_n N_D_c_258_n 0.00122128f $X=1.85 $Y=3.185 $X2=1.3
+ $Y2=2.425
cc_187 N_A_161_337#_c_177_n N_D_c_259_n 6.09588e-19 $X=0.905 $Y=2.805 $X2=1.3
+ $Y2=2.425
cc_188 N_A_161_337#_c_180_n N_D_c_259_n 0.0255006f $X=0.94 $Y=3.1 $X2=1.3
+ $Y2=2.425
cc_189 N_A_161_337#_c_181_n N_D_c_259_n 0.00476537f $X=1.4 $Y=1.85 $X2=1.3
+ $Y2=2.425
cc_190 N_A_161_337#_c_192_n N_D_c_259_n 0.00315222f $X=1.85 $Y=3.185 $X2=1.3
+ $Y2=2.425
cc_191 N_A_161_337#_c_180_n D 0.00743369f $X=0.94 $Y=3.1 $X2=1.3 $Y2=2.59
cc_192 N_A_161_337#_c_192_n D 0.0117787f $X=1.85 $Y=3.185 $X2=1.3 $Y2=2.59
cc_193 N_A_161_337#_c_192_n N_CK_M1000_g 0.015571f $X=1.85 $Y=3.185 $X2=1.72
+ $Y2=4.585
cc_194 N_A_161_337#_c_192_n N_CK_c_309_n 0.00158944f $X=1.85 $Y=3.185 $X2=1.78
+ $Y2=2.765
cc_195 N_A_161_337#_c_221_p N_CK_c_310_n 0.00158944f $X=1.85 $Y=1.43 $X2=2.26
+ $Y2=1.85
cc_196 N_A_161_337#_c_181_n N_CK_c_317_n 0.0122336f $X=1.4 $Y=1.85 $X2=1.945
+ $Y2=1.85
cc_197 N_A_161_337#_c_221_p N_CK_c_317_n 0.00917449f $X=1.85 $Y=1.43 $X2=1.945
+ $Y2=1.85
cc_198 N_A_161_337#_c_221_p N_CK_c_318_n 0.0121107f $X=1.85 $Y=1.43 $X2=2.26
+ $Y2=1.85
cc_199 N_A_161_337#_c_180_n N_CK_c_320_n 0.00496637f $X=0.94 $Y=3.1 $X2=1.86
+ $Y2=2.765
cc_200 N_A_161_337#_c_192_n N_CK_c_320_n 0.0153302f $X=1.85 $Y=3.185 $X2=1.86
+ $Y2=2.765
cc_201 N_A_161_337#_c_181_n N_CK_c_323_n 8.68647e-19 $X=1.4 $Y=1.85 $X2=2.41
+ $Y2=1.85
cc_202 N_A_161_337#_c_183_n N_CK_c_323_n 0.00101109f $X=1.485 $Y=1.765 $X2=2.41
+ $Y2=1.85
cc_203 N_A_161_337#_c_221_p N_CK_c_323_n 0.00487841f $X=1.85 $Y=1.43 $X2=2.41
+ $Y2=1.85
cc_204 N_A_161_337#_c_181_n N_A_329_89#_M1010_g 0.00127357f $X=1.4 $Y=1.85
+ $X2=1.72 $Y2=1.075
cc_205 N_A_161_337#_c_183_n N_A_329_89#_M1010_g 0.00554866f $X=1.485 $Y=1.765
+ $X2=1.72 $Y2=1.075
cc_206 N_A_161_337#_c_221_p N_A_329_89#_M1010_g 0.0165456f $X=1.85 $Y=1.43
+ $X2=1.72 $Y2=1.075
cc_207 N_A_161_337#_c_192_n N_A_329_89#_c_432_n 0.0025652f $X=1.85 $Y=3.185
+ $X2=2.26 $Y2=2.765
cc_208 N_A_161_337#_c_192_n N_A_329_89#_c_434_n 0.00103871f $X=1.85 $Y=3.185
+ $X2=2.26 $Y2=2.59
cc_209 N_A_161_337#_c_192_n N_A_329_89#_c_443_n 0.00257262f $X=1.85 $Y=3.185
+ $X2=2.405 $Y2=2.59
cc_210 N_A_161_337#_c_171_n N_A_118_115#_c_566_n 0.0266105f $X=0.94 $Y=1.85
+ $X2=0.6 $Y2=2.22
cc_211 N_A_161_337#_c_173_n N_A_118_115#_c_566_n 0.00700162f $X=0.94 $Y=1.685
+ $X2=0.6 $Y2=2.22
cc_212 N_A_161_337#_c_178_n N_A_118_115#_c_566_n 0.0128109f $X=0.905 $Y=2.975
+ $X2=0.6 $Y2=2.22
cc_213 N_A_161_337#_c_179_n N_A_118_115#_c_566_n 0.0193917f $X=0.94 $Y=1.935
+ $X2=0.6 $Y2=2.22
cc_214 N_A_161_337#_c_180_n N_A_118_115#_c_566_n 0.0810669f $X=0.94 $Y=3.1
+ $X2=0.6 $Y2=2.22
cc_215 N_A_161_337#_c_241_p N_A_118_115#_c_566_n 0.0133619f $X=1.025 $Y=3.185
+ $X2=0.6 $Y2=2.22
cc_216 N_A_161_337#_c_177_n N_A_118_115#_c_575_n 0.0022955f $X=0.905 $Y=2.805
+ $X2=0.745 $Y2=2.22
cc_217 N_A_161_337#_c_180_n N_A_118_115#_c_575_n 0.00271681f $X=0.94 $Y=3.1
+ $X2=0.745 $Y2=2.22
cc_218 N_A_161_337#_c_171_n N_A_118_115#_c_576_n 0.00127165f $X=0.94 $Y=1.85
+ $X2=2.595 $Y2=2.22
cc_219 N_A_161_337#_c_177_n N_A_118_115#_c_576_n 0.00576239f $X=0.905 $Y=2.805
+ $X2=2.595 $Y2=2.22
cc_220 N_A_161_337#_c_180_n N_A_118_115#_c_576_n 0.0226424f $X=0.94 $Y=3.1
+ $X2=2.595 $Y2=2.22
cc_221 N_A_161_337#_c_181_n N_A_118_115#_c_576_n 0.021201f $X=1.4 $Y=1.85
+ $X2=2.595 $Y2=2.22
cc_222 N_A_161_337#_c_221_p N_A_118_115#_c_576_n 0.00611528f $X=1.85 $Y=1.43
+ $X2=2.595 $Y2=2.22
cc_223 N_A_161_337#_c_192_n A_287_617# 0.0060995f $X=1.85 $Y=3.185 $X2=1.435
+ $Y2=3.085
cc_224 N_A_161_337#_c_183_n A_287_115# 6.51949e-19 $X=1.485 $Y=1.765 $X2=1.435
+ $Y2=0.575
cc_225 N_A_161_337#_c_221_p A_287_115# 9.96211e-19 $X=1.85 $Y=1.43 $X2=1.435
+ $Y2=0.575
cc_226 N_A_161_337#_c_204_p A_287_115# 0.0034593f $X=1.57 $Y=1.43 $X2=1.435
+ $Y2=0.575
cc_227 N_D_M1015_g N_CK_c_309_n 0.215574f $X=1.36 $Y=4.585 $X2=1.78 $Y2=2.765
cc_228 N_D_c_259_n N_CK_c_309_n 3.50159e-19 $X=1.3 $Y=2.425 $X2=1.78 $Y2=2.765
cc_229 D N_CK_c_309_n 0.00139761f $X=1.3 $Y=2.59 $X2=1.78 $Y2=2.765
cc_230 N_D_M1013_g N_CK_c_316_n 0.00234107f $X=1.36 $Y=1.075 $X2=1.86 $Y2=2.68
cc_231 N_D_c_258_n N_CK_c_316_n 0.00185841f $X=1.3 $Y=2.425 $X2=1.86 $Y2=2.68
cc_232 N_D_c_259_n N_CK_c_316_n 0.0124483f $X=1.3 $Y=2.425 $X2=1.86 $Y2=2.68
cc_233 D N_CK_c_316_n 0.00606314f $X=1.3 $Y=2.59 $X2=1.86 $Y2=2.68
cc_234 N_D_M1015_g N_CK_c_320_n 0.00165169f $X=1.36 $Y=4.585 $X2=1.86 $Y2=2.765
cc_235 D N_CK_c_320_n 0.00103938f $X=1.3 $Y=2.59 $X2=1.86 $Y2=2.765
cc_236 N_D_M1013_g N_A_329_89#_M1010_g 0.0581908f $X=1.36 $Y=1.075 $X2=1.72
+ $Y2=1.075
cc_237 N_D_c_258_n N_A_329_89#_c_431_n 0.0581908f $X=1.3 $Y=2.425 $X2=1.795
+ $Y2=2.3
cc_238 N_D_c_259_n N_A_329_89#_c_431_n 4.5169e-19 $X=1.3 $Y=2.425 $X2=1.795
+ $Y2=2.3
cc_239 N_D_c_258_n N_A_329_89#_c_433_n 0.00287606f $X=1.3 $Y=2.425 $X2=2.26
+ $Y2=2.6
cc_240 N_D_M1013_g N_A_118_115#_c_576_n 0.00314369f $X=1.36 $Y=1.075 $X2=2.595
+ $Y2=2.22
cc_241 N_D_c_258_n N_A_118_115#_c_576_n 0.00237496f $X=1.3 $Y=2.425 $X2=2.595
+ $Y2=2.22
cc_242 N_D_c_259_n N_A_118_115#_c_576_n 0.00482511f $X=1.3 $Y=2.425 $X2=2.595
+ $Y2=2.22
cc_243 D N_A_118_115#_c_576_n 0.0307072f $X=1.3 $Y=2.59 $X2=2.595 $Y2=2.22
cc_244 N_CK_c_310_n N_A_329_89#_M1010_g 0.0123786f $X=2.26 $Y=1.85 $X2=1.72
+ $Y2=1.075
cc_245 N_CK_c_311_n N_A_329_89#_M1010_g 0.0256778f $X=2.26 $Y=1.685 $X2=1.72
+ $Y2=1.075
cc_246 N_CK_c_316_n N_A_329_89#_M1010_g 0.00936286f $X=1.86 $Y=2.68 $X2=1.72
+ $Y2=1.075
cc_247 N_CK_c_317_n N_A_329_89#_M1010_g 0.00436832f $X=1.945 $Y=1.85 $X2=1.72
+ $Y2=1.075
cc_248 N_CK_c_323_n N_A_329_89#_M1010_g 4.21907e-19 $X=2.41 $Y=1.85 $X2=1.72
+ $Y2=1.075
cc_249 N_CK_c_310_n N_A_329_89#_c_430_n 0.0107061f $X=2.26 $Y=1.85 $X2=2.125
+ $Y2=2.3
cc_250 N_CK_c_316_n N_A_329_89#_c_430_n 0.00994433f $X=1.86 $Y=2.68 $X2=2.125
+ $Y2=2.3
cc_251 N_CK_c_318_n N_A_329_89#_c_430_n 0.00503591f $X=2.26 $Y=1.85 $X2=2.125
+ $Y2=2.3
cc_252 N_CK_c_323_n N_A_329_89#_c_430_n 7.09843e-19 $X=2.41 $Y=1.85 $X2=2.125
+ $Y2=2.3
cc_253 N_CK_c_309_n N_A_329_89#_c_431_n 0.0174061f $X=1.78 $Y=2.765 $X2=1.795
+ $Y2=2.3
cc_254 N_CK_c_316_n N_A_329_89#_c_431_n 0.00254254f $X=1.86 $Y=2.68 $X2=1.795
+ $Y2=2.3
cc_255 N_CK_c_320_n N_A_329_89#_c_431_n 9.11794e-19 $X=1.86 $Y=2.765 $X2=1.795
+ $Y2=2.3
cc_256 N_CK_M1000_g N_A_329_89#_M1004_g 0.0612056f $X=1.72 $Y=4.585 $X2=2.32
+ $Y2=4.585
cc_257 N_CK_c_309_n N_A_329_89#_c_432_n 0.0213338f $X=1.78 $Y=2.765 $X2=2.26
+ $Y2=2.765
cc_258 N_CK_c_310_n N_A_329_89#_c_432_n 0.00224211f $X=2.26 $Y=1.85 $X2=2.26
+ $Y2=2.765
cc_259 N_CK_c_318_n N_A_329_89#_c_432_n 3.82119e-19 $X=2.26 $Y=1.85 $X2=2.26
+ $Y2=2.765
cc_260 N_CK_c_320_n N_A_329_89#_c_432_n 0.00102234f $X=1.86 $Y=2.765 $X2=2.26
+ $Y2=2.765
cc_261 N_CK_c_316_n N_A_329_89#_c_433_n 0.00426729f $X=1.86 $Y=2.68 $X2=2.26
+ $Y2=2.6
cc_262 N_CK_c_309_n N_A_329_89#_c_434_n 8.47686e-19 $X=1.78 $Y=2.765 $X2=2.26
+ $Y2=2.59
cc_263 N_CK_c_310_n N_A_329_89#_c_434_n 8.65047e-19 $X=2.26 $Y=1.85 $X2=2.26
+ $Y2=2.59
cc_264 N_CK_c_316_n N_A_329_89#_c_434_n 0.00783596f $X=1.86 $Y=2.68 $X2=2.26
+ $Y2=2.59
cc_265 N_CK_c_318_n N_A_329_89#_c_434_n 0.00226605f $X=2.26 $Y=1.85 $X2=2.26
+ $Y2=2.59
cc_266 N_CK_c_320_n N_A_329_89#_c_434_n 0.00985033f $X=1.86 $Y=2.765 $X2=2.26
+ $Y2=2.59
cc_267 N_CK_M1014_g N_A_329_89#_c_438_n 0.0103827f $X=3.11 $Y=4.585 $X2=3.325
+ $Y2=2.59
cc_268 N_CK_c_314_n N_A_329_89#_c_438_n 0.0225165f $X=3.137 $Y=2.78 $X2=3.325
+ $Y2=2.59
cc_269 N_CK_c_304_n N_A_329_89#_c_439_n 0.00462924f $X=3.11 $Y=1.665 $X2=3.595
+ $Y2=2.185
cc_270 N_CK_c_308_n N_A_329_89#_c_439_n 0.00395023f $X=3.165 $Y=2.015 $X2=3.595
+ $Y2=2.185
cc_271 N_CK_c_314_n N_A_329_89#_c_439_n 0.00338699f $X=3.137 $Y=2.78 $X2=3.595
+ $Y2=2.185
cc_272 N_CK_c_319_n N_A_329_89#_c_439_n 0.0202148f $X=3.245 $Y=1.85 $X2=3.595
+ $Y2=2.185
cc_273 N_CK_c_321_n N_A_329_89#_c_439_n 0.00788984f $X=3.075 $Y=1.85 $X2=3.595
+ $Y2=2.185
cc_274 N_CK_c_308_n N_A_329_89#_c_440_n 0.00476435f $X=3.165 $Y=2.015 $X2=3.595
+ $Y2=1.42
cc_275 N_CK_c_319_n N_A_329_89#_c_440_n 0.00569038f $X=3.245 $Y=1.85 $X2=3.595
+ $Y2=1.42
cc_276 N_CK_c_321_n N_A_329_89#_c_440_n 0.00408779f $X=3.075 $Y=1.85 $X2=3.595
+ $Y2=1.42
cc_277 N_CK_c_308_n N_A_329_89#_c_441_n 0.00300965f $X=3.165 $Y=2.015 $X2=3.595
+ $Y2=2.27
cc_278 N_CK_c_314_n N_A_329_89#_c_441_n 0.00357453f $X=3.137 $Y=2.78 $X2=3.595
+ $Y2=2.27
cc_279 N_CK_c_319_n N_A_329_89#_c_441_n 0.00584453f $X=3.245 $Y=1.85 $X2=3.595
+ $Y2=2.27
cc_280 N_CK_c_321_n N_A_329_89#_c_441_n 6.56051e-19 $X=3.075 $Y=1.85 $X2=3.595
+ $Y2=2.27
cc_281 N_CK_c_314_n N_A_329_89#_c_442_n 0.00623084f $X=3.137 $Y=2.78 $X2=3.18
+ $Y2=2.59
cc_282 N_CK_c_315_n N_A_329_89#_c_442_n 0.0016292f $X=3.137 $Y=2.93 $X2=3.18
+ $Y2=2.59
cc_283 N_CK_c_316_n N_A_329_89#_c_443_n 0.00742331f $X=1.86 $Y=2.68 $X2=2.405
+ $Y2=2.59
cc_284 N_CK_c_320_n N_A_329_89#_c_443_n 7.22629e-19 $X=1.86 $Y=2.765 $X2=2.405
+ $Y2=2.59
cc_285 N_CK_c_314_n N_A_329_89#_c_444_n 0.00646645f $X=3.137 $Y=2.78 $X2=3.325
+ $Y2=2.59
cc_286 N_CK_c_304_n N_A_118_115#_M1008_g 0.0282002f $X=3.11 $Y=1.665 $X2=2.68
+ $Y2=1.075
cc_287 N_CK_c_308_n N_A_118_115#_M1008_g 0.00979265f $X=3.165 $Y=2.015 $X2=2.68
+ $Y2=1.075
cc_288 N_CK_c_311_n N_A_118_115#_M1008_g 0.096548f $X=2.26 $Y=1.685 $X2=2.68
+ $Y2=1.075
cc_289 N_CK_c_316_n N_A_118_115#_M1008_g 0.00249296f $X=1.86 $Y=2.68 $X2=2.68
+ $Y2=1.075
cc_290 N_CK_c_318_n N_A_118_115#_M1008_g 0.00300048f $X=2.26 $Y=1.85 $X2=2.68
+ $Y2=1.075
cc_291 N_CK_c_319_n N_A_118_115#_M1008_g 0.00230142f $X=3.245 $Y=1.85 $X2=2.68
+ $Y2=1.075
cc_292 N_CK_c_321_n N_A_118_115#_M1008_g 0.0109129f $X=3.075 $Y=1.85 $X2=2.68
+ $Y2=1.075
cc_293 N_CK_c_323_n N_A_118_115#_M1008_g 9.47095e-19 $X=2.41 $Y=1.85 $X2=2.68
+ $Y2=1.075
cc_294 N_CK_c_314_n N_A_118_115#_M1002_g 0.015555f $X=3.137 $Y=2.78 $X2=2.68
+ $Y2=4.585
cc_295 N_CK_c_315_n N_A_118_115#_M1002_g 0.0278012f $X=3.137 $Y=2.93 $X2=2.68
+ $Y2=4.585
cc_296 N_CK_c_314_n N_A_118_115#_c_560_n 0.0211647f $X=3.137 $Y=2.78 $X2=2.74
+ $Y2=2.22
cc_297 N_CK_c_316_n N_A_118_115#_c_560_n 6.23191e-19 $X=1.86 $Y=2.68 $X2=2.74
+ $Y2=2.22
cc_298 N_CK_c_321_n N_A_118_115#_c_560_n 0.00186852f $X=3.075 $Y=1.85 $X2=2.74
+ $Y2=2.22
cc_299 N_CK_c_314_n N_A_118_115#_c_562_n 0.00388214f $X=3.137 $Y=2.78 $X2=4.035
+ $Y2=2.22
cc_300 N_CK_c_308_n N_A_118_115#_c_564_n 0.00464402f $X=3.165 $Y=2.015 $X2=4.125
+ $Y2=1.8
cc_301 N_CK_c_314_n N_A_118_115#_c_570_n 0.0010711f $X=3.137 $Y=2.78 $X2=2.74
+ $Y2=2.22
cc_302 N_CK_c_316_n N_A_118_115#_c_570_n 0.00297176f $X=1.86 $Y=2.68 $X2=2.74
+ $Y2=2.22
cc_303 N_CK_c_321_n N_A_118_115#_c_570_n 0.00451788f $X=3.075 $Y=1.85 $X2=2.74
+ $Y2=2.22
cc_304 N_CK_c_308_n N_A_118_115#_c_573_n 0.00138853f $X=3.165 $Y=2.015 $X2=3.89
+ $Y2=2.22
cc_305 N_CK_c_314_n N_A_118_115#_c_573_n 0.00407354f $X=3.137 $Y=2.78 $X2=3.89
+ $Y2=2.22
cc_306 N_CK_c_319_n N_A_118_115#_c_573_n 0.00262273f $X=3.245 $Y=1.85 $X2=3.89
+ $Y2=2.22
cc_307 N_CK_c_321_n N_A_118_115#_c_573_n 0.0437997f $X=3.075 $Y=1.85 $X2=3.89
+ $Y2=2.22
cc_308 N_CK_c_314_n N_A_118_115#_c_574_n 9.27087e-19 $X=3.137 $Y=2.78 $X2=2.89
+ $Y2=2.22
cc_309 N_CK_c_321_n N_A_118_115#_c_574_n 0.0270759f $X=3.075 $Y=1.85 $X2=2.89
+ $Y2=2.22
cc_310 N_CK_c_309_n N_A_118_115#_c_576_n 7.03361e-19 $X=1.78 $Y=2.765 $X2=2.595
+ $Y2=2.22
cc_311 N_CK_c_310_n N_A_118_115#_c_576_n 0.00155223f $X=2.26 $Y=1.85 $X2=2.595
+ $Y2=2.22
cc_312 N_CK_c_316_n N_A_118_115#_c_576_n 0.0156918f $X=1.86 $Y=2.68 $X2=2.595
+ $Y2=2.22
cc_313 N_CK_c_318_n N_A_118_115#_c_576_n 0.00613294f $X=2.26 $Y=1.85 $X2=2.595
+ $Y2=2.22
cc_314 N_CK_c_320_n N_A_118_115#_c_576_n 0.00531735f $X=1.86 $Y=2.765 $X2=2.595
+ $Y2=2.22
cc_315 N_CK_c_321_n N_A_118_115#_c_576_n 0.0157447f $X=3.075 $Y=1.85 $X2=2.595
+ $Y2=2.22
cc_316 N_CK_c_323_n N_A_118_115#_c_576_n 0.0374821f $X=2.41 $Y=1.85 $X2=2.595
+ $Y2=2.22
cc_317 N_CK_c_304_n N_QN_c_710_n 0.0019799f $X=3.11 $Y=1.665 $X2=3.935 $Y2=0.865
cc_318 N_A_329_89#_c_432_n N_A_118_115#_M1002_g 0.214863f $X=2.26 $Y=2.765
+ $X2=2.68 $Y2=4.585
cc_319 N_A_329_89#_c_433_n N_A_118_115#_M1002_g 0.00761683f $X=2.26 $Y=2.6
+ $X2=2.68 $Y2=4.585
cc_320 N_A_329_89#_c_434_n N_A_118_115#_M1002_g 0.00367682f $X=2.26 $Y=2.59
+ $X2=2.68 $Y2=4.585
cc_321 N_A_329_89#_c_442_n N_A_118_115#_M1002_g 0.0105882f $X=3.18 $Y=2.59
+ $X2=2.68 $Y2=4.585
cc_322 N_A_329_89#_c_443_n N_A_118_115#_M1002_g 8.90723e-19 $X=2.405 $Y=2.59
+ $X2=2.68 $Y2=4.585
cc_323 N_A_329_89#_c_444_n N_A_118_115#_M1002_g 2.82435e-19 $X=3.325 $Y=2.59
+ $X2=2.68 $Y2=4.585
cc_324 N_A_329_89#_c_430_n N_A_118_115#_c_560_n 0.00761683f $X=2.125 $Y=2.3
+ $X2=2.74 $Y2=2.22
cc_325 N_A_329_89#_c_441_n N_A_118_115#_c_560_n 4.25625e-19 $X=3.595 $Y=2.27
+ $X2=2.74 $Y2=2.22
cc_326 N_A_329_89#_c_442_n N_A_118_115#_c_560_n 0.00186852f $X=3.18 $Y=2.59
+ $X2=2.74 $Y2=2.22
cc_327 N_A_329_89#_c_438_n N_A_118_115#_c_562_n 5.07664e-19 $X=3.325 $Y=2.59
+ $X2=4.035 $Y2=2.22
cc_328 N_A_329_89#_c_439_n N_A_118_115#_c_562_n 0.00201953f $X=3.595 $Y=2.185
+ $X2=4.035 $Y2=2.22
cc_329 N_A_329_89#_c_441_n N_A_118_115#_c_562_n 0.00174839f $X=3.595 $Y=2.27
+ $X2=4.035 $Y2=2.22
cc_330 N_A_329_89#_c_439_n N_A_118_115#_c_563_n 0.00266526f $X=3.595 $Y=2.185
+ $X2=4.037 $Y2=2.055
cc_331 N_A_329_89#_c_439_n N_A_118_115#_c_564_n 6.28573e-19 $X=3.595 $Y=2.185
+ $X2=4.125 $Y2=1.8
cc_332 N_A_329_89#_c_438_n N_A_118_115#_c_565_n 0.0279656f $X=3.325 $Y=2.59
+ $X2=4.125 $Y2=3.855
cc_333 N_A_329_89#_c_444_n N_A_118_115#_c_565_n 0.00495161f $X=3.325 $Y=2.59
+ $X2=4.125 $Y2=3.855
cc_334 N_A_329_89#_c_430_n N_A_118_115#_c_570_n 6.64388e-19 $X=2.125 $Y=2.3
+ $X2=2.74 $Y2=2.22
cc_335 N_A_329_89#_c_439_n N_A_118_115#_c_570_n 0.00105677f $X=3.595 $Y=2.185
+ $X2=2.74 $Y2=2.22
cc_336 N_A_329_89#_c_441_n N_A_118_115#_c_570_n 0.0040427f $X=3.595 $Y=2.27
+ $X2=2.74 $Y2=2.22
cc_337 N_A_329_89#_c_442_n N_A_118_115#_c_570_n 0.00487271f $X=3.18 $Y=2.59
+ $X2=2.74 $Y2=2.22
cc_338 N_A_329_89#_c_439_n N_A_118_115#_c_571_n 0.00317568f $X=3.595 $Y=2.185
+ $X2=4.035 $Y2=2.22
cc_339 N_A_329_89#_c_441_n N_A_118_115#_c_571_n 0.00780498f $X=3.595 $Y=2.27
+ $X2=4.035 $Y2=2.22
cc_340 N_A_329_89#_c_438_n N_A_118_115#_c_573_n 2.32884e-19 $X=3.325 $Y=2.59
+ $X2=3.89 $Y2=2.22
cc_341 N_A_329_89#_c_439_n N_A_118_115#_c_573_n 0.0108765f $X=3.595 $Y=2.185
+ $X2=3.89 $Y2=2.22
cc_342 N_A_329_89#_c_441_n N_A_118_115#_c_573_n 0.0224358f $X=3.595 $Y=2.27
+ $X2=3.89 $Y2=2.22
cc_343 N_A_329_89#_c_442_n N_A_118_115#_c_573_n 0.0233839f $X=3.18 $Y=2.59
+ $X2=3.89 $Y2=2.22
cc_344 N_A_329_89#_c_444_n N_A_118_115#_c_573_n 0.0236535f $X=3.325 $Y=2.59
+ $X2=3.89 $Y2=2.22
cc_345 N_A_329_89#_c_430_n N_A_118_115#_c_574_n 4.70316e-19 $X=2.125 $Y=2.3
+ $X2=2.89 $Y2=2.22
cc_346 N_A_329_89#_c_441_n N_A_118_115#_c_574_n 0.00136849f $X=3.595 $Y=2.27
+ $X2=2.89 $Y2=2.22
cc_347 N_A_329_89#_c_442_n N_A_118_115#_c_574_n 0.0270759f $X=3.18 $Y=2.59
+ $X2=2.89 $Y2=2.22
cc_348 N_A_329_89#_M1010_g N_A_118_115#_c_576_n 0.00255623f $X=1.72 $Y=1.075
+ $X2=2.595 $Y2=2.22
cc_349 N_A_329_89#_c_430_n N_A_118_115#_c_576_n 0.00985983f $X=2.125 $Y=2.3
+ $X2=2.595 $Y2=2.22
cc_350 N_A_329_89#_c_431_n N_A_118_115#_c_576_n 0.00164908f $X=1.795 $Y=2.3
+ $X2=2.595 $Y2=2.22
cc_351 N_A_329_89#_c_434_n N_A_118_115#_c_576_n 9.69764e-19 $X=2.26 $Y=2.59
+ $X2=2.595 $Y2=2.22
cc_352 N_A_329_89#_c_442_n N_A_118_115#_c_576_n 0.0147566f $X=3.18 $Y=2.59
+ $X2=2.595 $Y2=2.22
cc_353 N_A_329_89#_c_443_n N_A_118_115#_c_576_n 0.0242903f $X=2.405 $Y=2.59
+ $X2=2.595 $Y2=2.22
cc_354 N_A_329_89#_c_439_n N_A_118_115#_c_577_n 0.00155231f $X=3.595 $Y=2.185
+ $X2=4.035 $Y2=2.22
cc_355 N_A_329_89#_c_441_n N_A_118_115#_c_577_n 0.00170428f $X=3.595 $Y=2.27
+ $X2=4.035 $Y2=2.22
cc_356 N_A_329_89#_c_435_n N_QN_c_710_n 0.0274048f $X=3.325 $Y=0.825 $X2=3.935
+ $Y2=0.865
cc_357 N_A_329_89#_c_439_n N_QN_c_710_n 0.0194424f $X=3.595 $Y=2.185 $X2=3.935
+ $Y2=0.865
cc_358 N_A_329_89#_c_440_n N_QN_c_710_n 0.0136924f $X=3.595 $Y=1.42 $X2=3.935
+ $Y2=0.865
cc_359 N_A_329_89#_c_438_n N_QN_c_721_n 0.0775482f $X=3.325 $Y=2.59 $X2=3.935
+ $Y2=3.96
cc_360 N_A_329_89#_c_439_n N_QN_c_715_n 0.0136585f $X=3.595 $Y=2.185 $X2=4.02
+ $Y2=1.85
cc_361 N_A_329_89#_c_438_n N_QN_c_726_n 0.00707783f $X=3.325 $Y=2.59 $X2=4.02
+ $Y2=3.765
cc_362 N_A_329_89#_c_438_n QN 0.00668284f $X=3.325 $Y=2.59 $X2=3.94 $Y2=3.96
cc_363 N_A_118_115#_M1009_g N_QN_M1011_g 0.0386594f $X=4.15 $Y=0.945 $X2=4.58
+ $Y2=0.945
cc_364 N_A_118_115#_c_563_n N_QN_M1011_g 0.00883234f $X=4.037 $Y=2.055 $X2=4.58
+ $Y2=0.945
cc_365 N_A_118_115#_c_565_n N_QN_M1007_g 0.049185f $X=4.125 $Y=3.855 $X2=4.58
+ $Y2=5.085
cc_366 N_A_118_115#_c_583_n N_QN_M1007_g 0.0240502f $X=4.125 $Y=4.005 $X2=4.58
+ $Y2=5.085
cc_367 N_A_118_115#_c_562_n N_QN_c_709_n 0.0213149f $X=4.035 $Y=2.22 $X2=4.52
+ $Y2=2.22
cc_368 N_A_118_115#_c_571_n N_QN_c_709_n 0.00104076f $X=4.035 $Y=2.22 $X2=4.52
+ $Y2=2.22
cc_369 N_A_118_115#_c_577_n N_QN_c_709_n 9.12123e-19 $X=4.035 $Y=2.22 $X2=4.52
+ $Y2=2.22
cc_370 N_A_118_115#_M1009_g N_QN_c_710_n 0.0196674f $X=4.15 $Y=0.945 $X2=3.935
+ $Y2=0.865
cc_371 N_A_118_115#_c_564_n N_QN_c_710_n 0.00365097f $X=4.125 $Y=1.8 $X2=3.935
+ $Y2=0.865
cc_372 N_A_118_115#_c_565_n N_QN_c_721_n 0.00567875f $X=4.125 $Y=3.855 $X2=3.935
+ $Y2=3.96
cc_373 N_A_118_115#_c_583_n N_QN_c_721_n 0.00746388f $X=4.125 $Y=4.005 $X2=3.935
+ $Y2=3.96
cc_374 N_A_118_115#_c_563_n N_QN_c_713_n 0.00762363f $X=4.037 $Y=2.055 $X2=4.435
+ $Y2=1.85
cc_375 N_A_118_115#_c_564_n N_QN_c_713_n 0.0108917f $X=4.125 $Y=1.8 $X2=4.435
+ $Y2=1.85
cc_376 N_A_118_115#_c_571_n N_QN_c_713_n 0.0093039f $X=4.035 $Y=2.22 $X2=4.435
+ $Y2=1.85
cc_377 N_A_118_115#_c_577_n N_QN_c_713_n 0.0037949f $X=4.035 $Y=2.22 $X2=4.435
+ $Y2=1.85
cc_378 N_A_118_115#_c_562_n N_QN_c_715_n 0.00303508f $X=4.035 $Y=2.22 $X2=4.02
+ $Y2=1.85
cc_379 N_A_118_115#_c_571_n N_QN_c_715_n 0.00899348f $X=4.035 $Y=2.22 $X2=4.02
+ $Y2=1.85
cc_380 N_A_118_115#_c_573_n N_QN_c_715_n 0.0011692f $X=3.89 $Y=2.22 $X2=4.02
+ $Y2=1.85
cc_381 N_A_118_115#_c_577_n N_QN_c_715_n 0.00331526f $X=4.035 $Y=2.22 $X2=4.02
+ $Y2=1.85
cc_382 N_A_118_115#_c_565_n N_QN_c_724_n 0.0195604f $X=4.125 $Y=3.855 $X2=4.435
+ $Y2=3.765
cc_383 N_A_118_115#_c_583_n N_QN_c_724_n 0.00248624f $X=4.125 $Y=4.005 $X2=4.435
+ $Y2=3.765
cc_384 N_A_118_115#_c_562_n N_QN_c_716_n 0.00116148f $X=4.035 $Y=2.22 $X2=4.52
+ $Y2=2.22
cc_385 N_A_118_115#_c_563_n N_QN_c_716_n 0.0022611f $X=4.037 $Y=2.055 $X2=4.52
+ $Y2=2.22
cc_386 N_A_118_115#_c_565_n N_QN_c_716_n 0.0245871f $X=4.125 $Y=3.855 $X2=4.52
+ $Y2=2.22
cc_387 N_A_118_115#_c_571_n N_QN_c_716_n 0.00887114f $X=4.035 $Y=2.22 $X2=4.52
+ $Y2=2.22
cc_388 N_A_118_115#_c_577_n N_QN_c_716_n 0.0035858f $X=4.035 $Y=2.22 $X2=4.52
+ $Y2=2.22
cc_389 N_A_118_115#_c_583_n QN 0.00739895f $X=4.125 $Y=4.005 $X2=3.94 $Y2=3.96
cc_390 N_QN_M1007_g N_Q_c_777_n 0.00360944f $X=4.58 $Y=5.085 $X2=4.795 $Y2=4.33
cc_391 N_QN_M1011_g N_Q_c_775_n 0.00748977f $X=4.58 $Y=0.945 $X2=4.827 $Y2=1.335
cc_392 N_QN_M1011_g N_Q_c_776_n 0.06977f $X=4.58 $Y=0.945 $X2=4.827 $Y2=4.16
cc_393 N_QN_c_713_n N_Q_c_776_n 0.0135849f $X=4.435 $Y=1.85 $X2=4.827 $Y2=4.16
cc_394 N_QN_c_724_n N_Q_c_776_n 0.0135849f $X=4.435 $Y=3.765 $X2=4.827 $Y2=4.16
cc_395 N_QN_c_716_n N_Q_c_776_n 0.124235f $X=4.52 $Y=2.22 $X2=4.827 $Y2=4.16
cc_396 N_QN_M1007_g Q 0.0108355f $X=4.58 $Y=5.085 $X2=4.795 $Y2=4.33
cc_397 N_QN_c_724_n Q 0.00245821f $X=4.435 $Y=3.765 $X2=4.795 $Y2=4.33
