* File: sky130_osu_sc_12T_ms__and2_2.pxi.spice
* Created: Fri Nov 12 15:20:18 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__AND2_2%GND N_GND_M1002_d N_GND_M1007_s N_GND_M1003_b
+ N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p N_GND_c_22_p GND N_GND_c_3_p
+ PM_SKY130_OSU_SC_12T_MS__AND2_2%GND
x_PM_SKY130_OSU_SC_12T_MS__AND2_2%VDD N_VDD_M1001_s N_VDD_M1005_d N_VDD_M1006_d
+ N_VDD_M1001_b N_VDD_c_47_p N_VDD_c_48_p N_VDD_c_59_p N_VDD_c_66_p N_VDD_c_72_p
+ VDD N_VDD_c_49_p PM_SKY130_OSU_SC_12T_MS__AND2_2%VDD
x_PM_SKY130_OSU_SC_12T_MS__AND2_2%A N_A_M1003_g N_A_M1001_g N_A_c_85_n
+ N_A_c_86_n A PM_SKY130_OSU_SC_12T_MS__AND2_2%A
x_PM_SKY130_OSU_SC_12T_MS__AND2_2%B N_B_M1002_g N_B_M1005_g N_B_c_119_n
+ N_B_c_120_n B PM_SKY130_OSU_SC_12T_MS__AND2_2%B
x_PM_SKY130_OSU_SC_12T_MS__AND2_2%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1001_d N_A_27_115#_M1000_g N_A_27_115#_c_176_n
+ N_A_27_115#_M1004_g N_A_27_115#_c_159_n N_A_27_115#_c_160_n
+ N_A_27_115#_M1007_g N_A_27_115#_c_181_n N_A_27_115#_M1006_g
+ N_A_27_115#_c_165_n N_A_27_115#_c_166_n N_A_27_115#_c_167_n
+ N_A_27_115#_c_170_n N_A_27_115#_c_171_n N_A_27_115#_c_187_n
+ N_A_27_115#_c_172_n N_A_27_115#_c_174_n N_A_27_115#_c_175_n
+ N_A_27_115#_c_203_n PM_SKY130_OSU_SC_12T_MS__AND2_2%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__AND2_2%Y N_Y_M1000_d N_Y_M1004_s N_Y_c_242_n
+ N_Y_c_246_n Y N_Y_c_248_n N_Y_c_252_n PM_SKY130_OSU_SC_12T_MS__AND2_2%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.0806078f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1003_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_A_M1003_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=0.835
cc_4 N_GND_M1003_b N_A_c_85_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.285
cc_5 N_GND_M1003_b N_A_c_86_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.285
cc_6 N_GND_M1003_b N_B_M1002_g 0.0460664f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.835
cc_7 N_GND_c_2_p N_B_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.835
cc_8 N_GND_c_8_p N_B_M1002_g 0.00319969f $X=1.05 $Y=0.755 $X2=0.835 $Y2=0.835
cc_9 N_GND_c_3_p N_B_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.835 $Y2=0.835
cc_10 N_GND_M1003_b N_B_M1005_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_11 N_GND_M1003_b N_B_c_119_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.945
cc_12 N_GND_M1003_b N_B_c_120_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.945
cc_13 N_GND_M1003_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.48
cc_14 N_GND_M1003_b N_A_27_115#_M1000_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.835
cc_15 N_GND_c_8_p N_A_27_115#_M1000_g 0.00610843f $X=1.05 $Y=0.755 $X2=1.335
+ $Y2=0.835
cc_16 N_GND_c_16_p N_A_27_115#_M1000_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.835
cc_17 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335
+ $Y2=0.835
cc_18 N_GND_M1003_b N_A_27_115#_c_159_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.33
cc_19 N_GND_M1003_b N_A_27_115#_c_160_n 0.0244031f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.405
cc_20 N_GND_M1003_b N_A_27_115#_M1007_g 0.0264963f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.835
cc_21 N_GND_c_16_p N_A_27_115#_M1007_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.835
cc_22 N_GND_c_22_p N_A_27_115#_M1007_g 0.00502587f $X=1.98 $Y=0.755 $X2=1.765
+ $Y2=0.835
cc_23 N_GND_c_3_p N_A_27_115#_M1007_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765
+ $Y2=0.835
cc_24 N_GND_M1003_b N_A_27_115#_c_165_n 0.00567173f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.405
cc_25 N_GND_M1003_b N_A_27_115#_c_166_n 0.0547984f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_26 N_GND_M1003_b N_A_27_115#_c_167_n 0.0143389f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_27 N_GND_c_2_p N_A_27_115#_c_167_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_28 N_GND_c_3_p N_A_27_115#_c_167_n 0.00476261f $X=1.7 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_29 N_GND_M1003_b N_A_27_115#_c_170_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.455
cc_30 N_GND_M1003_b N_A_27_115#_c_171_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.455
cc_31 N_GND_M1003_b N_A_27_115#_c_172_n 0.0230268f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_32 N_GND_c_8_p N_A_27_115#_c_172_n 0.00704977f $X=1.05 $Y=0.755 $X2=1.43
+ $Y2=1.455
cc_33 N_GND_M1003_b N_A_27_115#_c_174_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.455
cc_34 N_GND_M1003_b N_A_27_115#_c_175_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.065
cc_35 N_GND_M1003_b N_Y_c_242_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_36 N_GND_c_8_p N_Y_c_242_n 0.00806382f $X=1.05 $Y=0.755 $X2=1.55 $Y2=0.755
cc_37 N_GND_c_16_p N_Y_c_242_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_38 N_GND_c_3_p N_Y_c_242_n 0.0047139f $X=1.7 $Y=0.19 $X2=1.55 $Y2=0.755
cc_39 N_GND_M1003_b N_Y_c_246_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_40 N_GND_M1003_b Y 0.0308484f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.74
cc_41 N_GND_M1003_b N_Y_c_248_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1
cc_42 N_GND_c_8_p N_Y_c_248_n 0.00119317f $X=1.05 $Y=0.755 $X2=1.55 $Y2=1
cc_43 N_GND_c_16_p N_Y_c_248_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.55 $Y2=1
cc_44 N_GND_c_22_p N_Y_c_248_n 0.00125659f $X=1.98 $Y=0.755 $X2=1.55 $Y2=1
cc_45 N_GND_M1003_b N_Y_c_252_n 0.0111067f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_46 N_VDD_M1001_b N_A_M1001_g 0.0189471f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_47 N_VDD_c_47_p N_A_M1001_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=3.235
cc_48 N_VDD_c_48_p N_A_M1001_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.235
cc_49 N_VDD_c_49_p N_A_M1001_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.475 $Y2=3.235
cc_50 N_VDD_M1001_b N_A_c_85_n 0.0111025f $X=-0.045 $Y=2.425 $X2=0.475 $Y2=2.285
cc_51 N_VDD_M1001_s N_A_c_86_n 0.0127298f $X=0.135 $Y=2.605 $X2=0.27 $Y2=2.285
cc_52 N_VDD_M1001_b N_A_c_86_n 0.00612103f $X=-0.045 $Y=2.425 $X2=0.27 $Y2=2.285
cc_53 N_VDD_c_47_p N_A_c_86_n 0.00370742f $X=0.26 $Y=3.635 $X2=0.27 $Y2=2.285
cc_54 N_VDD_M1001_s A 0.00742066f $X=0.135 $Y=2.605 $X2=0.275 $Y2=2.85
cc_55 N_VDD_M1001_b A 0.00970321f $X=-0.045 $Y=2.425 $X2=0.275 $Y2=2.85
cc_56 N_VDD_c_47_p A 0.00434783f $X=0.26 $Y=3.635 $X2=0.275 $Y2=2.85
cc_57 N_VDD_M1001_b N_B_M1005_g 0.0187476f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_58 N_VDD_c_48_p N_B_M1005_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.235
cc_59 N_VDD_c_59_p N_B_M1005_g 0.00337744f $X=1.12 $Y=3.295 $X2=0.905 $Y2=3.235
cc_60 N_VDD_c_49_p N_B_M1005_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.905 $Y2=3.235
cc_61 N_VDD_M1001_b N_B_c_120_n 0.00170274f $X=-0.045 $Y=2.425 $X2=0.95
+ $Y2=1.945
cc_62 N_VDD_M1001_b B 0.00856863f $X=-0.045 $Y=2.425 $X2=0.955 $Y2=2.48
cc_63 N_VDD_c_59_p B 0.00240671f $X=1.12 $Y=3.295 $X2=0.955 $Y2=2.48
cc_64 N_VDD_M1001_b N_A_27_115#_c_176_n 0.017104f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.48
cc_65 N_VDD_c_59_p N_A_27_115#_c_176_n 0.00337744f $X=1.12 $Y=3.295 $X2=1.335
+ $Y2=2.48
cc_66 N_VDD_c_66_p N_A_27_115#_c_176_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335
+ $Y2=2.48
cc_67 N_VDD_c_49_p N_A_27_115#_c_176_n 0.00468827f $X=1.7 $Y=4.25 $X2=1.335
+ $Y2=2.48
cc_68 N_VDD_M1001_b N_A_27_115#_c_160_n 0.00813142f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_69 N_VDD_M1001_b N_A_27_115#_c_181_n 0.0212198f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.48
cc_70 N_VDD_c_59_p N_A_27_115#_c_181_n 3.67508e-19 $X=1.12 $Y=3.295 $X2=1.765
+ $Y2=2.48
cc_71 N_VDD_c_66_p N_A_27_115#_c_181_n 0.00610567f $X=1.895 $Y=4.287 $X2=1.765
+ $Y2=2.48
cc_72 N_VDD_c_72_p N_A_27_115#_c_181_n 0.00656078f $X=1.98 $Y=2.955 $X2=1.765
+ $Y2=2.48
cc_73 N_VDD_c_49_p N_A_27_115#_c_181_n 0.00470215f $X=1.7 $Y=4.25 $X2=1.765
+ $Y2=2.48
cc_74 N_VDD_M1001_b N_A_27_115#_c_165_n 0.00216365f $X=-0.045 $Y=2.425 $X2=1.352
+ $Y2=2.405
cc_75 N_VDD_M1001_b N_A_27_115#_c_187_n 0.00155118f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=3.295
cc_76 N_VDD_c_48_p N_A_27_115#_c_187_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69
+ $Y2=3.295
cc_77 N_VDD_c_49_p N_A_27_115#_c_187_n 0.00475776f $X=1.7 $Y=4.25 $X2=0.69
+ $Y2=3.295
cc_78 N_VDD_M1001_b N_A_27_115#_c_175_n 8.22047e-19 $X=-0.045 $Y=2.425 $X2=0.65
+ $Y2=3.065
cc_79 N_VDD_M1001_b N_Y_c_246_n 0.00344954f $X=-0.045 $Y=2.425 $X2=1.55 $Y2=2.11
cc_80 N_VDD_c_66_p N_Y_c_246_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.11
cc_81 N_VDD_c_49_p N_Y_c_246_n 0.00475776f $X=1.7 $Y=4.25 $X2=1.55 $Y2=2.11
cc_82 N_A_M1003_g N_B_M1002_g 0.101204f $X=0.475 $Y=0.835 $X2=0.835 $Y2=0.835
cc_83 N_A_M1003_g N_B_M1005_g 0.048305f $X=0.475 $Y=0.835 $X2=0.905 $Y2=3.235
cc_84 N_A_M1003_g N_B_c_120_n 7.8234e-19 $X=0.475 $Y=0.835 $X2=0.95 $Y2=1.945
cc_85 N_A_M1003_g N_A_27_115#_c_167_n 0.0134114f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.755
cc_86 N_A_M1003_g N_A_27_115#_c_170_n 0.0160984f $X=0.475 $Y=0.835 $X2=0.525
+ $Y2=1.455
cc_87 N_A_c_85_n N_A_27_115#_c_170_n 0.00117122f $X=0.475 $Y=2.285 $X2=0.525
+ $Y2=1.455
cc_88 N_A_c_86_n N_A_27_115#_c_170_n 2.65873e-19 $X=0.27 $Y=2.285 $X2=0.525
+ $Y2=1.455
cc_89 N_A_c_85_n N_A_27_115#_c_171_n 0.00133457f $X=0.475 $Y=2.285 $X2=0.345
+ $Y2=1.455
cc_90 N_A_c_86_n N_A_27_115#_c_171_n 0.0055861f $X=0.27 $Y=2.285 $X2=0.345
+ $Y2=1.455
cc_91 N_A_M1003_g N_A_27_115#_c_174_n 0.00322084f $X=0.475 $Y=0.835 $X2=0.61
+ $Y2=1.455
cc_92 N_A_M1003_g N_A_27_115#_c_175_n 0.0265302f $X=0.475 $Y=0.835 $X2=0.65
+ $Y2=3.065
cc_93 N_A_M1001_g N_A_27_115#_c_175_n 0.0140172f $X=0.475 $Y=3.235 $X2=0.65
+ $Y2=3.065
cc_94 N_A_c_85_n N_A_27_115#_c_175_n 0.00766302f $X=0.475 $Y=2.285 $X2=0.65
+ $Y2=3.065
cc_95 N_A_c_86_n N_A_27_115#_c_175_n 0.0456533f $X=0.27 $Y=2.285 $X2=0.65
+ $Y2=3.065
cc_96 A N_A_27_115#_c_175_n 0.00758489f $X=0.275 $Y=2.85 $X2=0.65 $Y2=3.065
cc_97 N_A_M1001_g N_A_27_115#_c_203_n 0.00865855f $X=0.475 $Y=3.235 $X2=0.65
+ $Y2=3.235
cc_98 N_B_M1002_g N_A_27_115#_M1000_g 0.0271389f $X=0.835 $Y=0.835 $X2=1.335
+ $Y2=0.835
cc_99 N_B_M1005_g N_A_27_115#_c_159_n 0.00773101f $X=0.905 $Y=3.235 $X2=1.37
+ $Y2=2.33
cc_100 N_B_c_119_n N_A_27_115#_c_159_n 0.0206104f $X=0.95 $Y=1.945 $X2=1.37
+ $Y2=2.33
cc_101 N_B_c_120_n N_A_27_115#_c_159_n 0.0033451f $X=0.95 $Y=1.945 $X2=1.37
+ $Y2=2.33
cc_102 N_B_M1005_g N_A_27_115#_c_165_n 0.038666f $X=0.905 $Y=3.235 $X2=1.352
+ $Y2=2.405
cc_103 N_B_c_120_n N_A_27_115#_c_165_n 0.00170598f $X=0.95 $Y=1.945 $X2=1.352
+ $Y2=2.405
cc_104 B N_A_27_115#_c_165_n 0.00386686f $X=0.955 $Y=2.48 $X2=1.352 $Y2=2.405
cc_105 N_B_M1002_g N_A_27_115#_c_166_n 0.0104742f $X=0.835 $Y=0.835 $X2=1.43
+ $Y2=1.455
cc_106 N_B_M1002_g N_A_27_115#_c_172_n 0.0182215f $X=0.835 $Y=0.835 $X2=1.43
+ $Y2=1.455
cc_107 N_B_c_119_n N_A_27_115#_c_172_n 0.00258465f $X=0.95 $Y=1.945 $X2=1.43
+ $Y2=1.455
cc_108 N_B_c_120_n N_A_27_115#_c_172_n 0.0101796f $X=0.95 $Y=1.945 $X2=1.43
+ $Y2=1.455
cc_109 N_B_M1002_g N_A_27_115#_c_175_n 0.00755919f $X=0.835 $Y=0.835 $X2=0.65
+ $Y2=3.065
cc_110 N_B_M1005_g N_A_27_115#_c_175_n 0.0133197f $X=0.905 $Y=3.235 $X2=0.65
+ $Y2=3.065
cc_111 N_B_c_120_n N_A_27_115#_c_175_n 0.0541375f $X=0.95 $Y=1.945 $X2=0.65
+ $Y2=3.065
cc_112 B N_A_27_115#_c_175_n 0.00866797f $X=0.955 $Y=2.48 $X2=0.65 $Y2=3.065
cc_113 B N_A_27_115#_c_203_n 0.00286715f $X=0.955 $Y=2.48 $X2=0.65 $Y2=3.235
cc_114 N_B_c_120_n N_Y_c_246_n 0.0149875f $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_115 B N_Y_c_246_n 0.00649253f $X=0.955 $Y=2.48 $X2=1.55 $Y2=2.11
cc_116 N_B_M1002_g Y 6.71108e-19 $X=0.835 $Y=0.835 $X2=1.555 $Y2=1.74
cc_117 N_B_c_120_n Y 0.00695761f $X=0.95 $Y=1.945 $X2=1.555 $Y2=1.74
cc_118 N_B_M1002_g N_Y_c_248_n 7.71626e-19 $X=0.835 $Y=0.835 $X2=1.55 $Y2=1
cc_119 N_B_c_119_n N_Y_c_252_n 5.70769e-19 $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_120 N_B_c_120_n N_Y_c_252_n 0.00532157f $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_121 N_A_27_115#_M1000_g N_Y_c_242_n 0.00184843f $X=1.335 $Y=0.835 $X2=1.55
+ $Y2=0.755
cc_122 N_A_27_115#_M1007_g N_Y_c_242_n 0.00182852f $X=1.765 $Y=0.835 $X2=1.55
+ $Y2=0.755
cc_123 N_A_27_115#_c_166_n N_Y_c_242_n 0.0016986f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_124 N_A_27_115#_c_172_n N_Y_c_242_n 0.00498892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_125 N_A_27_115#_c_176_n N_Y_c_246_n 0.0026195f $X=1.335 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_126 N_A_27_115#_c_159_n N_Y_c_246_n 0.00744772f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_127 N_A_27_115#_c_160_n N_Y_c_246_n 0.0159823f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_128 N_A_27_115#_c_181_n N_Y_c_246_n 0.00375894f $X=1.765 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_129 N_A_27_115#_c_166_n N_Y_c_246_n 0.0013767f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_130 N_A_27_115#_c_172_n N_Y_c_246_n 0.00273485f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_131 N_A_27_115#_M1000_g Y 0.00251111f $X=1.335 $Y=0.835 $X2=1.555 $Y2=1.74
cc_132 N_A_27_115#_c_159_n Y 0.00892438f $X=1.37 $Y=2.33 $X2=1.555 $Y2=1.74
cc_133 N_A_27_115#_M1007_g Y 0.00251111f $X=1.765 $Y=0.835 $X2=1.555 $Y2=1.74
cc_134 N_A_27_115#_c_166_n Y 0.012094f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_135 N_A_27_115#_c_172_n Y 0.0148238f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_136 N_A_27_115#_M1000_g N_Y_c_248_n 0.00477951f $X=1.335 $Y=0.835 $X2=1.55
+ $Y2=1
cc_137 N_A_27_115#_M1007_g N_Y_c_248_n 0.0084691f $X=1.765 $Y=0.835 $X2=1.55
+ $Y2=1
cc_138 N_A_27_115#_c_172_n N_Y_c_248_n 0.00238892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1
cc_139 N_A_27_115#_c_159_n N_Y_c_252_n 0.00740115f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_140 N_A_27_115#_c_160_n N_Y_c_252_n 0.00229755f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_141 N_A_27_115#_c_166_n N_Y_c_252_n 0.00174847f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_142 N_A_27_115#_c_172_n N_Y_c_252_n 0.00181779f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
