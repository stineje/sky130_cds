* File: sky130_osu_sc_12T_ms__buf_2.pex.spice
* Created: Fri Nov 12 15:21:37 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__BUF_2%GND 1 2 21 23 30 32 40 44 47
r35 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r36 38 40 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.755
r37 33 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r38 32 38 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.305
r39 28 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r40 28 30 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r41 23 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r42 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r43 21 32 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r44 21 33 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r45 21 23 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r46 2 40 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41 $Y=0.575
+ $X2=1.55 $Y2=0.755
r47 1 30 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__BUF_2%VDD 1 2 17 19 25 27 34 40 43
r26 40 43 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r27 34 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r28 32 37 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.55 $Y=4.135 $X2=1.55
+ $Y2=3.635
r29 30 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r30 28 38 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r31 28 30 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r32 27 32 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.465 $Y=4.287
+ $X2=1.55 $Y2=4.135
r33 27 30 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=4.287
+ $X2=1.02 $Y2=4.287
r34 23 38 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r35 23 25 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135 $X2=0.69
+ $Y2=3.635
r36 19 38 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r37 19 21 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r38 17 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r39 17 21 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r40 2 37 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r41 2 34 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r42 1 25 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__BUF_2%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=2.85
+ $X2=0.635 $Y2=2.85
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2 $X2=0.635
+ $Y2=2.85
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635 $Y=2
+ $X2=0.635 $Y2=2
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=2.165
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=1.835
r45 7 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=2.165
r46 3 11 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__BUF_2%A_27_115# 1 3 11 13 15 17 20 22 24 28 33
+ 37 41 45 47 50
r69 46 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.455
+ $X2=0.26 $Y2=1.455
r70 45 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.965 $Y2=1.455
r71 45 46 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.345 $Y2=1.455
r72 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r73 39 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.54 $X2=0.26
+ $Y2=1.455
r74 39 41 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=0.26 $Y=1.54
+ $X2=0.26 $Y2=2.955
r75 35 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.37 $X2=0.26
+ $Y2=1.455
r76 35 37 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r77 32 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.455 $X2=0.965 $Y2=1.455
r78 32 33 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.455
+ $X2=1.18 $Y2=1.455
r79 30 32 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.455
+ $X2=0.965 $Y2=1.455
r80 27 28 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.455
+ $X2=1.335 $Y2=2.455
r81 25 27 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.455
+ $X2=1.18 $Y2=2.455
r82 22 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.53
+ $X2=1.335 $Y2=2.455
r83 22 24 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.335 $Y=2.53
+ $X2=1.335 $Y2=3.235
r84 18 33 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.18 $Y2=1.455
r85 18 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.835
r86 17 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.38
+ $X2=1.18 $Y2=2.455
r87 16 33 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=1.455
r88 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=2.38
r89 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=2.455
r90 13 15 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=3.235
r91 9 30 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=1.455
r92 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=0.835
r93 3 43 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r94 3 41 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r95 1 37 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__BUF_2%Y 1 3 10 16 26 29 32
r40 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=2.48
r41 24 26 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=1.79
r42 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1
r43 23 26 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1.79
r44 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r45 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.48
r46 16 19 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.955
r47 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1 $X2=1.12
+ $Y2=1
r48 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.12 $Y=0.755
+ $X2=1.12 $Y2=1
r49 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r50 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r51 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
.ends

