* File: sky130_osu_sc_18T_hs__tbufi_1.spice
* Created: Fri Nov 12 13:53:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_hs__tbufi_1.pex.spice"
.subckt sky130_osu_sc_18T_hs__tbufi_1  GND VDD OE A Y
* 
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_OE_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1001 A_196_115# N_OE_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g A_196_115# N_GND_M1003_b NLOWVT L=0.15 W=1
+ AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_VDD_M1002_d N_OE_M1002_g N_A_27_115#_M1002_s N_VDD_M1002_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1000 A_196_617# N_A_27_115#_M1000_g N_VDD_M1002_d N_VDD_M1002_b PSHORT L=0.15
+ W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.5 A=0.45 P=6.3 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_196_617# N_VDD_M1002_b PSHORT L=0.15 W=3
+ AD=0.795 AS=0.315 PD=6.53 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=7.296 P=11.44
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__tbufi_1.pxi.spice"
*
.ends
*
*
