* File: sky130_osu_sc_12T_ms__tbufi_1.pex.spice
* Created: Fri Nov 12 15:26:45 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__TBUFI_1%GND 1 17 19 26 35 38
r38 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r39 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r40 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r41 24 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r42 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r43 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r44 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r45 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r46 1 26 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__TBUFI_1%VDD 1 13 15 21 25 29 32
r21 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r22 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r23 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r24 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287 $X2=1.02
+ $Y2=4.287
r25 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r26 19 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.295
r27 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r28 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r29 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r30 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r31 1 21 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__TBUFI_1%OE 2 3 5 6 8 9 11 14 19 22 29 32
c65 29 0 2.60266e-19 $X=0.69 $Y=1.37
r66 26 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.485
+ $X2=0.69 $Y2=1.37
r67 26 32 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=0.69 $Y=1.485
+ $X2=0.69 $Y2=2.365
r68 22 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.37
+ $X2=0.69 $Y2=1.37
r69 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.37 $X2=0.69 $Y2=1.37
r70 12 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.455
+ $X2=0.475 $Y2=2.455
r71 9 19 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.905 $Y=1.17
+ $X2=0.69 $Y2=1.352
r72 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.905 $Y=1.17
+ $X2=0.905 $Y2=0.835
r73 6 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.53
+ $X2=0.475 $Y2=2.455
r74 6 8 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=2.53
+ $X2=0.475 $Y2=3.235
r75 3 19 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.475 $Y=1.17
+ $X2=0.69 $Y2=1.352
r76 3 5 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=1.17
+ $X2=0.475 $Y2=0.835
r77 2 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.38 $X2=0.27
+ $Y2=2.455
r78 1 3 44.3094 $w=2.23e-07 $l=2.69768e-07 $layer=POLY_cond $X=0.27 $Y=1.32
+ $X2=0.475 $Y2=1.17
r79 1 2 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.32 $X2=0.27
+ $Y2=2.38
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__TBUFI_1%A_27_115# 1 3 11 16 20 24 28 30 33
r50 29 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.26
+ $Y2=2
r51 28 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2 $X2=0.8
+ $Y2=2
r52 28 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=2 $X2=0.345
+ $Y2=2
r53 24 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r54 22 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2
r55 22 24 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2.955
r56 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.915
+ $X2=0.26 $Y2=2
r57 18 20 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=0.26 $Y=1.915
+ $X2=0.26 $Y2=0.755
r58 14 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8 $Y=2
+ $X2=0.8 $Y2=2
r59 14 16 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.8 $Y=2 $X2=0.905
+ $Y2=2
r60 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.165
+ $X2=0.905 $Y2=2
r61 9 11 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.905 $Y=2.165
+ $X2=0.905 $Y2=3.235
r62 3 26 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r63 3 24 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r64 1 20 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__TBUFI_1%A 3 7 10 15 20 23
c47 10 0 1.90743e-19 $X=1.325 $Y=1.61
c48 3 0 6.95226e-20 $X=1.265 $Y=0.835
r49 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.61
+ $X2=1.325 $Y2=1.61
r50 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=2.85
+ $X2=1.14 $Y2=2.85
r51 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.695
+ $X2=1.14 $Y2=1.61
r52 13 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=1.695
+ $X2=1.14 $Y2=2.85
r53 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.61 $X2=1.325 $Y2=1.61
r54 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.61
+ $X2=1.325 $Y2=1.775
r55 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.61
+ $X2=1.325 $Y2=1.445
r56 7 12 748.638 $w=1.5e-07 $l=1.46e-06 $layer=POLY_cond $X=1.265 $Y=3.235
+ $X2=1.265 $Y2=1.775
r57 3 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.265 $Y=0.835
+ $X2=1.265 $Y2=1.445
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__TBUFI_1%Y 1 3 10 16 26 29 32
r35 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.995
+ $X2=1.48 $Y2=2.11
r36 24 26 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=1.995
+ $X2=1.48 $Y2=1.34
r37 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.115
+ $X2=1.48 $Y2=1
r38 23 26 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.115
+ $X2=1.48 $Y2=1.34
r39 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.48 $Y=2.955
+ $X2=1.48 $Y2=3.635
r40 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.11
+ $X2=1.48 $Y2=2.11
r41 16 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.48 $Y=2.11
+ $X2=1.48 $Y2=2.955
r42 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1 $X2=1.48
+ $Y2=1
r43 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.48 $Y=0.755
+ $X2=1.48 $Y2=1
r44 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.48 $Y2=3.635
r45 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.48 $Y2=2.955
r46 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.34 $Y=0.575
+ $X2=1.48 $Y2=0.755
.ends

