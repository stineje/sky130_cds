magic
tech sky130A
magscale 1 2
timestamp 1606864613
<< checkpaint >>
rect -1209 -1243 1617 2575
<< nwell >>
rect -9 581 462 1341
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
rect 338 617 368 1217
<< nmoslvt >>
rect 80 115 110 315
rect 152 115 182 315
rect 252 115 282 315
rect 324 115 354 315
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 115 152 315
rect 182 267 252 315
rect 182 131 200 267
rect 234 131 252 267
rect 182 115 252 131
rect 282 115 324 315
rect 354 267 407 315
rect 354 131 365 267
rect 399 131 407 267
rect 354 115 407 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 166 1217
rect 110 861 121 1201
rect 155 861 166 1201
rect 110 617 166 861
rect 196 1201 252 1217
rect 196 793 207 1201
rect 241 793 252 1201
rect 196 617 252 793
rect 282 1133 338 1217
rect 282 793 293 1133
rect 327 793 338 1133
rect 282 617 338 793
rect 368 1201 421 1217
rect 368 793 379 1201
rect 413 793 421 1201
rect 368 617 421 793
<< ndiffc >>
rect 35 131 69 267
rect 200 131 234 267
rect 365 131 399 267
<< pdiffc >>
rect 35 793 69 1201
rect 121 861 155 1201
rect 207 793 241 1201
rect 293 793 327 1133
rect 379 793 413 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 338 1217 368 1243
rect 80 580 110 617
rect 44 570 110 580
rect 44 536 60 570
rect 94 536 110 570
rect 44 526 110 536
rect 44 370 74 526
rect 166 514 196 617
rect 152 484 196 514
rect 116 468 182 484
rect 116 434 128 468
rect 162 434 182 468
rect 116 418 182 434
rect 44 338 110 370
rect 80 315 110 338
rect 152 315 182 418
rect 252 413 282 617
rect 338 478 368 617
rect 338 462 416 478
rect 338 434 370 462
rect 224 397 282 413
rect 224 363 234 397
rect 268 363 282 397
rect 224 347 282 363
rect 252 315 282 347
rect 324 428 370 434
rect 404 428 416 462
rect 324 412 416 428
rect 324 404 368 412
rect 324 315 354 404
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
rect 324 89 354 115
<< polycont >>
rect 60 536 94 570
rect 128 434 162 468
rect 234 363 268 397
rect 370 428 404 462
<< locali >>
rect 0 1311 462 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 462 1311
rect 35 1201 69 1217
rect 121 1201 155 1271
rect 121 845 155 861
rect 207 1201 413 1217
rect 69 793 207 811
rect 241 1183 379 1201
rect 35 777 241 793
rect 293 1133 327 1149
rect 60 570 94 649
rect 293 666 327 793
rect 379 777 413 793
rect 293 632 336 666
rect 60 520 94 536
rect 128 468 162 575
rect 128 418 162 434
rect 216 413 250 501
rect 216 397 268 413
rect 216 363 234 397
rect 234 347 268 363
rect 302 387 336 632
rect 370 462 404 478
rect 370 412 404 428
rect 35 267 69 283
rect 35 61 69 131
rect 200 267 234 279
rect 200 115 234 131
rect 365 267 399 283
rect 365 61 399 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 462 61
rect 0 0 462 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 60 649 94 683
rect 128 575 162 609
rect 216 501 250 535
rect 370 428 404 462
rect 302 353 336 387
rect 200 279 234 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
<< metal1 >>
rect 0 1311 462 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 462 1311
rect 0 1271 462 1277
rect 48 683 106 689
rect 48 649 60 683
rect 94 649 128 683
rect 48 643 106 649
rect 116 609 174 615
rect 116 575 128 609
rect 162 575 196 609
rect 116 569 174 575
rect 204 535 262 541
rect 182 501 216 535
rect 250 501 262 535
rect 204 495 262 501
rect 358 462 416 468
rect 336 428 370 462
rect 404 428 416 462
rect 358 422 416 428
rect 290 387 348 393
rect 290 353 302 387
rect 336 353 348 387
rect 290 347 348 353
rect 188 313 246 319
rect 304 313 338 347
rect 188 279 200 313
rect 234 279 338 313
rect 188 273 246 279
rect 0 55 462 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 462 55
rect 0 0 462 21
<< labels >>
rlabel viali 77 666 77 666 1 A0
port 1 n
rlabel metal1 233 518 233 518 1 B0
port 2 n
rlabel viali 145 592 145 592 1 A1
port 4 n
rlabel viali 387 445 387 445 1 B1
rlabel metal1 321 340 321 340 1 Y
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
