* File: sky130_osu_sc_12T_ms__oai21_l.pxi.spice
* Created: Fri Nov 12 15:25:46 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%GND N_GND_M1003_d N_GND_M1003_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_MS__OAI21_L%GND
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%VDD N_VDD_M1005_d N_VDD_M1001_b N_VDD_c_41_p
+ N_VDD_c_47_p N_VDD_c_53_p VDD N_VDD_c_42_p
+ PM_SKY130_OSU_SC_12T_MS__OAI21_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%A0 N_A0_c_65_n N_A0_M1003_g N_A0_M1001_g
+ N_A0_c_69_n N_A0_c_70_n N_A0_c_71_n N_A0_c_72_n A0
+ PM_SKY130_OSU_SC_12T_MS__OAI21_L%A0
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%A1 N_A1_M1005_g N_A1_M1000_g N_A1_c_107_n
+ N_A1_c_108_n N_A1_c_109_n A1 PM_SKY130_OSU_SC_12T_MS__OAI21_L%A1
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%B0 N_B0_c_160_n N_B0_M1004_g N_B0_M1002_g
+ N_B0_c_164_n N_B0_c_165_n N_B0_c_166_n B0 PM_SKY130_OSU_SC_12T_MS__OAI21_L%B0
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%Y N_Y_M1002_d N_Y_M1001_s N_Y_M1004_d
+ N_Y_c_213_n N_Y_c_216_n N_Y_c_228_n N_Y_c_207_n N_Y_c_219_n N_Y_c_208_n Y
+ N_Y_c_211_n N_Y_c_212_n PM_SKY130_OSU_SC_12T_MS__OAI21_L%Y
x_PM_SKY130_OSU_SC_12T_MS__OAI21_L%A_27_114# N_A_27_114#_M1003_s
+ N_A_27_114#_M1000_d N_A_27_114#_c_261_n N_A_27_114#_c_264_n
+ N_A_27_114#_c_267_n N_A_27_114#_c_268_n
+ PM_SKY130_OSU_SC_12T_MS__OAI21_L%A_27_114#
cc_1 N_GND_M1003_b N_A0_c_65_n 0.0216251f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.215
cc_2 N_GND_c_2_p N_A0_c_65_n 0.00606f $X=0.605 $Y=0.15 $X2=0.475 $Y2=1.215
cc_3 N_GND_c_3_p N_A0_c_65_n 0.00308284f $X=0.69 $Y=0.735 $X2=0.475 $Y2=1.215
cc_4 N_GND_c_4_p N_A0_c_65_n 0.00467791f $X=1.02 $Y=0.185 $X2=0.475 $Y2=1.215
cc_5 N_GND_M1003_b N_A0_c_69_n 0.0245308f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.292
cc_6 N_GND_M1003_b N_A0_c_70_n 0.0342885f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.28
cc_7 N_GND_M1003_b N_A0_c_71_n 0.062092f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.115
cc_8 N_GND_M1003_b N_A0_c_72_n 0.0028102f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.28
cc_9 N_GND_M1003_b N_A1_M1005_g 0.0270518f $X=-0.045 $Y=0 $X2=0.835 $Y2=3.235
cc_10 N_GND_M1003_b N_A1_M1000_g 0.0438085f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.83
cc_11 N_GND_c_3_p N_A1_M1000_g 0.00308284f $X=0.69 $Y=0.735 $X2=0.905 $Y2=0.83
cc_12 N_GND_c_4_p N_A1_M1000_g 0.0046779f $X=1.02 $Y=0.185 $X2=0.905 $Y2=0.83
cc_13 N_GND_M1003_b N_A1_c_107_n 0.0312965f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.74
cc_14 N_GND_M1003_b N_A1_c_108_n 0.00417368f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.74
cc_15 N_GND_M1003_b N_A1_c_109_n 8.57225e-19 $X=-0.045 $Y=0 $X2=0.895 $Y2=2.48
cc_16 N_GND_M1003_b A1 0.00272305f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.48
cc_17 N_GND_M1003_b N_B0_c_160_n 0.0348025f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.665
cc_18 N_GND_M1003_b N_B0_M1004_g 0.049378f $X=-0.045 $Y=0 $X2=1.325 $Y2=3.445
cc_19 N_GND_M1003_b N_B0_M1002_g 0.0371969f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.83
cc_20 N_GND_c_4_p N_B0_M1002_g 0.0046779f $X=1.02 $Y=0.185 $X2=1.335 $Y2=0.83
cc_21 N_GND_M1003_b N_B0_c_164_n 0.00496231f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.11
cc_22 N_GND_M1003_b N_B0_c_165_n 0.00482746f $X=-0.045 $Y=0 $X2=1.285 $Y2=1.5
cc_23 N_GND_M1003_b N_B0_c_166_n 0.00272975f $X=-0.045 $Y=0 $X2=1.395 $Y2=1.5
cc_24 N_GND_M1003_b B0 0.0119375f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.11
cc_25 N_GND_M1003_b N_Y_c_207_n 0.00297509f $X=-0.045 $Y=0 $X2=1.54 $Y2=2.48
cc_26 N_GND_M1003_b N_Y_c_208_n 0.00897794f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.795
cc_27 N_GND_c_4_p N_Y_c_208_n 0.00470726f $X=1.02 $Y=0.185 $X2=1.55 $Y2=0.795
cc_28 N_GND_M1003_b Y 0.00749774f $X=-0.045 $Y=0 $X2=1.54 $Y2=2.48
cc_29 N_GND_M1003_b N_Y_c_211_n 0.0542512f $X=-0.045 $Y=0 $X2=1.542 $Y2=2.365
cc_30 N_GND_M1003_b N_Y_c_212_n 0.0145838f $X=-0.045 $Y=0 $X2=1.55 $Y2=1
cc_31 N_GND_M1003_b N_A_27_114#_c_261_n 0.0015601f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.75
cc_32 N_GND_c_2_p N_A_27_114#_c_261_n 0.00735313f $X=0.605 $Y=0.15 $X2=0.26
+ $Y2=0.75
cc_33 N_GND_c_4_p N_A_27_114#_c_261_n 0.00474759f $X=1.02 $Y=0.185 $X2=0.26
+ $Y2=0.75
cc_34 N_GND_M1003_d N_A_27_114#_c_264_n 0.00176461f $X=0.55 $Y=0.57 $X2=1.035
+ $Y2=1.155
cc_35 N_GND_M1003_b N_A_27_114#_c_264_n 0.0119928f $X=-0.045 $Y=0 $X2=1.035
+ $Y2=1.155
cc_36 N_GND_c_3_p N_A_27_114#_c_264_n 0.0135055f $X=0.69 $Y=0.735 $X2=1.035
+ $Y2=1.155
cc_37 N_GND_M1003_b N_A_27_114#_c_267_n 0.0103371f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.155
cc_38 N_GND_M1003_b N_A_27_114#_c_268_n 0.00888161f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.75
cc_39 N_GND_c_4_p N_A_27_114#_c_268_n 0.00474275f $X=1.02 $Y=0.185 $X2=1.12
+ $Y2=0.75
cc_40 N_VDD_M1001_b N_A0_M1001_g 0.0238089f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_41 N_VDD_c_41_p N_A0_M1001_g 0.00606474f $X=0.965 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_42 N_VDD_c_42_p N_A0_M1001_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.235
cc_43 N_VDD_M1001_b N_A0_c_70_n 0.00574563f $X=-0.045 $Y=2.425 $X2=0.415
+ $Y2=2.28
cc_44 N_VDD_M1001_b N_A0_c_72_n 0.00549657f $X=-0.045 $Y=2.425 $X2=0.415
+ $Y2=2.28
cc_45 N_VDD_M1001_b N_A1_M1005_g 0.0185298f $X=-0.045 $Y=2.425 $X2=0.835
+ $Y2=3.235
cc_46 N_VDD_c_41_p N_A1_M1005_g 0.00606474f $X=0.965 $Y=4.287 $X2=0.835
+ $Y2=3.235
cc_47 N_VDD_c_47_p N_A1_M1005_g 0.00333291f $X=1.05 $Y=3.655 $X2=0.835 $Y2=3.235
cc_48 N_VDD_c_42_p N_A1_M1005_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.835 $Y2=3.235
cc_49 N_VDD_M1001_b N_A1_c_109_n 0.00163533f $X=-0.045 $Y=2.425 $X2=0.895
+ $Y2=2.48
cc_50 N_VDD_M1001_b A1 0.00521027f $X=-0.045 $Y=2.425 $X2=0.895 $Y2=2.48
cc_51 N_VDD_M1001_b N_B0_M1004_g 0.0520054f $X=-0.045 $Y=2.425 $X2=1.325
+ $Y2=3.445
cc_52 N_VDD_c_47_p N_B0_M1004_g 0.00663655f $X=1.05 $Y=3.655 $X2=1.325 $Y2=3.445
cc_53 N_VDD_c_53_p N_B0_M1004_g 0.00606474f $X=1.02 $Y=4.25 $X2=1.325 $Y2=3.445
cc_54 N_VDD_c_42_p N_B0_M1004_g 0.00468827f $X=1.02 $Y=4.25 $X2=1.325 $Y2=3.445
cc_55 N_VDD_M1001_b N_Y_c_213_n 0.00156053f $X=-0.045 $Y=2.425 $X2=0.26 $Y2=3.63
cc_56 N_VDD_c_41_p N_Y_c_213_n 0.00736239f $X=0.965 $Y=4.287 $X2=0.26 $Y2=3.63
cc_57 N_VDD_c_42_p N_Y_c_213_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26 $Y2=3.63
cc_58 N_VDD_M1005_d N_Y_c_216_n 0.00912358f $X=0.91 $Y=2.605 $X2=1.455 $Y2=3.19
cc_59 N_VDD_c_47_p N_Y_c_216_n 0.0135869f $X=1.05 $Y=3.655 $X2=1.455 $Y2=3.19
cc_60 N_VDD_M1001_b N_Y_c_207_n 0.0255776f $X=-0.045 $Y=2.425 $X2=1.54 $Y2=2.48
cc_61 N_VDD_M1001_b N_Y_c_219_n 0.00156053f $X=-0.045 $Y=2.425 $X2=1.54
+ $Y2=3.275
cc_62 N_VDD_c_53_p N_Y_c_219_n 0.00757793f $X=1.02 $Y=4.25 $X2=1.54 $Y2=3.275
cc_63 N_VDD_c_42_p N_Y_c_219_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.54 $Y2=3.275
cc_64 N_VDD_M1001_b Y 0.00957382f $X=-0.045 $Y=2.425 $X2=1.54 $Y2=2.48
cc_65 N_A0_c_70_n N_A1_M1005_g 0.11491f $X=0.415 $Y=2.28 $X2=0.835 $Y2=3.235
cc_66 N_A0_c_71_n N_A1_M1005_g 0.00894734f $X=0.415 $Y=2.115 $X2=0.835 $Y2=3.235
cc_67 N_A0_c_72_n N_A1_M1005_g 0.00413298f $X=0.415 $Y=2.28 $X2=0.835 $Y2=3.235
cc_68 A0 N_A1_M1005_g 0.00376364f $X=0.415 $Y=2.85 $X2=0.835 $Y2=3.235
cc_69 N_A0_c_65_n N_A1_M1000_g 0.0249708f $X=0.475 $Y=1.215 $X2=0.905 $Y2=0.83
cc_70 N_A0_c_71_n N_A1_M1000_g 0.00763255f $X=0.415 $Y=2.115 $X2=0.905 $Y2=0.83
cc_71 N_A0_c_71_n N_A1_c_107_n 0.014675f $X=0.415 $Y=2.115 $X2=0.845 $Y2=1.74
cc_72 N_A0_c_70_n N_A1_c_108_n 8.44103e-19 $X=0.415 $Y=2.28 $X2=0.845 $Y2=1.74
cc_73 N_A0_c_71_n N_A1_c_108_n 0.00346793f $X=0.415 $Y=2.115 $X2=0.845 $Y2=1.74
cc_74 N_A0_c_72_n N_A1_c_108_n 0.0189532f $X=0.415 $Y=2.28 $X2=0.845 $Y2=1.74
cc_75 N_A0_M1001_g N_A1_c_109_n 8.44103e-19 $X=0.475 $Y=3.235 $X2=0.895 $Y2=2.48
cc_76 N_A0_c_70_n A1 0.00357623f $X=0.415 $Y=2.28 $X2=0.895 $Y2=2.48
cc_77 N_A0_c_72_n A1 0.00685942f $X=0.415 $Y=2.28 $X2=0.895 $Y2=2.48
cc_78 N_A0_c_72_n N_Y_M1001_s 0.00842425f $X=0.415 $Y=2.28 $X2=0.135 $Y2=2.605
cc_79 A0 N_Y_M1001_s 0.0119025f $X=0.415 $Y=2.85 $X2=0.135 $Y2=2.605
cc_80 N_A0_M1001_g N_Y_c_216_n 0.0157489f $X=0.475 $Y=3.235 $X2=1.455 $Y2=3.19
cc_81 N_A0_c_72_n N_Y_c_216_n 0.0069936f $X=0.415 $Y=2.28 $X2=1.455 $Y2=3.19
cc_82 A0 N_Y_c_216_n 0.0116431f $X=0.415 $Y=2.85 $X2=1.455 $Y2=3.19
cc_83 N_A0_c_70_n N_Y_c_228_n 0.00152768f $X=0.415 $Y=2.28 $X2=0.345 $Y2=3.19
cc_84 N_A0_c_72_n N_Y_c_228_n 9.01113e-19 $X=0.415 $Y=2.28 $X2=0.345 $Y2=3.19
cc_85 A0 N_Y_c_228_n 0.00385855f $X=0.415 $Y=2.85 $X2=0.345 $Y2=3.19
cc_86 A0 A_110_521# 0.0100173f $X=0.415 $Y=2.85 $X2=0.55 $Y2=2.605
cc_87 N_A0_c_65_n N_A_27_114#_c_264_n 0.0127824f $X=0.475 $Y=1.215 $X2=1.035
+ $Y2=1.155
cc_88 N_A0_c_69_n N_A_27_114#_c_264_n 0.00996929f $X=0.475 $Y=1.292 $X2=1.035
+ $Y2=1.155
cc_89 N_A0_c_69_n N_A_27_114#_c_267_n 0.00538489f $X=0.475 $Y=1.292 $X2=0.345
+ $Y2=1.155
cc_90 N_A1_M1000_g N_B0_c_160_n 8.29743e-19 $X=0.905 $Y=0.83 $X2=1.325 $Y2=1.665
cc_91 N_A1_c_107_n N_B0_c_160_n 0.0140152f $X=0.845 $Y=1.74 $X2=1.325 $Y2=1.665
cc_92 N_A1_c_108_n N_B0_c_160_n 2.71846e-19 $X=0.845 $Y=1.74 $X2=1.325 $Y2=1.665
cc_93 N_A1_M1005_g N_B0_M1004_g 0.0652523f $X=0.835 $Y=3.235 $X2=1.325 $Y2=3.445
cc_94 N_A1_c_108_n N_B0_M1004_g 0.00417871f $X=0.845 $Y=1.74 $X2=1.325 $Y2=3.445
cc_95 N_A1_c_109_n N_B0_M1004_g 0.00113925f $X=0.895 $Y=2.48 $X2=1.325 $Y2=3.445
cc_96 A1 N_B0_M1004_g 0.00127778f $X=0.895 $Y=2.48 $X2=1.325 $Y2=3.445
cc_97 N_A1_M1000_g N_B0_M1002_g 0.0328293f $X=0.905 $Y=0.83 $X2=1.335 $Y2=0.83
cc_98 N_A1_M1005_g N_B0_c_164_n 9.28322e-19 $X=0.835 $Y=3.235 $X2=1.2 $Y2=2.11
cc_99 N_A1_c_107_n N_B0_c_164_n 0.00180004f $X=0.845 $Y=1.74 $X2=1.2 $Y2=2.11
cc_100 N_A1_c_108_n N_B0_c_164_n 0.0387326f $X=0.845 $Y=1.74 $X2=1.2 $Y2=2.11
cc_101 A1 N_B0_c_164_n 2.28089e-19 $X=0.895 $Y=2.48 $X2=1.2 $Y2=2.11
cc_102 N_A1_M1000_g N_B0_c_165_n 0.00424671f $X=0.905 $Y=0.83 $X2=1.285 $Y2=1.5
cc_103 N_A1_c_108_n N_B0_c_165_n 7.09995e-19 $X=0.845 $Y=1.74 $X2=1.285 $Y2=1.5
cc_104 N_A1_c_107_n B0 0.00173697f $X=0.845 $Y=1.74 $X2=1.2 $Y2=2.11
cc_105 N_A1_c_108_n B0 0.008632f $X=0.845 $Y=1.74 $X2=1.2 $Y2=2.11
cc_106 N_A1_c_109_n B0 2.4196e-19 $X=0.895 $Y=2.48 $X2=1.2 $Y2=2.11
cc_107 A1 B0 0.0191116f $X=0.895 $Y=2.48 $X2=1.2 $Y2=2.11
cc_108 N_A1_M1005_g N_Y_c_216_n 0.0165071f $X=0.835 $Y=3.235 $X2=1.455 $Y2=3.19
cc_109 N_A1_c_109_n N_Y_c_216_n 0.00294448f $X=0.895 $Y=2.48 $X2=1.455 $Y2=3.19
cc_110 A1 N_Y_c_216_n 0.0102328f $X=0.895 $Y=2.48 $X2=1.455 $Y2=3.19
cc_111 N_A1_c_109_n N_Y_c_207_n 0.00408285f $X=0.895 $Y=2.48 $X2=1.54 $Y2=2.48
cc_112 A1 N_Y_c_207_n 9.93956e-19 $X=0.895 $Y=2.48 $X2=1.54 $Y2=2.48
cc_113 N_A1_c_109_n Y 5.19115e-19 $X=0.895 $Y=2.48 $X2=1.54 $Y2=2.48
cc_114 A1 Y 0.0182426f $X=0.895 $Y=2.48 $X2=1.54 $Y2=2.48
cc_115 N_A1_M1000_g N_Y_c_211_n 3.23152e-19 $X=0.905 $Y=0.83 $X2=1.542 $Y2=2.365
cc_116 N_A1_c_108_n N_Y_c_211_n 0.00507182f $X=0.845 $Y=1.74 $X2=1.542 $Y2=2.365
cc_117 N_A1_M1000_g N_A_27_114#_c_264_n 0.0163899f $X=0.905 $Y=0.83 $X2=1.035
+ $Y2=1.155
cc_118 N_A1_c_107_n N_A_27_114#_c_264_n 0.00370477f $X=0.845 $Y=1.74 $X2=1.035
+ $Y2=1.155
cc_119 N_A1_c_108_n N_A_27_114#_c_264_n 0.00800525f $X=0.845 $Y=1.74 $X2=1.035
+ $Y2=1.155
cc_120 N_B0_M1004_g N_Y_c_216_n 0.0176498f $X=1.325 $Y=3.445 $X2=1.455 $Y2=3.19
cc_121 N_B0_M1004_g N_Y_c_207_n 0.022499f $X=1.325 $Y=3.445 $X2=1.54 $Y2=2.48
cc_122 N_B0_c_160_n N_Y_c_208_n 0.0011207f $X=1.325 $Y=1.665 $X2=1.55 $Y2=0.795
cc_123 N_B0_M1002_g N_Y_c_208_n 0.00248617f $X=1.335 $Y=0.83 $X2=1.55 $Y2=0.795
cc_124 N_B0_c_166_n N_Y_c_208_n 0.00310915f $X=1.395 $Y=1.5 $X2=1.55 $Y2=0.795
cc_125 N_B0_M1004_g Y 0.0043049f $X=1.325 $Y=3.445 $X2=1.54 $Y2=2.48
cc_126 N_B0_c_160_n N_Y_c_211_n 0.00499921f $X=1.325 $Y=1.665 $X2=1.542
+ $Y2=2.365
cc_127 N_B0_M1004_g N_Y_c_211_n 0.0134421f $X=1.325 $Y=3.445 $X2=1.542 $Y2=2.365
cc_128 N_B0_M1002_g N_Y_c_211_n 0.0048469f $X=1.335 $Y=0.83 $X2=1.542 $Y2=2.365
cc_129 N_B0_c_164_n N_Y_c_211_n 0.0190824f $X=1.2 $Y=2.11 $X2=1.542 $Y2=2.365
cc_130 N_B0_c_166_n N_Y_c_211_n 0.0128496f $X=1.395 $Y=1.5 $X2=1.542 $Y2=2.365
cc_131 B0 N_Y_c_211_n 0.0235926f $X=1.2 $Y=2.11 $X2=1.542 $Y2=2.365
cc_132 N_B0_c_160_n N_Y_c_212_n 0.00189554f $X=1.325 $Y=1.665 $X2=1.55 $Y2=1
cc_133 N_B0_M1002_g N_Y_c_212_n 0.003655f $X=1.335 $Y=0.83 $X2=1.55 $Y2=1
cc_134 N_B0_c_166_n N_Y_c_212_n 0.0028145f $X=1.395 $Y=1.5 $X2=1.55 $Y2=1
cc_135 N_B0_M1002_g N_A_27_114#_c_264_n 0.00480345f $X=1.335 $Y=0.83 $X2=1.035
+ $Y2=1.155
cc_136 N_B0_c_165_n N_A_27_114#_c_264_n 0.00825083f $X=1.285 $Y=1.5 $X2=1.035
+ $Y2=1.155
cc_137 N_Y_c_216_n A_110_521# 0.00573878f $X=1.455 $Y=3.19 $X2=0.55 $Y2=2.605
cc_138 N_Y_c_211_n N_A_27_114#_c_264_n 0.00568156f $X=1.542 $Y=2.365 $X2=1.035
+ $Y2=1.155
cc_139 N_Y_c_212_n N_A_27_114#_c_264_n 0.00216548f $X=1.55 $Y=1 $X2=1.035
+ $Y2=1.155
cc_140 N_Y_c_212_n N_A_27_114#_c_268_n 0.0046453f $X=1.55 $Y=1 $X2=1.12 $Y2=0.75
