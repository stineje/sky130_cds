* File: sky130_osu_sc_15T_ls__aoi21_l.pxi.spice
* Created: Fri Nov 12 14:54:25 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%GND N_GND_M1003_s N_GND_M1005_d N_GND_M1003_b
+ N_GND_c_3_p N_GND_c_4_p N_GND_c_20_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_15T_LS__AOI21_L%GND
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%VDD N_VDD_M1000_d N_VDD_M1000_b N_VDD_c_43_p
+ N_VDD_c_44_p N_VDD_c_50_p VDD N_VDD_c_45_p
+ PM_SKY130_OSU_SC_15T_LS__AOI21_L%VDD
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%A0 N_A0_c_68_n N_A0_c_69_n N_A0_M1003_g
+ N_A0_M1000_g N_A0_c_73_n N_A0_c_75_n N_A0_c_76_n A0
+ PM_SKY130_OSU_SC_15T_LS__AOI21_L%A0
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%A1 N_A1_M1002_g N_A1_M1004_g N_A1_c_109_n
+ N_A1_c_110_n N_A1_c_111_n A1 PM_SKY130_OSU_SC_15T_LS__AOI21_L%A1
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%B0 N_B0_M1005_g N_B0_M1001_g N_B0_c_160_n
+ N_B0_c_161_n N_B0_c_162_n N_B0_c_164_n N_B0_c_165_n N_B0_c_166_n B0
+ PM_SKY130_OSU_SC_15T_LS__AOI21_L%B0
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%A_27_565# N_A_27_565#_M1000_s
+ N_A_27_565#_M1004_d N_A_27_565#_c_209_n N_A_27_565#_c_212_n
+ N_A_27_565#_c_222_n N_A_27_565#_c_214_n
+ PM_SKY130_OSU_SC_15T_LS__AOI21_L%A_27_565#
x_PM_SKY130_OSU_SC_15T_LS__AOI21_L%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_225_n
+ N_Y_c_228_n N_Y_c_229_n N_Y_c_231_n Y N_Y_c_234_n
+ PM_SKY130_OSU_SC_15T_LS__AOI21_L%Y
cc_1 N_GND_M1003_b N_A0_c_68_n 0.0660236f $X=-0.045 $Y=0 $X2=0.295 $Y2=2.37
cc_2 N_GND_M1003_b N_A0_c_69_n 0.0198745f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.43
cc_3 N_GND_c_3_p N_A0_c_69_n 0.00502587f $X=0.26 $Y=0.74 $X2=0.475 $Y2=1.43
cc_4 N_GND_c_4_p N_A0_c_69_n 0.00606474f $X=1.455 $Y=0.152 $X2=0.475 $Y2=1.43
cc_5 N_GND_c_5_p N_A0_c_69_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.43
cc_6 N_GND_M1003_b N_A0_c_73_n 0.0322892f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.51
cc_7 N_GND_c_3_p N_A0_c_73_n 0.00587964f $X=0.26 $Y=0.74 $X2=0.475 $Y2=1.51
cc_8 N_GND_M1003_b N_A0_c_75_n 0.0421132f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.505
cc_9 N_GND_M1003_b N_A0_c_76_n 0.00438599f $X=-0.045 $Y=0 $X2=0.385 $Y2=2.505
cc_10 N_GND_M1003_b N_A1_M1002_g 0.0407759f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_11 N_GND_c_4_p N_A1_M1002_g 0.00606474f $X=1.455 $Y=0.152 $X2=0.835 $Y2=0.945
cc_12 N_GND_c_5_p N_A1_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.945
cc_13 N_GND_M1003_b N_A1_M1004_g 0.0273376f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_14 N_GND_M1003_b N_A1_c_109_n 0.0355308f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.995
cc_15 N_GND_M1003_b N_A1_c_110_n 0.00889603f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.7
cc_16 N_GND_M1003_b N_A1_c_111_n 0.00478352f $X=-0.045 $Y=0 $X2=0.815 $Y2=1.995
cc_17 N_GND_M1003_b A1 0.00323672f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.7
cc_18 N_GND_M1003_b N_B0_M1005_g 0.0350932f $X=-0.045 $Y=0 $X2=1.325 $Y2=0.835
cc_19 N_GND_c_4_p N_B0_M1005_g 0.00606474f $X=1.455 $Y=0.152 $X2=1.325 $Y2=0.835
cc_20 N_GND_c_20_p N_B0_M1005_g 0.00502587f $X=1.54 $Y=0.74 $X2=1.325 $Y2=0.835
cc_21 N_GND_c_5_p N_B0_M1005_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.325 $Y2=0.835
cc_22 N_GND_M1003_b N_B0_M1001_g 5.06723e-19 $X=-0.045 $Y=0 $X2=1.335 $Y2=3.825
cc_23 N_GND_M1003_b N_B0_c_160_n 0.0493362f $X=-0.045 $Y=0 $X2=1.47 $Y2=2.485
cc_24 N_GND_M1003_b N_B0_c_161_n 0.0237317f $X=-0.045 $Y=0 $X2=1.47 $Y2=2.56
cc_25 N_GND_M1003_b N_B0_c_162_n 0.0498038f $X=-0.045 $Y=0 $X2=1.47 $Y2=1.6
cc_26 N_GND_c_20_p N_B0_c_162_n 0.0022951f $X=1.54 $Y=0.74 $X2=1.47 $Y2=1.6
cc_27 N_GND_M1003_b N_B0_c_164_n 0.0141127f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.33
cc_28 N_GND_M1003_b N_B0_c_165_n 0.00387834f $X=-0.045 $Y=0 $X2=1.25 $Y2=1.6
cc_29 N_GND_M1003_b N_B0_c_166_n 0.011995f $X=-0.045 $Y=0 $X2=1.53 $Y2=1.6
cc_30 N_GND_c_20_p N_B0_c_166_n 0.00200373f $X=1.54 $Y=0.74 $X2=1.53 $Y2=1.6
cc_31 N_GND_M1003_b B0 0.0176529f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.33
cc_32 N_GND_M1003_b N_Y_c_225_n 0.00156053f $X=-0.045 $Y=0 $X2=1.05 $Y2=0.74
cc_33 N_GND_c_4_p N_Y_c_225_n 0.00736239f $X=1.455 $Y=0.152 $X2=1.05 $Y2=0.74
cc_34 N_GND_c_5_p N_Y_c_225_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.05 $Y2=0.74
cc_35 N_GND_M1003_b N_Y_c_228_n 0.0225607f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.96
cc_36 N_GND_M1003_b N_Y_c_229_n 0.0136455f $X=-0.045 $Y=0 $X2=1.465 $Y2=1.22
cc_37 N_GND_c_20_p N_Y_c_229_n 0.00646494f $X=1.54 $Y=0.74 $X2=1.465 $Y2=1.22
cc_38 N_GND_M1003_b N_Y_c_231_n 0.00701376f $X=-0.045 $Y=0 $X2=1.195 $Y2=1.22
cc_39 N_GND_c_3_p N_Y_c_231_n 0.0029635f $X=0.26 $Y=0.74 $X2=1.195 $Y2=1.22
cc_40 N_GND_M1003_b Y 0.0092181f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.81
cc_41 N_GND_M1003_b N_Y_c_234_n 0.0114144f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.96
cc_42 N_VDD_M1000_b N_A0_M1000_g 0.0262808f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_43 N_VDD_c_43_p N_A0_M1000_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_44 N_VDD_c_44_p N_A0_M1000_g 0.00354579f $X=0.69 $Y=4.235 $X2=0.475 $Y2=3.825
cc_45 N_VDD_c_45_p N_A0_M1000_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=3.825
cc_46 N_VDD_M1000_b N_A0_c_76_n 0.00618364f $X=-0.045 $Y=2.645 $X2=0.385
+ $Y2=2.505
cc_47 N_VDD_M1000_d A0 0.00614677f $X=0.55 $Y=2.825 $X2=0.385 $Y2=3.07
cc_48 N_VDD_M1000_b N_A1_M1004_g 0.0193713f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_49 N_VDD_c_44_p N_A1_M1004_g 0.00354579f $X=0.69 $Y=4.235 $X2=0.905 $Y2=3.825
cc_50 N_VDD_c_50_p N_A1_M1004_g 0.00496961f $X=1.02 $Y=5.33 $X2=0.905 $Y2=3.825
cc_51 N_VDD_c_45_p N_A1_M1004_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.905 $Y2=3.825
cc_52 N_VDD_M1000_b N_A1_c_110_n 0.00476834f $X=-0.045 $Y=2.645 $X2=0.725
+ $Y2=2.7
cc_53 N_VDD_M1000_b A1 0.0103281f $X=-0.045 $Y=2.645 $X2=0.725 $Y2=2.7
cc_54 N_VDD_M1000_b N_B0_M1001_g 0.0250679f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=3.825
cc_55 N_VDD_c_50_p N_B0_M1001_g 0.00496961f $X=1.02 $Y=5.33 $X2=1.335 $Y2=3.825
cc_56 N_VDD_c_45_p N_B0_M1001_g 0.00429146f $X=1.02 $Y=5.36 $X2=1.335 $Y2=3.825
cc_57 N_VDD_M1000_b N_A_27_565#_c_209_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.895
cc_58 N_VDD_c_43_p N_A_27_565#_c_209_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.895
cc_59 N_VDD_c_45_p N_A_27_565#_c_209_n 0.00435496f $X=1.02 $Y=5.36 $X2=0.26
+ $Y2=3.895
cc_60 N_VDD_M1000_d N_A_27_565#_c_212_n 0.00744208f $X=0.55 $Y=2.825 $X2=1.035
+ $Y2=3.73
cc_61 N_VDD_c_44_p N_A_27_565#_c_212_n 0.0135055f $X=0.69 $Y=4.235 $X2=1.035
+ $Y2=3.73
cc_62 N_VDD_M1000_b N_A_27_565#_c_214_n 0.00198641f $X=-0.045 $Y=2.645 $X2=1.12
+ $Y2=3.895
cc_63 N_VDD_c_50_p N_A_27_565#_c_214_n 0.0045126f $X=1.02 $Y=5.33 $X2=1.12
+ $Y2=3.895
cc_64 N_VDD_c_45_p N_A_27_565#_c_214_n 0.00434939f $X=1.02 $Y=5.36 $X2=1.12
+ $Y2=3.895
cc_65 N_VDD_M1000_b N_Y_c_228_n 0.00960991f $X=-0.045 $Y=2.645 $X2=1.55 $Y2=1.96
cc_66 N_VDD_c_50_p N_Y_c_228_n 0.00477009f $X=1.02 $Y=5.33 $X2=1.55 $Y2=1.96
cc_67 N_VDD_c_45_p N_Y_c_228_n 0.00435496f $X=1.02 $Y=5.36 $X2=1.55 $Y2=1.96
cc_68 N_A0_c_68_n N_A1_M1002_g 0.00899556f $X=0.295 $Y=2.37 $X2=0.835 $Y2=0.945
cc_69 N_A0_c_69_n N_A1_M1002_g 0.069959f $X=0.475 $Y=1.43 $X2=0.835 $Y2=0.945
cc_70 N_A0_c_68_n N_A1_M1004_g 0.00367405f $X=0.295 $Y=2.37 $X2=0.905 $Y2=3.825
cc_71 N_A0_c_75_n N_A1_M1004_g 0.0814351f $X=0.475 $Y=2.505 $X2=0.905 $Y2=3.825
cc_72 N_A0_c_76_n N_A1_M1004_g 0.00277246f $X=0.385 $Y=2.505 $X2=0.905 $Y2=3.825
cc_73 A0 N_A1_M1004_g 0.00309207f $X=0.385 $Y=3.07 $X2=0.905 $Y2=3.825
cc_74 N_A0_c_68_n N_A1_c_109_n 0.0125472f $X=0.295 $Y=2.37 $X2=0.815 $Y2=1.995
cc_75 N_A0_c_68_n N_A1_c_110_n 0.00365573f $X=0.295 $Y=2.37 $X2=0.725 $Y2=2.7
cc_76 N_A0_c_75_n N_A1_c_110_n 0.00281397f $X=0.475 $Y=2.505 $X2=0.725 $Y2=2.7
cc_77 N_A0_c_76_n N_A1_c_110_n 0.0297299f $X=0.385 $Y=2.505 $X2=0.725 $Y2=2.7
cc_78 N_A0_c_68_n N_A1_c_111_n 0.00661569f $X=0.295 $Y=2.37 $X2=0.815 $Y2=1.995
cc_79 N_A0_c_75_n A1 0.00417236f $X=0.475 $Y=2.505 $X2=0.725 $Y2=2.7
cc_80 N_A0_c_76_n A1 0.00775911f $X=0.385 $Y=2.505 $X2=0.725 $Y2=2.7
cc_81 A0 A1 0.00560453f $X=0.385 $Y=3.07 $X2=0.725 $Y2=2.7
cc_82 N_A0_c_76_n N_A_27_565#_M1000_s 0.00883759f $X=0.385 $Y=2.505 $X2=0.135
+ $Y2=2.825
cc_83 A0 N_A_27_565#_M1000_s 0.0125212f $X=0.385 $Y=3.07 $X2=0.135 $Y2=2.825
cc_84 N_A0_M1000_g N_A_27_565#_c_212_n 0.0153088f $X=0.475 $Y=3.825 $X2=1.035
+ $Y2=3.73
cc_85 N_A0_c_76_n N_A_27_565#_c_212_n 0.00147075f $X=0.385 $Y=2.505 $X2=1.035
+ $Y2=3.73
cc_86 A0 N_A_27_565#_c_212_n 0.00792094f $X=0.385 $Y=3.07 $X2=1.035 $Y2=3.73
cc_87 N_A0_c_76_n N_A_27_565#_c_222_n 9.53261e-19 $X=0.385 $Y=2.505 $X2=0.345
+ $Y2=3.73
cc_88 A0 N_A_27_565#_c_222_n 0.00360346f $X=0.385 $Y=3.07 $X2=0.345 $Y2=3.73
cc_89 N_A0_c_69_n N_Y_c_231_n 0.00104729f $X=0.475 $Y=1.43 $X2=1.195 $Y2=1.22
cc_90 N_A1_M1002_g N_B0_M1005_g 0.0276778f $X=0.835 $Y=0.945 $X2=1.325 $Y2=0.835
cc_91 N_A1_c_109_n N_B0_c_160_n 0.0147459f $X=0.815 $Y=1.995 $X2=1.47 $Y2=2.485
cc_92 N_A1_M1004_g N_B0_c_161_n 0.0631994f $X=0.905 $Y=3.825 $X2=1.47 $Y2=2.56
cc_93 A1 N_B0_c_161_n 0.00105858f $X=0.725 $Y=2.7 $X2=1.47 $Y2=2.56
cc_94 N_A1_M1002_g N_B0_c_162_n 0.0039494f $X=0.835 $Y=0.945 $X2=1.47 $Y2=1.6
cc_95 N_A1_M1002_g N_B0_c_164_n 0.00326852f $X=0.835 $Y=0.945 $X2=1.165 $Y2=2.33
cc_96 N_A1_c_109_n N_B0_c_164_n 0.00506769f $X=0.815 $Y=1.995 $X2=1.165 $Y2=2.33
cc_97 N_A1_c_110_n N_B0_c_164_n 0.0109205f $X=0.725 $Y=2.7 $X2=1.165 $Y2=2.33
cc_98 N_A1_c_111_n N_B0_c_164_n 0.0226306f $X=0.815 $Y=1.995 $X2=1.165 $Y2=2.33
cc_99 N_A1_M1002_g N_B0_c_165_n 0.00477017f $X=0.835 $Y=0.945 $X2=1.25 $Y2=1.6
cc_100 N_A1_M1004_g B0 0.00717682f $X=0.905 $Y=3.825 $X2=1.165 $Y2=2.33
cc_101 N_A1_c_110_n B0 0.00705035f $X=0.725 $Y=2.7 $X2=1.165 $Y2=2.33
cc_102 A1 B0 0.00582284f $X=0.725 $Y=2.7 $X2=1.165 $Y2=2.33
cc_103 N_A1_M1004_g N_A_27_565#_c_212_n 0.0180368f $X=0.905 $Y=3.825 $X2=1.035
+ $Y2=3.73
cc_104 N_A1_M1002_g N_Y_c_225_n 0.00112545f $X=0.835 $Y=0.945 $X2=1.05 $Y2=0.74
cc_105 N_A1_c_109_n N_Y_c_225_n 3.56057e-19 $X=0.815 $Y=1.995 $X2=1.05 $Y2=0.74
cc_106 N_A1_M1004_g N_Y_c_228_n 8.50177e-19 $X=0.905 $Y=3.825 $X2=1.55 $Y2=1.96
cc_107 N_A1_c_110_n N_Y_c_228_n 0.00666053f $X=0.725 $Y=2.7 $X2=1.55 $Y2=1.96
cc_108 A1 N_Y_c_228_n 0.00511095f $X=0.725 $Y=2.7 $X2=1.55 $Y2=1.96
cc_109 N_A1_M1002_g N_Y_c_231_n 0.00407967f $X=0.835 $Y=0.945 $X2=1.195 $Y2=1.22
cc_110 N_A1_c_109_n N_Y_c_231_n 0.00171207f $X=0.815 $Y=1.995 $X2=1.195 $Y2=1.22
cc_111 N_A1_M1002_g Y 3.27704e-19 $X=0.835 $Y=0.945 $X2=1.55 $Y2=1.81
cc_112 N_B0_M1005_g N_Y_c_225_n 0.0112072f $X=1.325 $Y=0.835 $X2=1.05 $Y2=0.74
cc_113 N_B0_c_165_n N_Y_c_225_n 0.00317724f $X=1.25 $Y=1.6 $X2=1.05 $Y2=0.74
cc_114 N_B0_M1001_g N_Y_c_228_n 0.0169896f $X=1.335 $Y=3.825 $X2=1.55 $Y2=1.96
cc_115 N_B0_c_160_n N_Y_c_228_n 0.0192649f $X=1.47 $Y=2.485 $X2=1.55 $Y2=1.96
cc_116 N_B0_c_161_n N_Y_c_228_n 0.00834782f $X=1.47 $Y=2.56 $X2=1.55 $Y2=1.96
cc_117 N_B0_c_162_n N_Y_c_228_n 0.00170788f $X=1.47 $Y=1.6 $X2=1.55 $Y2=1.96
cc_118 N_B0_c_164_n N_Y_c_228_n 0.027719f $X=1.165 $Y=2.33 $X2=1.55 $Y2=1.96
cc_119 N_B0_c_166_n N_Y_c_228_n 0.0101032f $X=1.53 $Y=1.6 $X2=1.55 $Y2=1.96
cc_120 B0 N_Y_c_228_n 0.00715529f $X=1.165 $Y=2.33 $X2=1.55 $Y2=1.96
cc_121 N_B0_M1005_g N_Y_c_229_n 0.0119364f $X=1.325 $Y=0.835 $X2=1.465 $Y2=1.22
cc_122 N_B0_c_162_n N_Y_c_229_n 0.00145385f $X=1.47 $Y=1.6 $X2=1.465 $Y2=1.22
cc_123 N_B0_c_165_n N_Y_c_229_n 0.0028071f $X=1.25 $Y=1.6 $X2=1.465 $Y2=1.22
cc_124 N_B0_c_166_n N_Y_c_229_n 0.00718449f $X=1.53 $Y=1.6 $X2=1.465 $Y2=1.22
cc_125 N_B0_M1005_g N_Y_c_231_n 6.90188e-19 $X=1.325 $Y=0.835 $X2=1.195 $Y2=1.22
cc_126 N_B0_c_165_n N_Y_c_231_n 0.00487807f $X=1.25 $Y=1.6 $X2=1.195 $Y2=1.22
cc_127 N_B0_M1005_g Y 0.00272607f $X=1.325 $Y=0.835 $X2=1.55 $Y2=1.81
cc_128 N_B0_c_160_n Y 0.00138242f $X=1.47 $Y=2.485 $X2=1.55 $Y2=1.81
cc_129 N_B0_c_162_n Y 0.01116f $X=1.47 $Y=1.6 $X2=1.55 $Y2=1.81
cc_130 N_B0_c_164_n Y 0.00642461f $X=1.165 $Y=2.33 $X2=1.55 $Y2=1.81
cc_131 N_B0_c_166_n Y 0.0201061f $X=1.53 $Y=1.6 $X2=1.55 $Y2=1.81
cc_132 N_B0_c_160_n N_Y_c_234_n 0.00517151f $X=1.47 $Y=2.485 $X2=1.55 $Y2=1.96
cc_133 N_B0_c_162_n N_Y_c_234_n 8.18646e-19 $X=1.47 $Y=1.6 $X2=1.55 $Y2=1.96
cc_134 N_B0_c_164_n N_Y_c_234_n 0.00655582f $X=1.165 $Y=2.33 $X2=1.55 $Y2=1.96
cc_135 N_B0_c_166_n N_Y_c_234_n 0.00439213f $X=1.53 $Y=1.6 $X2=1.55 $Y2=1.96
