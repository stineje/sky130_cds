* File: sky130_osu_sc_18T_ls__mux2_1.pex.spice
* Created: Thu Oct 29 17:37:02 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%GND 1 20 24 30 32
r35 30 32 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r36 22 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r37 20 22 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r38 20 35 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r39 20 35 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r40 20 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.17
+ $X2=2.38 $Y2=0.17
r41 20 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r42 1 24 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%VDD 1 7 11 17 23
r30 17 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.38 $Y=6.49
+ $X2=2.38 $Y2=6.49
r31 15 23 76.8925 $w=3.03e-07 $l=2.035e-06 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=2.38 $Y2=6.507
r32 11 14 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r33 9 15 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.345 $Y2=6.507
r34 9 14 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r35 7 23 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r36 1 14 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r37 1 11 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%A_110_115# 1 2 7 9 13 17 21 24 27 34 40
+ 45 48
c69 7 0 3.63536e-20 $X=1.35 $Y=1.79
r70 41 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.69
+ $X2=1.09 $Y2=2.69
r71 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.69 $X2=0.925 $Y2=2.69
r72 37 40 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=2.69
+ $X2=0.925 $Y2=2.69
r73 35 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.85
+ $X2=1.09 $Y2=1.85
r74 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.85 $X2=0.925 $Y2=1.85
r75 31 34 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.925 $Y2=1.85
r76 27 29 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r77 25 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.855
+ $X2=0.69 $Y2=2.69
r78 25 27 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.69 $Y=2.855 $X2=0.69
+ $Y2=3.455
r79 24 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.525
+ $X2=0.69 $Y2=2.69
r80 23 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.015
+ $X2=0.69 $Y2=1.85
r81 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.69 $Y=2.015
+ $X2=0.69 $Y2=2.525
r82 19 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.685
+ $X2=0.69 $Y2=1.85
r83 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.69 $Y=1.685
+ $X2=0.69 $Y2=0.825
r84 15 17 964 $w=1.5e-07 $l=1.88e-06 $layer=POLY_cond $X=1.855 $Y=2.705
+ $X2=1.855 $Y2=4.585
r85 11 13 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.425 $Y=1.715
+ $X2=1.425 $Y2=1.075
r86 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.63
+ $X2=1.855 $Y2=2.705
r87 9 48 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.78 $Y=2.63 $X2=1.09
+ $Y2=2.63
r88 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=1.79
+ $X2=1.425 $Y2=1.715
r89 7 45 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.35 $Y=1.79 $X2=1.09
+ $Y2=1.79
r90 2 29 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r91 2 27 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r92 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%S0 3 8 9 11 12 13 15 18 21 26 30
c65 8 0 1.8854e-20 $X=0.475 $Y=4.585
r66 29 30 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.305
+ $X2=0.55 $Y2=2.305
r67 27 29 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.305
+ $X2=0.475 $Y2=2.305
r68 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.305 $X2=0.27 $Y2=2.305
r69 23 26 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=2.305
r70 21 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r71 16 18 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.855 $Y=2.195
+ $X2=1.855 $Y2=1.075
r72 13 15 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.425 $Y=6.16
+ $X2=1.425 $Y2=4.585
r73 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=6.235
+ $X2=1.425 $Y2=6.16
r74 11 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.35 $Y=6.235 $X2=0.55
+ $Y2=6.235
r75 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.27
+ $X2=1.855 $Y2=2.195
r76 9 30 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.78 $Y=2.27
+ $X2=0.55 $Y2=2.27
r77 6 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=6.16
+ $X2=0.55 $Y2=6.235
r78 6 8 807.606 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=6.16
+ $X2=0.475 $Y2=4.585
r79 5 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=2.305
r80 5 8 1084.5 $w=1.5e-07 $l=2.115e-06 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=4.585
r81 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.14
+ $X2=0.475 $Y2=2.305
r82 1 3 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=0.475 $Y=2.14
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%A0 1 2 9 13 19 22 24 26
c41 24 0 1.8854e-20 $X=1.265 $Y=2.96
r42 24 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.265 $Y=2.96
+ $X2=1.265 $Y2=2.96
r43 21 26 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.265 $Y=3.115
+ $X2=1.265 $Y2=2.96
r44 21 22 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=3.115
+ $X2=1.237 $Y2=3.285
r45 19 26 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=1.265 $Y=1.505
+ $X2=1.265 $Y2=2.96
r46 18 19 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=1.335
+ $X2=1.237 $Y2=1.505
r47 13 15 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.21 $Y=3.455
+ $X2=1.21 $Y2=5.835
r48 13 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.21 $Y=3.455
+ $X2=1.21 $Y2=3.285
r49 9 18 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.21 $Y=0.825
+ $X2=1.21 $Y2=1.335
r50 2 15 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=1.085
+ $Y=3.085 $X2=1.21 $Y2=5.835
r51 2 13 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=1.085
+ $Y=3.085 $X2=1.21 $Y2=3.455
r52 1 9 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%Y 1 2 8 10 14 16 20
c37 14 0 3.63536e-20 $X=1.64 $Y=2.22
r38 27 29 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.64 $Y=3.455
+ $X2=1.64 $Y2=5.835
r39 16 27 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.64 $Y=2.22
+ $X2=1.64 $Y2=3.455
r40 14 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=2.22
+ $X2=1.64 $Y2=2.22
r41 11 20 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.64 $Y=1.48
+ $X2=1.64 $Y2=0.825
r42 10 11 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.48
+ $X2=1.64 $Y2=1.48
r43 8 14 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=2.105
+ $X2=1.64 $Y2=2.22
r44 7 10 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=1.595
+ $X2=1.64 $Y2=1.48
r45 7 8 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=1.64 $Y=1.595 $X2=1.64
+ $Y2=2.105
r46 2 29 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=5.835
r47 2 27 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=3.455
r48 1 20 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__MUX2_1%A1 1 2 8 13
r17 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.07 $Y=3.455
+ $X2=2.07 $Y2=5.835
r18 10 17 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.07 $Y=2.59
+ $X2=2.07 $Y2=3.455
r19 10 13 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.07 $Y=2.59
+ $X2=2.07 $Y2=0.825
r20 8 10 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.59 $X2=2.07
+ $Y2=2.59
r21 2 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=5.835
r22 2 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=3.455
r23 1 13 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

