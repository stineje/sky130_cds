* File: sky130_osu_sc_12T_ls__nor2_l.spice
* Created: Fri Nov 12 15:39:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__nor2_l.pex.spice"
.subckt sky130_osu_sc_12T_ls__nor2_l  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_Y_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NSHORT L=0.15 W=0.36
+ AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4 SA=75000.2
+ SB=75000.6 A=0.054 P=1.02 MULT=1
MM1000 N_GND_M1000_d N_A_M1000_g N_Y_M1003_d N_GND_M1003_b NSHORT L=0.15 W=0.36
+ AD=0.0954 AS=0.0504 PD=1.25 PS=0.64 NRD=0 NRS=0 M=1 R=2.4 SA=75000.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1002 A_110_605# N_B_M1002_g N_Y_M1002_s N_VDD_M1002_b PHIGHVT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g A_110_605# N_VDD_M1002_b PHIGHVT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX4_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=2.49275 P=6.33
pX5_noxref noxref_7 Y Y PROBETYPE=1
pX6_noxref noxref_8 B B PROBETYPE=1
pX7_noxref noxref_9 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__nor2_l.pxi.spice"
*
.ends
*
*
