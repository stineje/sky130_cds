* File: sky130_osu_sc_18T_ms__oai22_l.pxi.spice
* Created: Fri Nov 12 14:05:53 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%GND N_GND_M1004_d N_GND_M1004_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_MS__OAI22_L%GND
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%VDD N_VDD_M1005_s N_VDD_M1007_d N_VDD_M1005_b
+ N_VDD_c_45_p N_VDD_c_46_p N_VDD_c_64_p VDD N_VDD_c_47_p
+ PM_SKY130_OSU_SC_18T_MS__OAI22_L%VDD
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%A0 N_A0_c_70_n N_A0_M1004_g N_A0_M1005_g
+ N_A0_c_74_n N_A0_c_75_n N_A0_c_76_n N_A0_c_77_n A0
+ PM_SKY130_OSU_SC_18T_MS__OAI22_L%A0
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%A1 N_A1_M1002_g N_A1_M1000_g N_A1_c_110_n
+ N_A1_c_111_n N_A1_c_112_n A1 PM_SKY130_OSU_SC_18T_MS__OAI22_L%A1
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%B0 N_B0_M1001_g N_B0_M1003_g N_B0_c_159_n
+ N_B0_c_160_n N_B0_c_161_n B0 PM_SKY130_OSU_SC_18T_MS__OAI22_L%B0
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%B1 N_B1_M1007_g N_B1_M1006_g N_B1_c_209_n
+ N_B1_c_210_n N_B1_c_211_n N_B1_c_212_n B1 PM_SKY130_OSU_SC_18T_MS__OAI22_L%B1
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_242_n
+ N_Y_c_254_n N_Y_c_246_n N_Y_c_257_n N_Y_c_285_p N_Y_c_238_n N_Y_c_239_n
+ N_Y_c_240_n Y PM_SKY130_OSU_SC_18T_MS__OAI22_L%Y
x_PM_SKY130_OSU_SC_18T_MS__OAI22_L%A_27_115# N_A_27_115#_M1004_s
+ N_A_27_115#_M1000_d N_A_27_115#_M1006_d N_A_27_115#_c_287_n
+ N_A_27_115#_c_290_n N_A_27_115#_c_297_n N_A_27_115#_c_292_n
+ N_A_27_115#_c_294_n PM_SKY130_OSU_SC_18T_MS__OAI22_L%A_27_115#
cc_1 N_GND_M1004_b N_A0_c_70_n 0.0246907f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.7
cc_2 N_GND_c_2_p N_A0_c_70_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.7
cc_3 N_GND_c_3_p N_A0_c_70_n 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.7
cc_4 N_GND_c_4_p N_A0_c_70_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=1.7
cc_5 N_GND_M1004_b N_A0_c_74_n 0.0245188f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.775
cc_6 N_GND_M1004_b N_A0_c_75_n 0.0342831f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.76
cc_7 N_GND_M1004_b N_A0_c_76_n 0.0617323f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.595
cc_8 N_GND_M1004_b N_A0_c_77_n 0.0028102f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.76
cc_9 N_GND_M1004_b N_A1_M1002_g 0.0270201f $X=-0.045 $Y=0 $X2=0.835 $Y2=4.585
cc_10 N_GND_M1004_b N_A1_M1000_g 0.0443528f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.075
cc_11 N_GND_c_3_p N_A1_M1000_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905 $Y2=1.075
cc_12 N_GND_c_4_p N_A1_M1000_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.905 $Y2=1.075
cc_13 N_GND_M1004_b N_A1_c_110_n 0.0318892f $X=-0.045 $Y=0 $X2=0.815 $Y2=2.22
cc_14 N_GND_M1004_b N_A1_c_111_n 0.00628302f $X=-0.045 $Y=0 $X2=0.815 $Y2=2.22
cc_15 N_GND_M1004_b N_A1_c_112_n 0.00134829f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.96
cc_16 N_GND_M1004_b A1 0.00271527f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.96
cc_17 N_GND_M1004_b N_B0_M1001_g 0.0226011f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.075
cc_18 N_GND_c_4_p N_B0_M1001_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335 $Y2=1.075
cc_19 N_GND_M1004_b N_B0_M1003_g 0.0437024f $X=-0.045 $Y=0 $X2=1.335 $Y2=4.585
cc_20 N_GND_M1004_b N_B0_c_159_n 0.028787f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.88
cc_21 N_GND_M1004_b N_B0_c_160_n 0.00518014f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.59
cc_22 N_GND_M1004_b N_B0_c_161_n 0.00424299f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.88
cc_23 N_GND_M1004_b B0 0.0129888f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.59
cc_24 N_GND_M1004_b N_B1_M1006_g 0.0549493f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.075
cc_25 N_GND_c_4_p N_B1_M1006_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765 $Y2=1.075
cc_26 N_GND_M1004_b N_B1_c_209_n 0.0319209f $X=-0.045 $Y=0 $X2=1.73 $Y2=2.81
cc_27 N_GND_M1004_b N_B1_c_210_n 0.00983533f $X=-0.045 $Y=0 $X2=1.73 $Y2=2.96
cc_28 N_GND_M1004_b N_B1_c_211_n 0.0576947f $X=-0.045 $Y=0 $X2=2.005 $Y2=2.225
cc_29 N_GND_M1004_b N_B1_c_212_n 0.0125315f $X=-0.045 $Y=0 $X2=2.005 $Y2=2.225
cc_30 N_GND_M1004_b B1 0.00895888f $X=-0.045 $Y=0 $X2=2.005 $Y2=2.225
cc_31 N_GND_M1004_b N_Y_c_238_n 0.00764938f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.85
cc_32 N_GND_M1004_b N_Y_c_239_n 0.00181926f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.735
cc_33 N_GND_M1004_b N_Y_c_240_n 5.70233e-19 $X=-0.045 $Y=0 $X2=1.665 $Y2=1.48
cc_34 N_GND_M1004_b Y 0.00397674f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.85
cc_35 N_GND_M1004_b N_A_27_115#_c_287_n 0.00156053f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_36 N_GND_c_2_p N_A_27_115#_c_287_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_37 N_GND_c_4_p N_A_27_115#_c_287_n 0.00476261f $X=1.7 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_38 N_GND_M1004_d N_A_27_115#_c_290_n 0.00580138f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.42
cc_39 N_GND_c_3_p N_A_27_115#_c_290_n 0.00986105f $X=0.69 $Y=0.825 $X2=1.035
+ $Y2=1.42
cc_40 N_GND_M1004_b N_A_27_115#_c_292_n 0.0321475f $X=-0.045 $Y=0 $X2=1.895
+ $Y2=0.66
cc_41 N_GND_c_4_p N_A_27_115#_c_292_n 0.0233363f $X=1.7 $Y=0.19 $X2=1.895
+ $Y2=0.66
cc_42 N_GND_M1004_b N_A_27_115#_c_294_n 0.00893451f $X=-0.045 $Y=0 $X2=1.205
+ $Y2=0.66
cc_43 N_GND_c_4_p N_A_27_115#_c_294_n 0.0048048f $X=1.7 $Y=0.19 $X2=1.205
+ $Y2=0.66
cc_44 N_VDD_M1005_b N_A0_M1005_g 0.0204563f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_45 N_VDD_c_45_p N_A0_M1005_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_46 N_VDD_c_46_p N_A0_M1005_g 0.00606474f $X=1.825 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_47 N_VDD_c_47_p N_A0_M1005_g 0.00468827f $X=1.7 $Y=6.47 $X2=0.475 $Y2=4.585
cc_48 N_VDD_M1005_b N_A0_c_75_n 0.0059005f $X=-0.045 $Y=2.905 $X2=0.415 $Y2=2.76
cc_49 N_VDD_M1005_s N_A0_c_77_n 0.00849866f $X=0.135 $Y=3.085 $X2=0.415 $Y2=2.76
cc_50 N_VDD_M1005_b N_A0_c_77_n 0.00549657f $X=-0.045 $Y=2.905 $X2=0.415
+ $Y2=2.76
cc_51 N_VDD_c_45_p N_A0_c_77_n 2.89251e-19 $X=0.26 $Y=4.135 $X2=0.415 $Y2=2.76
cc_52 N_VDD_M1005_s A0 0.0139414f $X=0.135 $Y=3.085 $X2=0.415 $Y2=3.33
cc_53 N_VDD_c_45_p A0 0.00289954f $X=0.26 $Y=4.135 $X2=0.415 $Y2=3.33
cc_54 N_VDD_M1005_b N_A1_M1002_g 0.0186099f $X=-0.045 $Y=2.905 $X2=0.835
+ $Y2=4.585
cc_55 N_VDD_c_46_p N_A1_M1002_g 0.00606474f $X=1.825 $Y=6.507 $X2=0.835
+ $Y2=4.585
cc_56 N_VDD_c_47_p N_A1_M1002_g 0.00468827f $X=1.7 $Y=6.47 $X2=0.835 $Y2=4.585
cc_57 N_VDD_M1005_b N_A1_c_112_n 0.00395559f $X=-0.045 $Y=2.905 $X2=0.895
+ $Y2=2.96
cc_58 N_VDD_M1005_b A1 0.00722999f $X=-0.045 $Y=2.905 $X2=0.895 $Y2=2.96
cc_59 N_VDD_M1005_b N_B0_M1003_g 0.0205368f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=4.585
cc_60 N_VDD_c_46_p N_B0_M1003_g 0.00606474f $X=1.825 $Y=6.507 $X2=1.335
+ $Y2=4.585
cc_61 N_VDD_c_47_p N_B0_M1003_g 0.00468827f $X=1.7 $Y=6.47 $X2=1.335 $Y2=4.585
cc_62 N_VDD_M1005_b N_B1_c_210_n 0.028286f $X=-0.045 $Y=2.905 $X2=1.73 $Y2=2.96
cc_63 N_VDD_c_46_p N_B1_c_210_n 0.00606474f $X=1.825 $Y=6.507 $X2=1.73 $Y2=2.96
cc_64 N_VDD_c_64_p N_B1_c_210_n 0.00713292f $X=1.91 $Y=4.135 $X2=1.73 $Y2=2.96
cc_65 N_VDD_c_47_p N_B1_c_210_n 0.00468827f $X=1.7 $Y=6.47 $X2=1.73 $Y2=2.96
cc_66 N_VDD_M1005_b N_Y_c_242_n 0.00156987f $X=-0.045 $Y=2.905 $X2=1.085
+ $Y2=3.795
cc_67 N_VDD_c_46_p N_Y_c_242_n 0.00738471f $X=1.825 $Y=6.507 $X2=1.085 $Y2=3.795
cc_68 N_VDD_c_47_p N_Y_c_242_n 0.00476747f $X=1.7 $Y=6.47 $X2=1.085 $Y2=3.795
cc_69 N_VDD_M1005_b N_Y_c_238_n 0.00136067f $X=-0.045 $Y=2.905 $X2=1.665
+ $Y2=1.85
cc_70 N_A0_c_75_n N_A1_M1002_g 0.216534f $X=0.415 $Y=2.76 $X2=0.835 $Y2=4.585
cc_71 N_A0_c_76_n N_A1_M1002_g 0.00799469f $X=0.415 $Y=2.595 $X2=0.835 $Y2=4.585
cc_72 N_A0_c_77_n N_A1_M1002_g 0.00302464f $X=0.415 $Y=2.76 $X2=0.835 $Y2=4.585
cc_73 A0 N_A1_M1002_g 0.00376364f $X=0.415 $Y=3.33 $X2=0.835 $Y2=4.585
cc_74 N_A0_c_70_n N_A1_M1000_g 0.0442543f $X=0.475 $Y=1.7 $X2=0.905 $Y2=1.075
cc_75 N_A0_c_76_n N_A1_M1000_g 0.00745307f $X=0.415 $Y=2.595 $X2=0.905 $Y2=1.075
cc_76 N_A0_c_76_n N_A1_c_110_n 0.0167307f $X=0.415 $Y=2.595 $X2=0.815 $Y2=2.22
cc_77 N_A0_c_75_n N_A1_c_111_n 0.00128494f $X=0.415 $Y=2.76 $X2=0.815 $Y2=2.22
cc_78 N_A0_c_76_n N_A1_c_111_n 0.00640175f $X=0.415 $Y=2.595 $X2=0.815 $Y2=2.22
cc_79 N_A0_c_77_n N_A1_c_111_n 0.0241512f $X=0.415 $Y=2.76 $X2=0.815 $Y2=2.22
cc_80 N_A0_M1005_g N_A1_c_112_n 0.00128494f $X=0.475 $Y=4.585 $X2=0.895 $Y2=2.96
cc_81 N_A0_M1005_g A1 4.3358e-19 $X=0.475 $Y=4.585 $X2=0.895 $Y2=2.96
cc_82 N_A0_c_77_n A1 0.00249278f $X=0.415 $Y=2.76 $X2=0.895 $Y2=2.96
cc_83 A0 A_110_617# 0.0129699f $X=0.415 $Y=3.33 $X2=0.55 $Y2=3.085
cc_84 N_A0_c_77_n N_Y_c_246_n 0.00152664f $X=0.415 $Y=2.76 $X2=1.17 $Y2=3.415
cc_85 A0 N_Y_c_246_n 0.00392194f $X=0.415 $Y=3.33 $X2=1.17 $Y2=3.415
cc_86 N_A0_c_70_n N_A_27_115#_c_290_n 0.0198204f $X=0.475 $Y=1.7 $X2=1.035
+ $Y2=1.42
cc_87 N_A0_c_74_n N_A_27_115#_c_297_n 0.0030143f $X=0.475 $Y=1.775 $X2=0.345
+ $Y2=1.42
cc_88 N_A1_M1000_g N_B0_M1001_g 0.0242274f $X=0.905 $Y=1.075 $X2=1.335 $Y2=1.075
cc_89 N_A1_M1002_g N_B0_M1003_g 0.046277f $X=0.835 $Y=4.585 $X2=1.335 $Y2=4.585
cc_90 N_A1_M1000_g N_B0_M1003_g 0.0130769f $X=0.905 $Y=1.075 $X2=1.335 $Y2=4.585
cc_91 N_A1_c_111_n N_B0_M1003_g 0.00185146f $X=0.815 $Y=2.22 $X2=1.335 $Y2=4.585
cc_92 N_A1_c_112_n N_B0_M1003_g 0.00125927f $X=0.895 $Y=2.96 $X2=1.335 $Y2=4.585
cc_93 A1 N_B0_M1003_g 0.0039398f $X=0.895 $Y=2.96 $X2=1.335 $Y2=4.585
cc_94 N_A1_M1000_g N_B0_c_159_n 0.0194179f $X=0.905 $Y=1.075 $X2=1.325 $Y2=1.88
cc_95 N_A1_M1002_g N_B0_c_160_n 0.00190813f $X=0.835 $Y=4.585 $X2=1.2 $Y2=2.59
cc_96 N_A1_M1000_g N_B0_c_160_n 0.00235131f $X=0.905 $Y=1.075 $X2=1.2 $Y2=2.59
cc_97 N_A1_c_111_n N_B0_c_160_n 0.0346786f $X=0.815 $Y=2.22 $X2=1.2 $Y2=2.59
cc_98 N_A1_M1000_g N_B0_c_161_n 0.00763077f $X=0.905 $Y=1.075 $X2=1.325 $Y2=1.88
cc_99 N_A1_M1002_g B0 0.00416458f $X=0.835 $Y=4.585 $X2=1.2 $Y2=2.59
cc_100 N_A1_c_110_n B0 0.00100952f $X=0.815 $Y=2.22 $X2=1.2 $Y2=2.59
cc_101 N_A1_c_111_n B0 0.00821238f $X=0.815 $Y=2.22 $X2=1.2 $Y2=2.59
cc_102 N_A1_c_112_n B0 2.4196e-19 $X=0.895 $Y=2.96 $X2=1.2 $Y2=2.59
cc_103 A1 B0 0.0191116f $X=0.895 $Y=2.96 $X2=1.2 $Y2=2.59
cc_104 N_A1_M1002_g N_Y_c_242_n 0.0258582f $X=0.835 $Y=4.585 $X2=1.085 $Y2=3.795
cc_105 N_A1_M1002_g N_Y_c_246_n 0.00383489f $X=0.835 $Y=4.585 $X2=1.17 $Y2=3.415
cc_106 A1 N_Y_c_246_n 0.00669635f $X=0.895 $Y=2.96 $X2=1.17 $Y2=3.415
cc_107 N_A1_c_112_n N_Y_c_238_n 0.00278415f $X=0.895 $Y=2.96 $X2=1.665 $Y2=1.85
cc_108 A1 N_Y_c_238_n 0.00663666f $X=0.895 $Y=2.96 $X2=1.665 $Y2=1.85
cc_109 N_A1_M1000_g N_A_27_115#_c_290_n 0.0176072f $X=0.905 $Y=1.075 $X2=1.035
+ $Y2=1.42
cc_110 N_A1_c_110_n N_A_27_115#_c_290_n 0.0022598f $X=0.815 $Y=2.22 $X2=1.035
+ $Y2=1.42
cc_111 N_A1_c_111_n N_A_27_115#_c_290_n 0.0046765f $X=0.815 $Y=2.22 $X2=1.035
+ $Y2=1.42
cc_112 N_B0_M1001_g N_B1_M1006_g 0.0388095f $X=1.335 $Y=1.075 $X2=1.765
+ $Y2=1.075
cc_113 N_B0_M1003_g N_B1_M1006_g 0.0310455f $X=1.335 $Y=4.585 $X2=1.765
+ $Y2=1.075
cc_114 N_B0_c_159_n N_B1_M1006_g 0.0183044f $X=1.325 $Y=1.88 $X2=1.765 $Y2=1.075
cc_115 N_B0_c_160_n N_B1_M1006_g 6.89792e-19 $X=1.2 $Y=2.59 $X2=1.765 $Y2=1.075
cc_116 N_B0_c_161_n N_B1_M1006_g 5.25213e-19 $X=1.325 $Y=1.88 $X2=1.765
+ $Y2=1.075
cc_117 N_B0_M1003_g N_B1_c_210_n 0.20245f $X=1.335 $Y=4.585 $X2=1.73 $Y2=2.96
cc_118 N_B0_M1003_g N_Y_c_242_n 0.0258582f $X=1.335 $Y=4.585 $X2=1.085 $Y2=3.795
cc_119 N_B0_M1003_g N_Y_c_254_n 0.018662f $X=1.335 $Y=4.585 $X2=1.58 $Y2=3.415
cc_120 N_B0_c_160_n N_Y_c_254_n 0.00149518f $X=1.2 $Y=2.59 $X2=1.58 $Y2=3.415
cc_121 N_B0_c_160_n N_Y_c_246_n 9.67699e-19 $X=1.2 $Y=2.59 $X2=1.17 $Y2=3.415
cc_122 N_B0_M1001_g N_Y_c_257_n 0.00163819f $X=1.335 $Y=1.075 $X2=1.55 $Y2=1.245
cc_123 N_B0_M1003_g N_Y_c_238_n 0.0114207f $X=1.335 $Y=4.585 $X2=1.665 $Y2=1.85
cc_124 N_B0_c_159_n N_Y_c_238_n 0.00159117f $X=1.325 $Y=1.88 $X2=1.665 $Y2=1.85
cc_125 N_B0_c_160_n N_Y_c_238_n 0.0260605f $X=1.2 $Y=2.59 $X2=1.665 $Y2=1.85
cc_126 N_B0_c_161_n N_Y_c_238_n 0.0188911f $X=1.325 $Y=1.88 $X2=1.665 $Y2=1.85
cc_127 B0 N_Y_c_238_n 0.00640554f $X=1.2 $Y=2.59 $X2=1.665 $Y2=1.85
cc_128 N_B0_M1001_g N_Y_c_239_n 0.00157615f $X=1.335 $Y=1.075 $X2=1.665
+ $Y2=1.735
cc_129 N_B0_c_159_n N_Y_c_239_n 2.63601e-19 $X=1.325 $Y=1.88 $X2=1.665 $Y2=1.735
cc_130 N_B0_c_161_n N_Y_c_239_n 8.33805e-19 $X=1.325 $Y=1.88 $X2=1.665 $Y2=1.735
cc_131 N_B0_M1001_g N_Y_c_240_n 0.00286422f $X=1.335 $Y=1.075 $X2=1.665 $Y2=1.48
cc_132 N_B0_c_159_n Y 0.00379994f $X=1.325 $Y=1.88 $X2=1.665 $Y2=1.85
cc_133 N_B0_c_161_n Y 0.00762114f $X=1.325 $Y=1.88 $X2=1.665 $Y2=1.85
cc_134 N_B0_c_159_n N_A_27_115#_c_290_n 3.35424e-19 $X=1.325 $Y=1.88 $X2=1.035
+ $Y2=1.42
cc_135 N_B0_c_161_n N_A_27_115#_c_290_n 0.00655381f $X=1.325 $Y=1.88 $X2=1.035
+ $Y2=1.42
cc_136 N_B0_M1001_g N_A_27_115#_c_292_n 0.0130261f $X=1.335 $Y=1.075 $X2=1.895
+ $Y2=0.66
cc_137 N_B1_c_210_n N_Y_c_254_n 0.0176551f $X=1.73 $Y=2.96 $X2=1.58 $Y2=3.415
cc_138 N_B1_M1006_g N_Y_c_257_n 0.0137941f $X=1.765 $Y=1.075 $X2=1.55 $Y2=1.245
cc_139 N_B1_M1006_g N_Y_c_238_n 0.0109293f $X=1.765 $Y=1.075 $X2=1.665 $Y2=1.85
cc_140 N_B1_c_209_n N_Y_c_238_n 0.0207198f $X=1.73 $Y=2.81 $X2=1.665 $Y2=1.85
cc_141 N_B1_c_210_n N_Y_c_238_n 0.0284849f $X=1.73 $Y=2.96 $X2=1.665 $Y2=1.85
cc_142 N_B1_c_211_n N_Y_c_238_n 0.00828193f $X=2.005 $Y=2.225 $X2=1.665 $Y2=1.85
cc_143 N_B1_c_212_n N_Y_c_238_n 0.0203078f $X=2.005 $Y=2.225 $X2=1.665 $Y2=1.85
cc_144 B1 N_Y_c_238_n 0.00704472f $X=2.005 $Y=2.225 $X2=1.665 $Y2=1.85
cc_145 N_B1_M1006_g N_Y_c_239_n 0.00516527f $X=1.765 $Y=1.075 $X2=1.665
+ $Y2=1.735
cc_146 N_B1_M1006_g N_Y_c_240_n 0.0116229f $X=1.765 $Y=1.075 $X2=1.665 $Y2=1.48
cc_147 N_B1_M1006_g Y 0.00959795f $X=1.765 $Y=1.075 $X2=1.665 $Y2=1.85
cc_148 B1 Y 0.00540133f $X=2.005 $Y=2.225 $X2=1.665 $Y2=1.85
cc_149 N_B1_M1006_g N_A_27_115#_c_292_n 0.0123847f $X=1.765 $Y=1.075 $X2=1.895
+ $Y2=0.66
cc_150 N_Y_c_254_n A_282_617# 0.00732587f $X=1.58 $Y=3.415 $X2=1.41 $Y2=3.085
cc_151 N_Y_c_240_n N_A_27_115#_c_290_n 0.0029159f $X=1.665 $Y=1.48 $X2=1.035
+ $Y2=1.42
cc_152 N_Y_M1001_d N_A_27_115#_c_292_n 0.00376923f $X=1.41 $Y=0.575 $X2=1.895
+ $Y2=0.66
cc_153 N_Y_c_257_n N_A_27_115#_c_292_n 0.00176198f $X=1.55 $Y=1.245 $X2=1.895
+ $Y2=0.66
cc_154 N_Y_c_285_p N_A_27_115#_c_292_n 0.0129297f $X=1.55 $Y=1.165 $X2=1.895
+ $Y2=0.66
