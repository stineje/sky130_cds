* File: sky130_osu_sc_12T_hs__xnor2_l.pxi.spice
* Created: Fri Nov 12 15:14:07 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%GND N_GND_M1006_d N_GND_M1010_d N_GND_M1006_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_14_p N_GND_c_54_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_HS__XNOR2_L%GND
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%VDD N_VDD_M1000_d N_VDD_M1004_d N_VDD_M1000_b
+ N_VDD_c_79_p N_VDD_c_80_p N_VDD_c_76_p N_VDD_c_94_p N_VDD_c_96_p VDD
+ N_VDD_c_77_p PM_SKY130_OSU_SC_12T_HS__XNOR2_L%VDD
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A N_A_c_115_n N_A_M1006_g N_A_M1000_g
+ N_A_c_119_n N_A_M1002_g N_A_M1003_g N_A_c_122_n N_A_c_123_n N_A_c_124_n
+ N_A_c_125_n N_A_c_126_n N_A_c_130_n N_A_c_131_n N_A_c_133_n N_A_c_134_n
+ N_A_c_136_n N_A_c_137_n A N_A_c_142_n N_A_c_143_n
+ PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A_27_115# N_A_27_115#_M1006_s
+ N_A_27_115#_M1000_s N_A_27_115#_M1009_g N_A_27_115#_c_237_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_240_n N_A_27_115#_c_241_n
+ N_A_27_115#_c_242_n N_A_27_115#_c_245_n N_A_27_115#_c_246_n
+ N_A_27_115#_c_247_n N_A_27_115#_c_248_n
+ PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A_27_115#
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A_238_89# N_A_238_89#_M1007_d
+ N_A_238_89#_M1001_d N_A_238_89#_M1011_g N_A_238_89#_M1005_g
+ N_A_238_89#_c_323_n N_A_238_89#_c_324_n N_A_238_89#_c_325_n
+ N_A_238_89#_c_327_n N_A_238_89#_c_328_n
+ PM_SKY130_OSU_SC_12T_HS__XNOR2_L%A_238_89#
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%B N_B_c_384_n N_B_M1010_g N_B_c_401_n
+ N_B_M1004_g N_B_c_388_n N_B_c_389_n N_B_c_390_n N_B_M1007_g N_B_c_393_n
+ N_B_c_408_n N_B_M1001_g N_B_c_394_n N_B_c_396_n N_B_c_397_n B
+ PM_SKY130_OSU_SC_12T_HS__XNOR2_L%B
x_PM_SKY130_OSU_SC_12T_HS__XNOR2_L%Y N_Y_M1011_d N_Y_M1005_d N_Y_c_441_n
+ N_Y_c_475_n N_Y_c_447_n N_Y_c_442_n Y N_Y_c_446_n N_Y_c_451_n
+ PM_SKY130_OSU_SC_12T_HS__XNOR2_L%Y
cc_1 N_GND_M1006_b N_A_c_115_n 0.0183287f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.2
cc_2 N_GND_c_2_p N_A_c_115_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.2
cc_3 N_GND_c_3_p N_A_c_115_n 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=1.2
cc_4 N_GND_c_4_p N_A_c_115_n 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=1.2
cc_5 N_GND_M1006_b N_A_c_119_n 0.00547593f $X=-0.045 $Y=0 $X2=0.71 $Y2=1.275
cc_6 N_GND_c_3_p N_A_c_119_n 0.00412096f $X=0.69 $Y=0.74 $X2=0.71 $Y2=1.275
cc_7 N_GND_M1006_b N_A_M1003_g 0.0192964f $X=-0.045 $Y=0 $X2=1.865 $Y2=3.235
cc_8 N_GND_M1006_b N_A_c_122_n 0.00962022f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.275
cc_9 N_GND_M1006_b N_A_c_123_n 0.0590857f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.38
cc_10 N_GND_M1006_b N_A_c_124_n 0.00429392f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.53
cc_11 N_GND_M1006_b N_A_c_125_n 0.0219799f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.275
cc_12 N_GND_M1006_b N_A_c_126_n 0.0136685f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.2
cc_13 N_GND_c_3_p N_A_c_126_n 0.00308284f $X=0.69 $Y=0.74 $X2=0.845 $Y2=1.2
cc_14 N_GND_c_14_p N_A_c_126_n 0.00606474f $X=2.355 $Y=0.152 $X2=0.845 $Y2=1.2
cc_15 N_GND_c_4_p N_A_c_126_n 0.00468827f $X=2.38 $Y=0.19 $X2=0.845 $Y2=1.2
cc_16 N_GND_M1006_b N_A_c_130_n 0.0506697f $X=-0.045 $Y=0 $X2=1.865 $Y2=1.955
cc_17 N_GND_M1006_b N_A_c_131_n 0.00124261f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.37
cc_18 N_GND_c_3_p N_A_c_131_n 3.74727e-19 $X=0.69 $Y=0.74 $X2=0.845 $Y2=1.37
cc_19 N_GND_M1006_b N_A_c_133_n 0.00659141f $X=-0.045 $Y=0 $X2=2.105 $Y2=1.74
cc_20 N_GND_M1006_d N_A_c_134_n 4.23026e-19 $X=0.55 $Y=0.575 $X2=0.845 $Y2=1.255
cc_21 N_GND_M1006_b N_A_c_134_n 7.09331e-19 $X=-0.045 $Y=0 $X2=0.845 $Y2=1.255
cc_22 N_GND_c_14_p N_A_c_136_n 0.0087746f $X=2.355 $Y=0.152 $X2=2.02 $Y2=1
cc_23 N_GND_M1006_d N_A_c_137_n 0.00299484f $X=0.55 $Y=0.575 $X2=0.93 $Y2=1
cc_24 N_GND_c_3_p N_A_c_137_n 6.34087e-19 $X=0.69 $Y=0.74 $X2=0.93 $Y2=1
cc_25 N_GND_c_14_p N_A_c_137_n 0.00921136f $X=2.355 $Y=0.152 $X2=0.93 $Y2=1
cc_26 N_GND_M1006_b A 0.00270604f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.37
cc_27 N_GND_c_3_p A 0.00252415f $X=0.69 $Y=0.74 $X2=0.845 $Y2=1.37
cc_28 N_GND_M1006_b N_A_c_142_n 0.0049133f $X=-0.045 $Y=0 $X2=2.105 $Y2=1.74
cc_29 N_GND_M1006_b N_A_c_143_n 0.00512637f $X=-0.045 $Y=0 $X2=2.107 $Y2=1.625
cc_30 N_GND_M1006_b N_A_27_115#_M1009_g 0.0168741f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=3.235
cc_31 N_GND_M1006_b N_A_27_115#_c_237_n 0.0174971f $X=-0.045 $Y=0 $X2=1.865
+ $Y2=1.235
cc_32 N_GND_c_14_p N_A_27_115#_c_237_n 0.00606474f $X=2.355 $Y=0.152 $X2=1.865
+ $Y2=1.235
cc_33 N_GND_c_4_p N_A_27_115#_c_237_n 0.00468827f $X=2.38 $Y=0.19 $X2=1.865
+ $Y2=1.235
cc_34 N_GND_M1006_b N_A_27_115#_c_240_n 0.0277533f $X=-0.045 $Y=0 $X2=0.845
+ $Y2=1.94
cc_35 N_GND_M1006_b N_A_27_115#_c_241_n 0.0364542f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.4
cc_36 N_GND_M1006_b N_A_27_115#_c_242_n 0.0353523f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_37 N_GND_c_2_p N_A_27_115#_c_242_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_38 N_GND_c_4_p N_A_27_115#_c_242_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_39 N_GND_M1006_b N_A_27_115#_c_245_n 0.0186783f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.955
cc_40 N_GND_M1006_b N_A_27_115#_c_246_n 0.0348304f $X=-0.045 $Y=0 $X2=1.68
+ $Y2=1.94
cc_41 N_GND_M1006_b N_A_27_115#_c_247_n 0.00464186f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.4
cc_42 N_GND_M1006_b N_A_27_115#_c_248_n 0.00692367f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.94
cc_43 N_GND_M1006_b N_A_238_89#_M1011_g 0.0686775f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=0.85
cc_44 N_GND_c_14_p N_A_238_89#_M1011_g 0.00606474f $X=2.355 $Y=0.152 $X2=1.265
+ $Y2=0.85
cc_45 N_GND_c_4_p N_A_238_89#_M1011_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.265
+ $Y2=0.85
cc_46 N_GND_M1006_b N_A_238_89#_c_323_n 0.021482f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=2.285
cc_47 N_GND_M1006_b N_A_238_89#_c_324_n 0.0319502f $X=-0.045 $Y=0 $X2=2.785
+ $Y2=2.285
cc_48 N_GND_M1006_b N_A_238_89#_c_325_n 0.0587121f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=0.755
cc_49 N_GND_c_4_p N_A_238_89#_c_325_n 0.00476261f $X=2.38 $Y=0.19 $X2=2.87
+ $Y2=0.755
cc_50 N_GND_M1006_b N_A_238_89#_c_327_n 0.00243339f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=2.955
cc_51 N_GND_M1006_b N_A_238_89#_c_328_n 0.00720662f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=2.285
cc_52 N_GND_M1006_b N_B_c_384_n 0.0135598f $X=-0.045 $Y=0 $X2=2.225 $Y2=1.2
cc_53 N_GND_c_14_p N_B_c_384_n 0.00606474f $X=2.355 $Y=0.152 $X2=2.225 $Y2=1.2
cc_54 N_GND_c_54_p N_B_c_384_n 0.00308284f $X=2.44 $Y=0.74 $X2=2.225 $Y2=1.2
cc_55 N_GND_c_4_p N_B_c_384_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.225 $Y2=1.2
cc_56 N_GND_M1006_b N_B_c_388_n 0.00754663f $X=-0.045 $Y=0 $X2=2.58 $Y2=2.455
cc_57 N_GND_M1006_b N_B_c_389_n 0.00440456f $X=-0.045 $Y=0 $X2=2.3 $Y2=2.455
cc_58 N_GND_M1006_b N_B_c_390_n 0.0243936f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.2
cc_59 N_GND_c_54_p N_B_c_390_n 0.00308284f $X=2.44 $Y=0.74 $X2=2.655 $Y2=1.2
cc_60 N_GND_c_4_p N_B_c_390_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.655 $Y2=1.2
cc_61 N_GND_M1006_b N_B_c_393_n 0.045354f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.38
cc_62 N_GND_M1006_b N_B_c_394_n 0.0482504f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.382
cc_63 N_GND_c_54_p N_B_c_394_n 0.00317391f $X=2.44 $Y=0.74 $X2=2.655 $Y2=1.382
cc_64 N_GND_M1006_b N_B_c_396_n 0.00181559f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.455
cc_65 N_GND_M1006_b N_B_c_397_n 0.00222287f $X=-0.045 $Y=0 $X2=2.53 $Y2=1.37
cc_66 N_GND_c_54_p N_B_c_397_n 0.0031552f $X=2.44 $Y=0.74 $X2=2.53 $Y2=1.37
cc_67 N_GND_M1006_b B 0.00608496f $X=-0.045 $Y=0 $X2=2.53 $Y2=1.4
cc_68 N_GND_c_54_p B 0.00319733f $X=2.44 $Y=0.74 $X2=2.53 $Y2=1.4
cc_69 N_GND_M1006_b N_Y_c_441_n 0.00636628f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.37
cc_70 N_GND_M1006_b N_Y_c_442_n 0.00311548f $X=-0.045 $Y=0 $X2=1.425 $Y2=0.755
cc_71 N_GND_c_14_p N_Y_c_442_n 0.0145361f $X=2.355 $Y=0.152 $X2=1.425 $Y2=0.755
cc_72 N_GND_c_4_p N_Y_c_442_n 0.0108897f $X=2.38 $Y=0.19 $X2=1.425 $Y2=0.755
cc_73 N_GND_M1006_b Y 0.00613557f $X=-0.045 $Y=0 $X2=1.42 $Y2=1.655
cc_74 N_GND_M1006_b N_Y_c_446_n 0.001892f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.37
cc_75 N_VDD_M1000_b N_A_M1003_g 0.0215143f $X=-0.045 $Y=2.425 $X2=1.865
+ $Y2=3.235
cc_76 N_VDD_c_76_p N_A_M1003_g 0.00606474f $X=2.355 $Y=4.287 $X2=1.865 $Y2=3.235
cc_77 N_VDD_c_77_p N_A_M1003_g 0.00468827f $X=2.38 $Y=4.25 $X2=1.865 $Y2=3.235
cc_78 N_VDD_M1000_b N_A_c_124_n 0.0279802f $X=-0.045 $Y=2.425 $X2=0.45 $Y2=2.53
cc_79 N_VDD_c_79_p N_A_c_124_n 0.00606474f $X=0.605 $Y=4.287 $X2=0.45 $Y2=2.53
cc_80 N_VDD_c_80_p N_A_c_124_n 0.00337744f $X=0.69 $Y=2.955 $X2=0.45 $Y2=2.53
cc_81 N_VDD_c_77_p N_A_c_124_n 0.00468827f $X=2.38 $Y=4.25 $X2=0.45 $Y2=2.53
cc_82 N_VDD_M1000_b N_A_27_115#_M1009_g 0.0197604f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_83 N_VDD_c_80_p N_A_27_115#_M1009_g 0.00337744f $X=0.69 $Y=2.955 $X2=0.905
+ $Y2=3.235
cc_84 N_VDD_c_76_p N_A_27_115#_M1009_g 0.00606474f $X=2.355 $Y=4.287 $X2=0.905
+ $Y2=3.235
cc_85 N_VDD_c_77_p N_A_27_115#_M1009_g 0.00468827f $X=2.38 $Y=4.25 $X2=0.905
+ $Y2=3.235
cc_86 N_VDD_c_80_p N_A_27_115#_c_240_n 0.00176917f $X=0.69 $Y=2.955 $X2=0.845
+ $Y2=1.94
cc_87 N_VDD_M1000_b N_A_27_115#_c_245_n 0.0104815f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=2.955
cc_88 N_VDD_c_79_p N_A_27_115#_c_245_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=2.955
cc_89 N_VDD_c_77_p N_A_27_115#_c_245_n 0.00476261f $X=2.38 $Y=4.25 $X2=0.26
+ $Y2=2.955
cc_90 N_VDD_M1000_b N_A_238_89#_M1005_g 0.0192967f $X=-0.045 $Y=2.425 $X2=1.265
+ $Y2=3.235
cc_91 N_VDD_c_76_p N_A_238_89#_M1005_g 0.00606474f $X=2.355 $Y=4.287 $X2=1.265
+ $Y2=3.235
cc_92 N_VDD_c_77_p N_A_238_89#_M1005_g 0.00468827f $X=2.38 $Y=4.25 $X2=1.265
+ $Y2=3.235
cc_93 N_VDD_M1000_b N_A_238_89#_c_323_n 0.00559382f $X=-0.045 $Y=2.425 $X2=1.325
+ $Y2=2.285
cc_94 N_VDD_c_94_p N_A_238_89#_c_324_n 0.00811678f $X=2.44 $Y=2.955 $X2=2.785
+ $Y2=2.285
cc_95 N_VDD_M1000_b N_A_238_89#_c_327_n 0.00991954f $X=-0.045 $Y=2.425 $X2=2.87
+ $Y2=2.955
cc_96 N_VDD_c_96_p N_A_238_89#_c_327_n 0.00757793f $X=2.38 $Y=4.25 $X2=2.87
+ $Y2=2.955
cc_97 N_VDD_c_77_p N_A_238_89#_c_327_n 0.00476261f $X=2.38 $Y=4.25 $X2=2.87
+ $Y2=2.955
cc_98 N_VDD_M1000_b N_B_c_401_n 0.0139689f $X=-0.045 $Y=2.425 $X2=2.225 $Y2=2.53
cc_99 N_VDD_c_76_p N_B_c_401_n 0.00606474f $X=2.355 $Y=4.287 $X2=2.225 $Y2=2.53
cc_100 N_VDD_c_94_p N_B_c_401_n 0.00337744f $X=2.44 $Y=2.955 $X2=2.225 $Y2=2.53
cc_101 N_VDD_c_77_p N_B_c_401_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.225 $Y2=2.53
cc_102 N_VDD_M1000_b N_B_c_388_n 0.00535962f $X=-0.045 $Y=2.425 $X2=2.58
+ $Y2=2.455
cc_103 N_VDD_c_94_p N_B_c_388_n 0.00221017f $X=2.44 $Y=2.955 $X2=2.58 $Y2=2.455
cc_104 N_VDD_M1000_b N_B_c_389_n 0.00345657f $X=-0.045 $Y=2.425 $X2=2.3
+ $Y2=2.455
cc_105 N_VDD_M1000_b N_B_c_408_n 0.0183291f $X=-0.045 $Y=2.425 $X2=2.655
+ $Y2=2.53
cc_106 N_VDD_c_94_p N_B_c_408_n 0.00337744f $X=2.44 $Y=2.955 $X2=2.655 $Y2=2.53
cc_107 N_VDD_c_96_p N_B_c_408_n 0.00606474f $X=2.38 $Y=4.25 $X2=2.655 $Y2=2.53
cc_108 N_VDD_c_77_p N_B_c_408_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.655 $Y2=2.53
cc_109 N_VDD_M1000_b N_B_c_396_n 0.00423637f $X=-0.045 $Y=2.425 $X2=2.655
+ $Y2=2.455
cc_110 N_VDD_M1000_b N_Y_c_447_n 0.00313975f $X=-0.045 $Y=2.425 $X2=1.565
+ $Y2=3.635
cc_111 N_VDD_c_76_p N_Y_c_447_n 0.0149397f $X=2.355 $Y=4.287 $X2=1.565 $Y2=3.635
cc_112 N_VDD_c_77_p N_Y_c_447_n 0.00958198f $X=2.38 $Y=4.25 $X2=1.565 $Y2=3.635
cc_113 N_VDD_M1000_b Y 0.00321849f $X=-0.045 $Y=2.425 $X2=1.42 $Y2=1.655
cc_114 N_VDD_c_80_p N_Y_c_451_n 0.0045586f $X=0.69 $Y=2.955 $X2=1.425 $Y2=2.85
cc_115 N_A_c_123_n N_A_27_115#_M1009_g 0.0100216f $X=0.45 $Y=2.38 $X2=0.905
+ $Y2=3.235
cc_116 N_A_c_124_n N_A_27_115#_M1009_g 0.0231282f $X=0.45 $Y=2.53 $X2=0.905
+ $Y2=3.235
cc_117 N_A_c_136_n N_A_27_115#_c_237_n 0.00921346f $X=2.02 $Y=1 $X2=1.865
+ $Y2=1.235
cc_118 N_A_c_143_n N_A_27_115#_c_237_n 0.00289059f $X=2.107 $Y=1.625 $X2=1.865
+ $Y2=1.235
cc_119 N_A_c_123_n N_A_27_115#_c_240_n 0.0212638f $X=0.45 $Y=2.38 $X2=0.845
+ $Y2=1.94
cc_120 N_A_c_125_n N_A_27_115#_c_240_n 0.018362f $X=0.845 $Y=1.275 $X2=0.845
+ $Y2=1.94
cc_121 N_A_c_131_n N_A_27_115#_c_240_n 6.77205e-19 $X=0.845 $Y=1.37 $X2=0.845
+ $Y2=1.94
cc_122 A N_A_27_115#_c_240_n 5.38486e-19 $X=0.845 $Y=1.37 $X2=0.845 $Y2=1.94
cc_123 N_A_c_130_n N_A_27_115#_c_241_n 0.00513787f $X=1.865 $Y=1.955 $X2=1.765
+ $Y2=1.4
cc_124 N_A_c_136_n N_A_27_115#_c_241_n 0.00127901f $X=2.02 $Y=1 $X2=1.765
+ $Y2=1.4
cc_125 N_A_c_143_n N_A_27_115#_c_241_n 0.00175248f $X=2.107 $Y=1.625 $X2=1.765
+ $Y2=1.4
cc_126 N_A_c_115_n N_A_27_115#_c_242_n 0.0062242f $X=0.475 $Y=1.2 $X2=0.26
+ $Y2=0.755
cc_127 N_A_c_122_n N_A_27_115#_c_242_n 0.0233638f $X=0.45 $Y=1.275 $X2=0.26
+ $Y2=0.755
cc_128 N_A_c_131_n N_A_27_115#_c_242_n 0.00858616f $X=0.845 $Y=1.37 $X2=0.26
+ $Y2=0.755
cc_129 N_A_c_137_n N_A_27_115#_c_242_n 0.0128571f $X=0.93 $Y=1 $X2=0.26
+ $Y2=0.755
cc_130 A N_A_27_115#_c_242_n 0.00564707f $X=0.845 $Y=1.37 $X2=0.26 $Y2=0.755
cc_131 N_A_c_123_n N_A_27_115#_c_245_n 0.0208779f $X=0.45 $Y=2.38 $X2=0.26
+ $Y2=2.955
cc_132 N_A_c_124_n N_A_27_115#_c_245_n 0.00651153f $X=0.45 $Y=2.53 $X2=0.26
+ $Y2=2.955
cc_133 N_A_c_119_n N_A_27_115#_c_246_n 8.76512e-19 $X=0.71 $Y=1.275 $X2=1.68
+ $Y2=1.94
cc_134 N_A_c_123_n N_A_27_115#_c_246_n 0.019959f $X=0.45 $Y=2.38 $X2=1.68
+ $Y2=1.94
cc_135 N_A_c_124_n N_A_27_115#_c_246_n 0.00170478f $X=0.45 $Y=2.53 $X2=1.68
+ $Y2=1.94
cc_136 N_A_c_125_n N_A_27_115#_c_246_n 8.34298e-19 $X=0.845 $Y=1.275 $X2=1.68
+ $Y2=1.94
cc_137 N_A_c_130_n N_A_27_115#_c_246_n 0.00505743f $X=1.865 $Y=1.955 $X2=1.68
+ $Y2=1.94
cc_138 N_A_c_131_n N_A_27_115#_c_246_n 0.00683916f $X=0.845 $Y=1.37 $X2=1.68
+ $Y2=1.94
cc_139 N_A_c_133_n N_A_27_115#_c_246_n 0.0141647f $X=2.105 $Y=1.74 $X2=1.68
+ $Y2=1.94
cc_140 A N_A_27_115#_c_246_n 0.00489601f $X=0.845 $Y=1.37 $X2=1.68 $Y2=1.94
cc_141 N_A_c_130_n N_A_27_115#_c_247_n 4.6714e-19 $X=1.865 $Y=1.955 $X2=1.765
+ $Y2=1.4
cc_142 N_A_c_133_n N_A_27_115#_c_247_n 0.0130621f $X=2.105 $Y=1.74 $X2=1.765
+ $Y2=1.4
cc_143 N_A_c_136_n N_A_27_115#_c_247_n 0.00713168f $X=2.02 $Y=1 $X2=1.765
+ $Y2=1.4
cc_144 N_A_c_142_n N_A_27_115#_c_247_n 0.00336273f $X=2.105 $Y=1.74 $X2=1.765
+ $Y2=1.4
cc_145 N_A_c_143_n N_A_27_115#_c_247_n 0.00689669f $X=2.107 $Y=1.625 $X2=1.765
+ $Y2=1.4
cc_146 N_A_c_123_n N_A_238_89#_M1011_g 0.00462097f $X=0.45 $Y=2.38 $X2=1.265
+ $Y2=0.85
cc_147 N_A_c_126_n N_A_238_89#_M1011_g 0.0696135f $X=0.845 $Y=1.2 $X2=1.265
+ $Y2=0.85
cc_148 N_A_c_130_n N_A_238_89#_M1011_g 0.00442887f $X=1.865 $Y=1.955 $X2=1.265
+ $Y2=0.85
cc_149 N_A_c_131_n N_A_238_89#_M1011_g 0.00168579f $X=0.845 $Y=1.37 $X2=1.265
+ $Y2=0.85
cc_150 N_A_c_133_n N_A_238_89#_M1011_g 4.13594e-19 $X=2.105 $Y=1.74 $X2=1.265
+ $Y2=0.85
cc_151 N_A_c_134_n N_A_238_89#_M1011_g 8.13035e-19 $X=0.845 $Y=1.255 $X2=1.265
+ $Y2=0.85
cc_152 N_A_c_136_n N_A_238_89#_M1011_g 0.0089629f $X=2.02 $Y=1 $X2=1.265
+ $Y2=0.85
cc_153 A N_A_238_89#_M1011_g 9.48751e-19 $X=0.845 $Y=1.37 $X2=1.265 $Y2=0.85
cc_154 N_A_M1003_g N_A_238_89#_M1005_g 0.0320513f $X=1.865 $Y=3.235 $X2=1.265
+ $Y2=3.235
cc_155 N_A_M1003_g N_A_238_89#_c_323_n 0.0126871f $X=1.865 $Y=3.235 $X2=1.325
+ $Y2=2.285
cc_156 N_A_M1003_g N_A_238_89#_c_324_n 0.0182294f $X=1.865 $Y=3.235 $X2=2.785
+ $Y2=2.285
cc_157 N_A_c_130_n N_A_238_89#_c_324_n 0.00741834f $X=1.865 $Y=1.955 $X2=2.785
+ $Y2=2.285
cc_158 N_A_c_133_n N_A_238_89#_c_324_n 0.0257565f $X=2.105 $Y=1.74 $X2=2.785
+ $Y2=2.285
cc_159 N_A_c_142_n N_A_238_89#_c_324_n 0.00356792f $X=2.105 $Y=1.74 $X2=2.785
+ $Y2=2.285
cc_160 N_A_c_133_n N_A_238_89#_c_325_n 0.0107692f $X=2.105 $Y=1.74 $X2=2.87
+ $Y2=0.755
cc_161 N_A_c_136_n N_A_238_89#_c_325_n 0.0115282f $X=2.02 $Y=1 $X2=2.87
+ $Y2=0.755
cc_162 N_A_c_142_n N_A_238_89#_c_325_n 0.00537064f $X=2.105 $Y=1.74 $X2=2.87
+ $Y2=0.755
cc_163 N_A_c_136_n N_B_c_384_n 0.00416726f $X=2.02 $Y=1 $X2=2.225 $Y2=1.2
cc_164 N_A_c_143_n N_B_c_384_n 0.00173913f $X=2.107 $Y=1.625 $X2=2.225 $Y2=1.2
cc_165 N_A_M1003_g N_B_c_389_n 0.0980212f $X=1.865 $Y=3.235 $X2=2.3 $Y2=2.455
cc_166 N_A_c_130_n N_B_c_389_n 0.00900867f $X=1.865 $Y=1.955 $X2=2.3 $Y2=2.455
cc_167 N_A_c_136_n N_B_c_390_n 0.0012955f $X=2.02 $Y=1 $X2=2.655 $Y2=1.2
cc_168 N_A_M1003_g N_B_c_393_n 0.00331379f $X=1.865 $Y=3.235 $X2=2.655 $Y2=2.38
cc_169 N_A_c_130_n N_B_c_393_n 0.0193364f $X=1.865 $Y=1.955 $X2=2.655 $Y2=2.38
cc_170 N_A_c_133_n N_B_c_393_n 0.00361324f $X=2.105 $Y=1.74 $X2=2.655 $Y2=2.38
cc_171 N_A_c_142_n N_B_c_393_n 0.00298898f $X=2.105 $Y=1.74 $X2=2.655 $Y2=2.38
cc_172 N_A_c_130_n N_B_c_394_n 0.00684403f $X=1.865 $Y=1.955 $X2=2.655 $Y2=1.382
cc_173 N_A_c_133_n N_B_c_394_n 0.00265313f $X=2.105 $Y=1.74 $X2=2.655 $Y2=1.382
cc_174 N_A_c_142_n N_B_c_394_n 0.00102425f $X=2.105 $Y=1.74 $X2=2.655 $Y2=1.382
cc_175 N_A_c_143_n N_B_c_394_n 0.00355806f $X=2.107 $Y=1.625 $X2=2.655 $Y2=1.382
cc_176 N_A_c_143_n N_B_c_397_n 0.0041324f $X=2.107 $Y=1.625 $X2=2.53 $Y2=1.37
cc_177 N_A_c_143_n B 0.020637f $X=2.107 $Y=1.625 $X2=2.53 $Y2=1.4
cc_178 N_A_c_136_n N_Y_M1011_d 0.0052569f $X=2.02 $Y=1 $X2=1.34 $Y2=0.575
cc_179 N_A_c_131_n N_Y_c_441_n 0.00551701f $X=0.845 $Y=1.37 $X2=1.425 $Y2=1.37
cc_180 N_A_c_134_n N_Y_c_441_n 0.00530076f $X=0.845 $Y=1.255 $X2=1.425 $Y2=1.37
cc_181 N_A_c_136_n N_Y_c_441_n 0.014779f $X=2.02 $Y=1 $X2=1.425 $Y2=1.37
cc_182 A N_Y_c_441_n 9.01697e-19 $X=0.845 $Y=1.37 $X2=1.425 $Y2=1.37
cc_183 N_A_c_143_n N_Y_c_441_n 0.00503144f $X=2.107 $Y=1.625 $X2=1.425 $Y2=1.37
cc_184 N_A_c_126_n N_Y_c_442_n 5.92936e-19 $X=0.845 $Y=1.2 $X2=1.425 $Y2=0.755
cc_185 N_A_c_136_n N_Y_c_442_n 0.014597f $X=2.02 $Y=1 $X2=1.425 $Y2=0.755
cc_186 N_A_c_125_n Y 3.61257e-19 $X=0.845 $Y=1.275 $X2=1.42 $Y2=1.655
cc_187 N_A_c_130_n Y 0.00702394f $X=1.865 $Y=1.955 $X2=1.42 $Y2=1.655
cc_188 N_A_c_131_n Y 0.00234899f $X=0.845 $Y=1.37 $X2=1.42 $Y2=1.655
cc_189 N_A_c_133_n Y 6.59307e-19 $X=2.105 $Y=1.74 $X2=1.42 $Y2=1.655
cc_190 N_A_c_142_n Y 0.0130548f $X=2.105 $Y=1.74 $X2=1.42 $Y2=1.655
cc_191 N_A_c_143_n Y 0.00703362f $X=2.107 $Y=1.625 $X2=1.42 $Y2=1.655
cc_192 N_A_c_125_n N_Y_c_446_n 2.49214e-19 $X=0.845 $Y=1.275 $X2=1.425 $Y2=1.37
cc_193 N_A_c_131_n N_Y_c_446_n 0.00145163f $X=0.845 $Y=1.37 $X2=1.425 $Y2=1.37
cc_194 N_A_c_136_n N_Y_c_446_n 0.0259322f $X=2.02 $Y=1 $X2=1.425 $Y2=1.37
cc_195 A N_Y_c_446_n 0.0172747f $X=0.845 $Y=1.37 $X2=1.425 $Y2=1.37
cc_196 N_A_c_143_n N_Y_c_446_n 0.0130404f $X=2.107 $Y=1.625 $X2=1.425 $Y2=1.37
cc_197 N_A_c_136_n A_196_115# 0.0106358f $X=2.02 $Y=1 $X2=0.98 $Y2=0.575
cc_198 N_A_c_136_n A_388_115# 0.00450984f $X=2.02 $Y=1 $X2=1.94 $Y2=0.575
cc_199 N_A_c_143_n A_388_115# 4.72742e-19 $X=2.107 $Y=1.625 $X2=1.94 $Y2=0.575
cc_200 N_A_27_115#_c_237_n N_A_238_89#_M1011_g 0.0180699f $X=1.865 $Y=1.235
+ $X2=1.265 $Y2=0.85
cc_201 N_A_27_115#_c_240_n N_A_238_89#_M1011_g 0.067895f $X=0.845 $Y=1.94
+ $X2=1.265 $Y2=0.85
cc_202 N_A_27_115#_c_241_n N_A_238_89#_M1011_g 0.0145931f $X=1.765 $Y=1.4
+ $X2=1.265 $Y2=0.85
cc_203 N_A_27_115#_c_246_n N_A_238_89#_M1011_g 0.0144815f $X=1.68 $Y=1.94
+ $X2=1.265 $Y2=0.85
cc_204 N_A_27_115#_c_247_n N_A_238_89#_M1011_g 0.00769245f $X=1.765 $Y=1.4
+ $X2=1.265 $Y2=0.85
cc_205 N_A_27_115#_M1009_g N_A_238_89#_c_323_n 0.067895f $X=0.905 $Y=3.235
+ $X2=1.325 $Y2=2.285
cc_206 N_A_27_115#_c_246_n N_A_238_89#_c_323_n 0.002291f $X=1.68 $Y=1.94
+ $X2=1.325 $Y2=2.285
cc_207 N_A_27_115#_M1009_g N_A_238_89#_c_324_n 0.00444529f $X=0.905 $Y=3.235
+ $X2=2.785 $Y2=2.285
cc_208 N_A_27_115#_c_241_n N_A_238_89#_c_324_n 6.35071e-19 $X=1.765 $Y=1.4
+ $X2=2.785 $Y2=2.285
cc_209 N_A_27_115#_c_246_n N_A_238_89#_c_324_n 0.0495257f $X=1.68 $Y=1.94
+ $X2=2.785 $Y2=2.285
cc_210 N_A_27_115#_c_237_n N_B_c_384_n 0.02878f $X=1.865 $Y=1.235 $X2=2.225
+ $Y2=1.2
cc_211 N_A_27_115#_c_241_n N_B_c_394_n 0.0337502f $X=1.765 $Y=1.4 $X2=2.655
+ $Y2=1.382
cc_212 N_A_27_115#_c_247_n N_B_c_394_n 9.96331e-19 $X=1.765 $Y=1.4 $X2=2.655
+ $Y2=1.382
cc_213 N_A_27_115#_c_241_n N_B_c_397_n 0.0012687f $X=1.765 $Y=1.4 $X2=2.53
+ $Y2=1.37
cc_214 N_A_27_115#_c_247_n N_B_c_397_n 0.00326486f $X=1.765 $Y=1.4 $X2=2.53
+ $Y2=1.37
cc_215 N_A_27_115#_c_237_n N_Y_c_441_n 0.0050539f $X=1.865 $Y=1.235 $X2=1.425
+ $Y2=1.37
cc_216 N_A_27_115#_c_241_n N_Y_c_441_n 0.00141648f $X=1.765 $Y=1.4 $X2=1.425
+ $Y2=1.37
cc_217 N_A_27_115#_c_246_n N_Y_c_441_n 0.00508766f $X=1.68 $Y=1.94 $X2=1.425
+ $Y2=1.37
cc_218 N_A_27_115#_c_247_n N_Y_c_441_n 0.0137932f $X=1.765 $Y=1.4 $X2=1.425
+ $Y2=1.37
cc_219 N_A_27_115#_M1009_g N_Y_c_475_n 7.92921e-19 $X=0.905 $Y=3.235 $X2=1.565
+ $Y2=2.965
cc_220 N_A_27_115#_c_237_n N_Y_c_442_n 0.00244041f $X=1.865 $Y=1.235 $X2=1.425
+ $Y2=0.755
cc_221 N_A_27_115#_c_241_n N_Y_c_442_n 0.00181308f $X=1.765 $Y=1.4 $X2=1.425
+ $Y2=0.755
cc_222 N_A_27_115#_c_247_n N_Y_c_442_n 0.00192723f $X=1.765 $Y=1.4 $X2=1.425
+ $Y2=0.755
cc_223 N_A_27_115#_M1009_g Y 0.00191867f $X=0.905 $Y=3.235 $X2=1.42 $Y2=1.655
cc_224 N_A_27_115#_c_240_n Y 7.98026e-19 $X=0.845 $Y=1.94 $X2=1.42 $Y2=1.655
cc_225 N_A_27_115#_c_241_n Y 5.37513e-19 $X=1.765 $Y=1.4 $X2=1.42 $Y2=1.655
cc_226 N_A_27_115#_c_246_n Y 0.0158271f $X=1.68 $Y=1.94 $X2=1.42 $Y2=1.655
cc_227 N_A_27_115#_c_247_n Y 0.0108798f $X=1.765 $Y=1.4 $X2=1.42 $Y2=1.655
cc_228 N_A_27_115#_c_241_n N_Y_c_446_n 0.00177952f $X=1.765 $Y=1.4 $X2=1.425
+ $Y2=1.37
cc_229 N_A_27_115#_c_246_n N_Y_c_446_n 0.00426863f $X=1.68 $Y=1.94 $X2=1.425
+ $Y2=1.37
cc_230 N_A_27_115#_c_247_n N_Y_c_446_n 0.00314875f $X=1.765 $Y=1.4 $X2=1.425
+ $Y2=1.37
cc_231 N_A_27_115#_M1009_g N_Y_c_451_n 0.00108503f $X=0.905 $Y=3.235 $X2=1.425
+ $Y2=2.85
cc_232 N_A_238_89#_c_324_n N_B_c_389_n 0.0131927f $X=2.785 $Y=2.285 $X2=2.3
+ $Y2=2.455
cc_233 N_A_238_89#_c_325_n N_B_c_390_n 0.0364201f $X=2.87 $Y=0.755 $X2=2.655
+ $Y2=1.2
cc_234 N_A_238_89#_c_324_n N_B_c_393_n 0.0200313f $X=2.785 $Y=2.285 $X2=2.655
+ $Y2=2.38
cc_235 N_A_238_89#_c_327_n N_B_c_393_n 0.0137951f $X=2.87 $Y=2.955 $X2=2.655
+ $Y2=2.38
cc_236 N_A_238_89#_c_324_n N_B_c_394_n 0.00185828f $X=2.785 $Y=2.285 $X2=2.655
+ $Y2=1.382
cc_237 N_A_238_89#_c_324_n N_B_c_397_n 0.00451293f $X=2.785 $Y=2.285 $X2=2.53
+ $Y2=1.37
cc_238 N_A_238_89#_c_325_n N_B_c_397_n 0.0211625f $X=2.87 $Y=0.755 $X2=2.53
+ $Y2=1.37
cc_239 N_A_238_89#_c_325_n B 0.00784554f $X=2.87 $Y=0.755 $X2=2.53 $Y2=1.4
cc_240 N_A_238_89#_M1011_g N_Y_c_441_n 0.00793259f $X=1.265 $Y=0.85 $X2=1.425
+ $Y2=1.37
cc_241 N_A_238_89#_M1005_g N_Y_c_475_n 0.0034761f $X=1.265 $Y=3.235 $X2=1.565
+ $Y2=2.965
cc_242 N_A_238_89#_c_323_n N_Y_c_475_n 0.00170549f $X=1.325 $Y=2.285 $X2=1.565
+ $Y2=2.965
cc_243 N_A_238_89#_c_324_n N_Y_c_475_n 0.015078f $X=2.785 $Y=2.285 $X2=1.565
+ $Y2=2.965
cc_244 N_A_238_89#_M1011_g N_Y_c_442_n 0.00333621f $X=1.265 $Y=0.85 $X2=1.425
+ $Y2=0.755
cc_245 N_A_238_89#_M1011_g Y 0.00978463f $X=1.265 $Y=0.85 $X2=1.42 $Y2=1.655
cc_246 N_A_238_89#_M1005_g Y 0.00464698f $X=1.265 $Y=3.235 $X2=1.42 $Y2=1.655
cc_247 N_A_238_89#_c_323_n Y 0.00651733f $X=1.325 $Y=2.285 $X2=1.42 $Y2=1.655
cc_248 N_A_238_89#_c_324_n Y 0.0162812f $X=2.785 $Y=2.285 $X2=1.42 $Y2=1.655
cc_249 N_A_238_89#_M1011_g N_Y_c_446_n 0.00296721f $X=1.265 $Y=0.85 $X2=1.425
+ $Y2=1.37
cc_250 N_A_238_89#_M1005_g N_Y_c_451_n 0.00624758f $X=1.265 $Y=3.235 $X2=1.425
+ $Y2=2.85
cc_251 N_A_238_89#_c_324_n N_Y_c_451_n 0.00233457f $X=2.785 $Y=2.285 $X2=1.425
+ $Y2=2.85
