magic
tech sky130A
magscale 1 2
timestamp 1612372269
<< nwell >>
rect -9 529 199 1119
<< nmoslvt >>
rect 80 115 110 445
<< pmos >>
rect 80 713 110 965
<< ndiff >>
rect 27 335 80 445
rect 27 131 35 335
rect 69 131 80 335
rect 27 115 80 131
rect 110 335 163 445
rect 110 131 121 335
rect 155 131 163 335
rect 110 115 163 131
<< pdiff >>
rect 27 949 80 965
rect 27 745 35 949
rect 69 745 80 949
rect 27 713 80 745
rect 110 949 163 965
rect 110 745 121 949
rect 155 745 163 949
rect 110 713 163 745
<< ndiffc >>
rect 35 131 69 335
rect 121 131 155 335
<< pdiffc >>
rect 35 745 69 949
rect 121 745 155 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1049 85 1083
<< poly >>
rect 80 965 110 991
rect 80 445 110 713
rect 80 80 110 115
<< locali >>
rect 0 1089 198 1110
rect 0 1049 51 1089
rect 85 1049 198 1089
rect 35 949 69 1049
rect 35 729 69 745
rect 121 949 155 1049
rect 121 729 155 745
rect 35 335 69 351
rect 35 61 69 131
rect 121 335 155 351
rect 121 61 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1089 198 1110
rect 0 1055 51 1089
rect 85 1055 198 1089
rect 0 1049 198 1055
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
