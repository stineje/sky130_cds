magic
tech sky130A
magscale 1 2
timestamp 1606864593
<< checkpaint >>
rect -1209 -1243 2569 2575
<< nwell >>
rect -9 581 1456 1341
<< nmos >>
rect 85 115 115 315
rect 171 115 201 315
rect 243 115 273 315
rect 363 115 393 315
rect 435 115 465 315
rect 521 115 551 315
rect 593 115 623 315
rect 713 115 743 315
rect 785 115 815 315
rect 871 115 901 315
rect 1061 115 1091 315
rect 1251 115 1281 315
rect 1337 115 1367 315
<< pmoshvt >>
rect 85 617 115 1217
rect 171 617 201 1217
rect 243 617 273 1217
rect 363 617 393 1217
rect 435 617 465 1217
rect 521 617 551 1217
rect 593 617 623 1217
rect 713 617 743 1217
rect 785 617 815 1217
rect 871 617 901 1217
rect 1061 617 1091 1217
rect 1251 617 1281 1217
rect 1337 617 1367 1217
<< ndiff >>
rect 32 267 85 315
rect 32 131 40 267
rect 74 131 85 267
rect 32 115 85 131
rect 115 267 171 315
rect 115 131 126 267
rect 160 131 171 267
rect 115 115 171 131
rect 201 115 243 315
rect 273 267 363 315
rect 273 131 284 267
rect 352 131 363 267
rect 273 115 363 131
rect 393 115 435 315
rect 465 199 521 315
rect 465 131 476 199
rect 510 131 521 199
rect 465 115 521 131
rect 551 115 593 315
rect 623 267 713 315
rect 623 131 634 267
rect 702 131 713 267
rect 623 115 713 131
rect 743 115 785 315
rect 815 267 871 315
rect 815 131 826 267
rect 860 131 871 267
rect 815 115 871 131
rect 901 267 954 315
rect 901 131 912 267
rect 946 131 954 267
rect 901 115 954 131
rect 1008 267 1061 315
rect 1008 131 1016 267
rect 1050 131 1061 267
rect 1008 115 1061 131
rect 1091 267 1144 315
rect 1091 131 1102 267
rect 1136 131 1144 267
rect 1091 115 1144 131
rect 1198 267 1251 315
rect 1198 131 1206 267
rect 1240 131 1251 267
rect 1198 115 1251 131
rect 1281 267 1337 315
rect 1281 131 1292 267
rect 1326 131 1337 267
rect 1281 115 1337 131
rect 1367 267 1420 315
rect 1367 131 1378 267
rect 1412 131 1420 267
rect 1367 115 1420 131
<< pdiff >>
rect 32 1201 85 1217
rect 32 657 40 1201
rect 74 657 85 1201
rect 32 617 85 657
rect 115 1201 171 1217
rect 115 725 126 1201
rect 160 725 171 1201
rect 115 617 171 725
rect 201 617 243 1217
rect 273 1201 363 1217
rect 273 657 284 1201
rect 352 657 363 1201
rect 273 617 363 657
rect 393 617 435 1217
rect 465 1201 521 1217
rect 465 725 476 1201
rect 510 725 521 1201
rect 465 617 521 725
rect 551 617 593 1217
rect 623 1201 713 1217
rect 623 657 634 1201
rect 702 657 713 1201
rect 623 617 713 657
rect 743 617 785 1217
rect 815 1201 871 1217
rect 815 657 826 1201
rect 860 657 871 1201
rect 815 617 871 657
rect 901 1201 954 1217
rect 901 657 912 1201
rect 946 657 954 1201
rect 901 617 954 657
rect 1008 1201 1061 1217
rect 1008 725 1016 1201
rect 1050 725 1061 1201
rect 1008 617 1061 725
rect 1091 1201 1144 1217
rect 1091 657 1102 1201
rect 1136 657 1144 1201
rect 1091 617 1144 657
rect 1198 1201 1251 1217
rect 1198 657 1206 1201
rect 1240 657 1251 1201
rect 1198 617 1251 657
rect 1281 1201 1337 1217
rect 1281 657 1292 1201
rect 1326 657 1337 1201
rect 1281 617 1337 657
rect 1367 1201 1420 1217
rect 1367 657 1378 1201
rect 1412 657 1420 1201
rect 1367 617 1420 657
<< ndiffc >>
rect 40 131 74 267
rect 126 131 160 267
rect 284 131 352 267
rect 476 131 510 199
rect 634 131 702 267
rect 826 131 860 267
rect 912 131 946 267
rect 1016 131 1050 267
rect 1102 131 1136 267
rect 1206 131 1240 267
rect 1292 131 1326 267
rect 1378 131 1412 267
<< pdiffc >>
rect 40 657 74 1201
rect 126 725 160 1201
rect 284 657 352 1201
rect 476 725 510 1201
rect 634 657 702 1201
rect 826 657 860 1201
rect 912 657 946 1201
rect 1016 725 1050 1201
rect 1102 657 1136 1201
rect 1206 657 1240 1201
rect 1292 657 1326 1201
rect 1378 657 1412 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
rect 979 27 1003 61
rect 1037 27 1061 61
rect 1115 27 1139 61
rect 1173 27 1197 61
rect 1251 27 1275 61
rect 1309 27 1333 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
rect 707 1271 731 1305
rect 765 1271 789 1305
rect 843 1271 867 1305
rect 901 1271 925 1305
rect 979 1271 1003 1305
rect 1037 1271 1061 1305
rect 1115 1271 1139 1305
rect 1173 1271 1197 1305
rect 1251 1271 1275 1305
rect 1309 1271 1333 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
rect 1003 27 1037 61
rect 1139 27 1173 61
rect 1275 27 1309 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
rect 731 1271 765 1305
rect 867 1271 901 1305
rect 1003 1271 1037 1305
rect 1139 1271 1173 1305
rect 1275 1271 1309 1305
<< poly >>
rect 85 1217 115 1243
rect 171 1217 201 1243
rect 243 1217 273 1243
rect 363 1217 393 1243
rect 435 1217 465 1243
rect 521 1217 551 1243
rect 593 1217 623 1243
rect 713 1217 743 1243
rect 785 1217 815 1243
rect 871 1217 901 1243
rect 1061 1217 1091 1243
rect 1251 1217 1281 1243
rect 1337 1217 1367 1243
rect 85 586 115 617
rect 75 570 129 586
rect 75 536 85 570
rect 119 536 129 570
rect 75 520 129 536
rect 75 374 105 520
rect 171 477 201 617
rect 243 586 273 617
rect 243 570 297 586
rect 243 536 253 570
rect 287 536 297 570
rect 243 520 297 536
rect 171 461 225 477
rect 363 475 393 617
rect 435 580 465 617
rect 521 580 551 617
rect 435 570 551 580
rect 435 536 467 570
rect 501 536 551 570
rect 435 526 551 536
rect 593 475 623 617
rect 713 586 743 617
rect 689 570 743 586
rect 689 536 699 570
rect 733 536 743 570
rect 689 520 743 536
rect 171 427 181 461
rect 215 427 225 461
rect 171 411 225 427
rect 267 445 719 475
rect 75 344 115 374
rect 85 315 115 344
rect 171 315 201 411
rect 267 367 297 445
rect 689 403 719 445
rect 785 471 815 617
rect 871 586 901 617
rect 871 570 942 586
rect 871 556 898 570
rect 882 536 898 556
rect 932 536 942 570
rect 882 520 942 536
rect 785 455 839 471
rect 785 421 795 455
rect 829 421 839 455
rect 785 405 839 421
rect 243 337 297 367
rect 339 387 393 403
rect 339 353 349 387
rect 383 353 393 387
rect 339 337 393 353
rect 243 315 273 337
rect 363 315 393 337
rect 435 387 551 397
rect 435 353 467 387
rect 501 353 551 387
rect 435 343 551 353
rect 435 315 465 343
rect 521 315 551 343
rect 593 387 647 403
rect 593 353 603 387
rect 637 353 647 387
rect 593 337 647 353
rect 689 387 743 403
rect 689 353 699 387
rect 733 353 743 387
rect 689 337 743 353
rect 593 315 623 337
rect 713 315 743 337
rect 785 315 815 405
rect 882 367 912 520
rect 1061 403 1091 617
rect 1251 601 1281 617
rect 1241 571 1281 601
rect 1241 471 1271 571
rect 1337 512 1367 617
rect 1216 455 1271 471
rect 1216 421 1226 455
rect 1260 421 1271 455
rect 1313 496 1367 512
rect 1313 462 1323 496
rect 1357 462 1367 496
rect 1313 446 1367 462
rect 1216 405 1271 421
rect 871 337 912 367
rect 1008 387 1091 403
rect 1008 353 1018 387
rect 1052 353 1091 387
rect 1008 337 1091 353
rect 871 315 901 337
rect 1061 315 1091 337
rect 1241 360 1271 405
rect 1241 330 1281 360
rect 1251 315 1281 330
rect 1337 315 1367 446
rect 85 89 115 115
rect 171 89 201 115
rect 243 89 273 115
rect 363 89 393 115
rect 435 89 465 115
rect 521 89 551 115
rect 593 89 623 115
rect 713 89 743 115
rect 785 89 815 115
rect 871 89 901 115
rect 1061 89 1091 115
rect 1251 89 1281 115
rect 1337 89 1367 115
<< polycont >>
rect 85 536 119 570
rect 253 536 287 570
rect 467 536 501 570
rect 699 536 733 570
rect 181 427 215 461
rect 898 536 932 570
rect 795 421 829 455
rect 349 353 383 387
rect 467 353 501 387
rect 603 353 637 387
rect 699 353 733 387
rect 1226 421 1260 455
rect 1323 462 1357 496
rect 1018 353 1052 387
<< locali >>
rect 0 1311 1452 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 595 1311
rect 629 1271 731 1311
rect 765 1271 867 1311
rect 901 1271 1003 1311
rect 1037 1271 1139 1311
rect 1173 1271 1275 1311
rect 1309 1271 1452 1311
rect 40 1201 74 1217
rect 17 657 40 669
rect 126 1201 160 1271
rect 126 709 160 725
rect 284 1201 352 1217
rect 17 628 74 657
rect 476 1201 510 1271
rect 476 709 510 725
rect 634 1201 702 1217
rect 352 657 355 675
rect 284 654 355 657
rect 634 654 702 657
rect 17 387 51 628
rect 108 620 355 654
rect 535 620 702 654
rect 826 1201 860 1271
rect 826 641 860 657
rect 912 1201 946 1217
rect 1016 1201 1050 1271
rect 1016 709 1050 725
rect 1102 1201 1136 1217
rect 912 654 946 657
rect 912 620 1000 654
rect 108 586 142 620
rect 85 570 142 586
rect 119 536 142 570
rect 85 520 142 536
rect 17 353 40 387
rect 17 332 74 353
rect 108 370 142 520
rect 253 570 287 586
rect 253 535 287 536
rect 467 570 501 586
rect 287 501 383 535
rect 181 461 215 477
rect 181 411 215 427
rect 349 387 383 501
rect 467 387 501 536
rect 108 336 315 370
rect 349 337 383 353
rect 467 337 501 353
rect 535 387 569 620
rect 699 570 733 586
rect 699 535 733 536
rect 40 267 74 332
rect 281 283 315 336
rect 535 303 569 353
rect 603 501 699 535
rect 898 570 932 586
rect 898 535 932 536
rect 603 387 637 501
rect 966 455 1000 620
rect 779 421 795 455
rect 829 421 845 455
rect 912 421 1000 455
rect 1102 455 1136 657
rect 1206 1201 1240 1217
rect 1206 609 1240 657
rect 1292 1201 1326 1271
rect 1292 641 1326 657
rect 1378 1201 1412 1217
rect 1412 649 1435 666
rect 1378 632 1435 649
rect 1206 570 1240 575
rect 1206 536 1357 570
rect 1323 496 1357 536
rect 1102 421 1226 455
rect 1260 421 1276 455
rect 912 387 946 421
rect 683 353 699 387
rect 733 353 946 387
rect 1002 353 1018 387
rect 1052 353 1068 387
rect 603 337 637 353
rect 40 115 74 131
rect 126 267 160 283
rect 281 267 352 283
rect 535 269 702 303
rect 281 249 284 267
rect 126 61 160 131
rect 634 267 702 269
rect 284 115 352 131
rect 476 199 510 215
rect 476 61 510 131
rect 634 115 702 131
rect 826 267 860 283
rect 826 61 860 131
rect 912 267 946 353
rect 912 115 946 131
rect 1016 267 1050 283
rect 1016 61 1050 131
rect 1102 267 1136 421
rect 1323 387 1357 462
rect 1102 115 1136 131
rect 1206 353 1357 387
rect 1206 267 1240 353
rect 1401 322 1435 632
rect 1378 286 1435 322
rect 1206 115 1240 131
rect 1292 267 1326 283
rect 1292 61 1326 131
rect 1378 267 1412 286
rect 1378 115 1412 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1003 61
rect 1037 21 1139 61
rect 1173 21 1275 61
rect 1309 21 1452 61
rect 0 0 1452 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 595 1305 629 1311
rect 595 1277 629 1305
rect 731 1305 765 1311
rect 731 1277 765 1305
rect 867 1305 901 1311
rect 867 1277 901 1305
rect 1003 1305 1037 1311
rect 1003 1277 1037 1305
rect 1139 1305 1173 1311
rect 1139 1277 1173 1305
rect 1275 1305 1309 1311
rect 1275 1277 1309 1305
rect 40 353 74 387
rect 253 501 287 535
rect 181 427 215 461
rect 449 353 467 387
rect 467 353 483 387
rect 535 353 569 387
rect 699 501 733 535
rect 898 501 932 535
rect 795 421 829 455
rect 1378 657 1412 683
rect 1378 649 1412 657
rect 1206 575 1240 609
rect 1226 421 1260 455
rect 1018 353 1052 387
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
rect 1003 27 1037 55
rect 1003 21 1037 27
rect 1139 27 1173 55
rect 1139 21 1173 27
rect 1275 27 1309 55
rect 1275 21 1309 27
<< metal1 >>
rect 0 1311 1452 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 595 1311
rect 629 1277 731 1311
rect 765 1277 867 1311
rect 901 1277 1003 1311
rect 1037 1277 1139 1311
rect 1173 1277 1275 1311
rect 1309 1277 1452 1311
rect 0 1271 1452 1277
rect 1366 683 1424 689
rect 1343 649 1378 683
rect 1412 649 1424 683
rect 1366 643 1424 649
rect 1194 609 1252 615
rect 1172 575 1206 609
rect 1240 575 1252 609
rect 1194 569 1252 575
rect 241 535 299 541
rect 687 535 745 541
rect 886 535 944 541
rect 241 501 253 535
rect 287 501 699 535
rect 733 501 898 535
rect 932 501 944 535
rect 241 495 299 501
rect 687 495 745 501
rect 886 495 944 501
rect 169 461 227 467
rect 169 427 181 461
rect 215 427 249 461
rect 783 455 841 461
rect 1214 455 1272 461
rect 169 421 227 427
rect 783 421 795 455
rect 829 421 1226 455
rect 1260 421 1272 455
rect 783 415 841 421
rect 1214 415 1272 421
rect 28 387 86 393
rect 437 387 495 393
rect 28 353 40 387
rect 74 353 449 387
rect 483 353 495 387
rect 28 347 86 353
rect 437 347 495 353
rect 523 387 581 393
rect 1006 387 1064 393
rect 523 353 535 387
rect 569 353 1018 387
rect 1052 353 1064 387
rect 523 347 581 353
rect 1006 347 1064 353
rect 0 55 1452 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1003 55
rect 1037 21 1139 55
rect 1173 21 1275 55
rect 1309 21 1452 55
rect 0 0 1452 21
<< labels >>
rlabel metal1 198 444 198 444 1 D
port 1 n
rlabel metal1 915 518 915 518 1 CK
port 3 n
rlabel metal1 1395 666 1395 666 1 Q
port 4 n
rlabel metal1 1224 592 1224 592 1 QN
port 2 n
rlabel viali 68 49 68 49 1 gnd
rlabel viali 68 1285 68 1285 1 vdd
<< end >>
