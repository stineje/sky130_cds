* File: sky130_osu_sc_15T_ls__and2_8.spice
* Created: Fri Nov 12 14:53:56 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__and2_8.pex.spice"
.subckt sky130_osu_sc_15T_ls__and2_8  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1007 A_110_115# N_A_M1007_g N_A_27_115#_M1007_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75004.1 A=0.111 P=1.78 MULT=1
MM1003 N_GND_M1003_d N_B_M1003_g A_110_115# N_GND_M1007_b NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.0777 PD=1.09 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1003_d N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.1 SB=75003.2 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1001_d N_A_27_115#_M1008_g N_GND_M1008_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_A_27_115#_M1009_g N_GND_M1008_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1009_d N_A_27_115#_M1012_g N_GND_M1012_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.3 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_A_27_115#_M1013_g N_GND_M1012_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1013_d N_A_27_115#_M1014_g N_GND_M1014_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1016_d N_A_27_115#_M1016_g N_GND_M1014_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1016_d N_A_27_115#_M1018_g N_GND_M1018_s N_GND_M1007_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75004.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75004.1 A=0.3 P=4.3 MULT=1
MM1010 N_VDD_M1010_d N_B_M1010_g N_A_27_115#_M1000_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75003.6 A=0.3 P=4.3 MULT=1
MM1002 N_Y_M1002_d N_A_27_115#_M1002_g N_VDD_M1010_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75003.2 A=0.3 P=4.3 MULT=1
MM1004 N_Y_M1002_d N_A_27_115#_M1004_g N_VDD_M1004_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001.5 SB=75002.8 A=0.3 P=4.3 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_VDD_M1004_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001.9 SB=75002.3 A=0.3 P=4.3 MULT=1
MM1006 N_Y_M1005_d N_A_27_115#_M1006_g N_VDD_M1006_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.3 SB=75001.9 A=0.3 P=4.3 MULT=1
MM1011 N_Y_M1011_d N_A_27_115#_M1011_g N_VDD_M1006_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.8 SB=75001.5 A=0.3 P=4.3 MULT=1
MM1015 N_Y_M1011_d N_A_27_115#_M1015_g N_VDD_M1015_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1017 N_Y_M1017_d N_A_27_115#_M1017_g N_VDD_M1015_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.6 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1019 N_Y_M1017_d N_A_27_115#_M1019_g N_VDD_M1019_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75004.1 SB=75000.2 A=0.3 P=4.3 MULT=1
DX20_noxref N_GND_M1007_b N_VDD_M1000_b NWDIODE A=14.7352 P=15.89
pX21_noxref noxref_8 A A PROBETYPE=1
pX22_noxref noxref_9 B B PROBETYPE=1
pX23_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__and2_8.pxi.spice"
*
.ends
*
*
