* File: sky130_osu_sc_18T_ms__and2_2.pxi.spice
* Created: Thu Oct 29 17:27:21 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__AND2_2%GND N_GND_M1002_d N_GND_M1006_s N_GND_M1004_b
+ N_GND_c_7_p N_GND_c_21_p N_GND_c_2_p N_GND_c_16_p GND N_GND_c_3_p
+ PM_SKY130_OSU_SC_18T_MS__AND2_2%GND
x_PM_SKY130_OSU_SC_18T_MS__AND2_2%VDD N_VDD_M1005_s N_VDD_M1000_d N_VDD_M1007_s
+ N_VDD_M1005_b N_VDD_c_46_p N_VDD_c_47_p N_VDD_c_58_p N_VDD_c_70_p N_VDD_c_65_p
+ VDD N_VDD_c_48_p PM_SKY130_OSU_SC_18T_MS__AND2_2%VDD
x_PM_SKY130_OSU_SC_18T_MS__AND2_2%A N_A_M1004_g N_A_M1005_g A N_A_c_84_n
+ N_A_c_85_n PM_SKY130_OSU_SC_18T_MS__AND2_2%A
x_PM_SKY130_OSU_SC_18T_MS__AND2_2%B N_B_M1002_g N_B_M1000_g B N_B_c_119_n
+ N_B_c_120_n PM_SKY130_OSU_SC_18T_MS__AND2_2%B
x_PM_SKY130_OSU_SC_18T_MS__AND2_2%A_27_115# N_A_27_115#_M1004_s
+ N_A_27_115#_M1005_d N_A_27_115#_M1001_g N_A_27_115#_c_175_n
+ N_A_27_115#_M1003_g N_A_27_115#_c_158_n N_A_27_115#_c_159_n
+ N_A_27_115#_M1006_g N_A_27_115#_c_180_n N_A_27_115#_M1007_g
+ N_A_27_115#_c_164_n N_A_27_115#_c_165_n N_A_27_115#_c_168_n
+ N_A_27_115#_c_169_n N_A_27_115#_c_186_n N_A_27_115#_c_170_n
+ N_A_27_115#_c_172_n N_A_27_115#_c_173_n N_A_27_115#_c_174_n
+ N_A_27_115#_c_202_n PM_SKY130_OSU_SC_18T_MS__AND2_2%A_27_115#
x_PM_SKY130_OSU_SC_18T_MS__AND2_2%Y N_Y_M1001_d N_Y_M1003_d Y N_Y_c_242_n
+ N_Y_c_245_n N_Y_c_246_n N_Y_c_247_n PM_SKY130_OSU_SC_18T_MS__AND2_2%Y
cc_1 N_GND_M1004_b N_A_M1004_g 0.0806078f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1004_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1004_g 0.00468827f $X=1.7 $Y=0.17 $X2=0.475 $Y2=1.075
cc_4 N_GND_M1004_b N_A_c_84_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.765
cc_5 N_GND_M1004_b N_A_c_85_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_6 N_GND_M1004_b N_B_M1002_g 0.0460664f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_7 N_GND_c_7_p N_B_M1002_g 0.00376152f $X=1.05 $Y=0.825 $X2=0.835 $Y2=1.075
cc_8 N_GND_c_2_p N_B_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=1.075
cc_9 N_GND_c_3_p N_B_M1002_g 0.00468827f $X=1.7 $Y=0.17 $X2=0.835 $Y2=1.075
cc_10 N_GND_M1004_b N_B_M1000_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_11 N_GND_M1004_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.96
cc_12 N_GND_M1004_b N_B_c_119_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_13 N_GND_M1004_b N_B_c_120_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_14 N_GND_M1004_b N_A_27_115#_M1001_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_15 N_GND_c_7_p N_A_27_115#_M1001_g 0.0103278f $X=1.05 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_16 N_GND_c_16_p N_A_27_115#_M1001_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_c_3_p N_A_27_115#_M1001_g 0.00468827f $X=1.7 $Y=0.17 $X2=1.335
+ $Y2=1.075
cc_18 N_GND_M1004_b N_A_27_115#_c_158_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.81
cc_19 N_GND_M1004_b N_A_27_115#_c_159_n 0.0244031f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.885
cc_20 N_GND_M1004_b N_A_27_115#_M1006_g 0.0264963f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_21 N_GND_c_21_p N_A_27_115#_M1006_g 0.00713292f $X=1.98 $Y=0.825 $X2=1.765
+ $Y2=1.075
cc_22 N_GND_c_16_p N_A_27_115#_M1006_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=1.075
cc_23 N_GND_c_3_p N_A_27_115#_M1006_g 0.00468827f $X=1.7 $Y=0.17 $X2=1.765
+ $Y2=1.075
cc_24 N_GND_M1004_b N_A_27_115#_c_164_n 0.00567173f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.885
cc_25 N_GND_M1004_b N_A_27_115#_c_165_n 0.0143389f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_26 N_GND_c_2_p N_A_27_115#_c_165_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_27 N_GND_c_3_p N_A_27_115#_c_165_n 0.00476261f $X=1.7 $Y=0.17 $X2=0.26
+ $Y2=0.825
cc_28 N_GND_M1004_b N_A_27_115#_c_168_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.935
cc_29 N_GND_M1004_b N_A_27_115#_c_169_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.935
cc_30 N_GND_M1004_b N_A_27_115#_c_170_n 0.0230268f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_31 N_GND_c_7_p N_A_27_115#_c_170_n 0.00704977f $X=1.05 $Y=0.825 $X2=1.43
+ $Y2=1.935
cc_32 N_GND_M1004_b N_A_27_115#_c_172_n 0.0547984f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_33 N_GND_M1004_b N_A_27_115#_c_173_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.935
cc_34 N_GND_M1004_b N_A_27_115#_c_174_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.545
cc_35 N_GND_M1004_b Y 0.0308484f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_36 N_GND_M1004_b N_Y_c_242_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.48
cc_37 N_GND_c_7_p N_Y_c_242_n 0.00119317f $X=1.05 $Y=0.825 $X2=1.55 $Y2=1.48
cc_38 N_GND_c_21_p N_Y_c_242_n 0.00125659f $X=1.98 $Y=0.825 $X2=1.55 $Y2=1.48
cc_39 N_GND_M1004_b N_Y_c_245_n 0.0111067f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_40 N_GND_M1004_b N_Y_c_246_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_41 N_GND_M1004_b N_Y_c_247_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_42 N_GND_c_7_p N_Y_c_247_n 0.0187614f $X=1.05 $Y=0.825 $X2=1.55 $Y2=0.825
cc_43 N_GND_c_16_p N_Y_c_247_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.825
cc_44 N_GND_c_3_p N_Y_c_247_n 0.00475776f $X=1.7 $Y=0.17 $X2=1.55 $Y2=0.825
cc_45 N_VDD_M1005_b N_A_M1005_g 0.0189471f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_46 N_VDD_c_46_p N_A_M1005_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_47 N_VDD_c_47_p N_A_M1005_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=4.585
cc_48 N_VDD_c_48_p N_A_M1005_g 0.00468827f $X=1.7 $Y=6.49 $X2=0.475 $Y2=4.585
cc_49 N_VDD_M1005_s A 0.00742066f $X=0.135 $Y=3.085 $X2=0.275 $Y2=3.33
cc_50 N_VDD_M1005_b A 0.00970321f $X=-0.045 $Y=2.905 $X2=0.275 $Y2=3.33
cc_51 N_VDD_c_46_p A 0.00434783f $X=0.26 $Y=4.135 $X2=0.275 $Y2=3.33
cc_52 N_VDD_M1005_s N_A_c_84_n 0.0127298f $X=0.135 $Y=3.085 $X2=0.27 $Y2=2.765
cc_53 N_VDD_M1005_b N_A_c_84_n 0.00612103f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.765
cc_54 N_VDD_c_46_p N_A_c_84_n 0.00370742f $X=0.26 $Y=4.135 $X2=0.27 $Y2=2.765
cc_55 N_VDD_M1005_b N_A_c_85_n 0.0111025f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=2.765
cc_56 N_VDD_M1005_b N_B_M1000_g 0.0187476f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_57 N_VDD_c_47_p N_B_M1000_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=4.585
cc_58 N_VDD_c_58_p N_B_M1000_g 0.00354579f $X=1.12 $Y=3.795 $X2=0.905 $Y2=4.585
cc_59 N_VDD_c_48_p N_B_M1000_g 0.00468827f $X=1.7 $Y=6.49 $X2=0.905 $Y2=4.585
cc_60 N_VDD_M1005_b B 0.00856863f $X=-0.045 $Y=2.905 $X2=0.955 $Y2=2.96
cc_61 N_VDD_c_58_p B 0.00240671f $X=1.12 $Y=3.795 $X2=0.955 $Y2=2.96
cc_62 N_VDD_M1005_b N_B_c_119_n 0.00170274f $X=-0.045 $Y=2.905 $X2=0.95
+ $Y2=2.425
cc_63 N_VDD_M1005_b N_A_27_115#_c_175_n 0.017104f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.96
cc_64 N_VDD_c_58_p N_A_27_115#_c_175_n 0.00354579f $X=1.12 $Y=3.795 $X2=1.335
+ $Y2=2.96
cc_65 N_VDD_c_65_p N_A_27_115#_c_175_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.335
+ $Y2=2.96
cc_66 N_VDD_c_48_p N_A_27_115#_c_175_n 0.00468827f $X=1.7 $Y=6.49 $X2=1.335
+ $Y2=2.96
cc_67 N_VDD_M1005_b N_A_27_115#_c_159_n 0.00813142f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.885
cc_68 N_VDD_M1005_b N_A_27_115#_c_180_n 0.0212198f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.96
cc_69 N_VDD_c_58_p N_A_27_115#_c_180_n 3.67508e-19 $X=1.12 $Y=3.795 $X2=1.765
+ $Y2=2.96
cc_70 N_VDD_c_70_p N_A_27_115#_c_180_n 0.00732698f $X=1.98 $Y=3.455 $X2=1.765
+ $Y2=2.96
cc_71 N_VDD_c_65_p N_A_27_115#_c_180_n 0.00610567f $X=1.895 $Y=6.507 $X2=1.765
+ $Y2=2.96
cc_72 N_VDD_c_48_p N_A_27_115#_c_180_n 0.00470215f $X=1.7 $Y=6.49 $X2=1.765
+ $Y2=2.96
cc_73 N_VDD_M1005_b N_A_27_115#_c_164_n 0.00216365f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.885
cc_74 N_VDD_M1005_b N_A_27_115#_c_186_n 0.00155118f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=3.795
cc_75 N_VDD_c_47_p N_A_27_115#_c_186_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69
+ $Y2=3.795
cc_76 N_VDD_c_48_p N_A_27_115#_c_186_n 0.00475776f $X=1.7 $Y=6.49 $X2=0.69
+ $Y2=3.795
cc_77 N_VDD_M1005_b N_A_27_115#_c_174_n 8.22047e-19 $X=-0.045 $Y=2.905 $X2=0.65
+ $Y2=3.545
cc_78 N_VDD_M1005_b N_Y_c_246_n 0.00344954f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.59
cc_79 N_VDD_c_65_p N_Y_c_246_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55 $Y2=2.59
cc_80 N_VDD_c_48_p N_Y_c_246_n 0.00475776f $X=1.7 $Y=6.49 $X2=1.55 $Y2=2.59
cc_81 N_A_M1004_g N_B_M1002_g 0.129148f $X=0.475 $Y=1.075 $X2=0.835 $Y2=1.075
cc_82 N_A_M1004_g N_B_M1000_g 0.0498038f $X=0.475 $Y=1.075 $X2=0.905 $Y2=4.585
cc_83 N_A_M1004_g N_B_c_119_n 7.8234e-19 $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.425
cc_84 N_A_M1004_g N_A_27_115#_c_165_n 0.0158058f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_85 N_A_M1004_g N_A_27_115#_c_168_n 0.0160984f $X=0.475 $Y=1.075 $X2=0.525
+ $Y2=1.935
cc_86 N_A_c_84_n N_A_27_115#_c_168_n 2.65873e-19 $X=0.27 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_87 N_A_c_85_n N_A_27_115#_c_168_n 0.00117122f $X=0.475 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_88 N_A_c_84_n N_A_27_115#_c_169_n 0.0055861f $X=0.27 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_89 N_A_c_85_n N_A_27_115#_c_169_n 0.00133457f $X=0.475 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_90 N_A_M1004_g N_A_27_115#_c_173_n 0.00322084f $X=0.475 $Y=1.075 $X2=0.61
+ $Y2=1.935
cc_91 N_A_M1004_g N_A_27_115#_c_174_n 0.0265302f $X=0.475 $Y=1.075 $X2=0.65
+ $Y2=3.545
cc_92 N_A_M1005_g N_A_27_115#_c_174_n 0.0140172f $X=0.475 $Y=4.585 $X2=0.65
+ $Y2=3.545
cc_93 A N_A_27_115#_c_174_n 0.00758489f $X=0.275 $Y=3.33 $X2=0.65 $Y2=3.545
cc_94 N_A_c_84_n N_A_27_115#_c_174_n 0.0456533f $X=0.27 $Y=2.765 $X2=0.65
+ $Y2=3.545
cc_95 N_A_c_85_n N_A_27_115#_c_174_n 0.00766302f $X=0.475 $Y=2.765 $X2=0.65
+ $Y2=3.545
cc_96 N_A_M1005_g N_A_27_115#_c_202_n 0.00884152f $X=0.475 $Y=4.585 $X2=0.65
+ $Y2=3.715
cc_97 N_B_M1002_g N_A_27_115#_M1001_g 0.0349266f $X=0.835 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_98 N_B_M1000_g N_A_27_115#_c_158_n 0.00773101f $X=0.905 $Y=4.585 $X2=1.37
+ $Y2=2.81
cc_99 N_B_c_119_n N_A_27_115#_c_158_n 0.0033451f $X=0.95 $Y=2.425 $X2=1.37
+ $Y2=2.81
cc_100 N_B_c_120_n N_A_27_115#_c_158_n 0.0206104f $X=0.95 $Y=2.425 $X2=1.37
+ $Y2=2.81
cc_101 N_B_M1000_g N_A_27_115#_c_164_n 0.0400641f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.885
cc_102 B N_A_27_115#_c_164_n 0.00386686f $X=0.955 $Y=2.96 $X2=1.352 $Y2=2.885
cc_103 N_B_c_119_n N_A_27_115#_c_164_n 0.00170598f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.885
cc_104 N_B_M1002_g N_A_27_115#_c_170_n 0.0182215f $X=0.835 $Y=1.075 $X2=1.43
+ $Y2=1.935
cc_105 N_B_c_119_n N_A_27_115#_c_170_n 0.0101796f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_106 N_B_c_120_n N_A_27_115#_c_170_n 0.00258465f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_107 N_B_M1002_g N_A_27_115#_c_172_n 0.0104742f $X=0.835 $Y=1.075 $X2=1.43
+ $Y2=1.935
cc_108 N_B_M1002_g N_A_27_115#_c_174_n 0.00755919f $X=0.835 $Y=1.075 $X2=0.65
+ $Y2=3.545
cc_109 N_B_M1000_g N_A_27_115#_c_174_n 0.0133197f $X=0.905 $Y=4.585 $X2=0.65
+ $Y2=3.545
cc_110 B N_A_27_115#_c_174_n 0.00866797f $X=0.955 $Y=2.96 $X2=0.65 $Y2=3.545
cc_111 N_B_c_119_n N_A_27_115#_c_174_n 0.0541375f $X=0.95 $Y=2.425 $X2=0.65
+ $Y2=3.545
cc_112 B N_A_27_115#_c_202_n 0.00286715f $X=0.955 $Y=2.96 $X2=0.65 $Y2=3.715
cc_113 N_B_M1002_g Y 6.71108e-19 $X=0.835 $Y=1.075 $X2=1.555 $Y2=2.22
cc_114 N_B_c_119_n Y 0.00695761f $X=0.95 $Y=2.425 $X2=1.555 $Y2=2.22
cc_115 N_B_M1002_g N_Y_c_242_n 7.96664e-19 $X=0.835 $Y=1.075 $X2=1.55 $Y2=1.48
cc_116 N_B_c_119_n N_Y_c_245_n 0.00532157f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_117 N_B_c_120_n N_Y_c_245_n 5.70769e-19 $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_118 B N_Y_c_246_n 0.00649253f $X=0.955 $Y=2.96 $X2=1.55 $Y2=2.59
cc_119 N_B_c_119_n N_Y_c_246_n 0.0149875f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_120 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_121 N_A_27_115#_c_158_n Y 0.00892438f $X=1.37 $Y=2.81 $X2=1.555 $Y2=2.22
cc_122 N_A_27_115#_M1006_g Y 0.00251111f $X=1.765 $Y=1.075 $X2=1.555 $Y2=2.22
cc_123 N_A_27_115#_c_170_n Y 0.0148238f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_124 N_A_27_115#_c_172_n Y 0.012094f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_125 N_A_27_115#_M1001_g N_Y_c_242_n 0.0053924f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.48
cc_126 N_A_27_115#_M1006_g N_Y_c_242_n 0.00908199f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=1.48
cc_127 N_A_27_115#_c_170_n N_Y_c_242_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.48
cc_128 N_A_27_115#_c_158_n N_Y_c_245_n 0.00740115f $X=1.37 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_129 N_A_27_115#_c_159_n N_Y_c_245_n 0.00229755f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.59
cc_130 N_A_27_115#_c_170_n N_Y_c_245_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_131 N_A_27_115#_c_172_n N_Y_c_245_n 0.00174847f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_132 N_A_27_115#_c_175_n N_Y_c_246_n 0.00278785f $X=1.335 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_133 N_A_27_115#_c_158_n N_Y_c_246_n 0.00744772f $X=1.37 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_134 N_A_27_115#_c_159_n N_Y_c_246_n 0.0159823f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.59
cc_135 N_A_27_115#_c_180_n N_Y_c_246_n 0.00392729f $X=1.765 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_136 N_A_27_115#_c_170_n N_Y_c_246_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_137 N_A_27_115#_c_172_n N_Y_c_246_n 0.0013767f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_138 N_A_27_115#_M1001_g N_Y_c_247_n 0.00233629f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_139 N_A_27_115#_M1006_g N_Y_c_247_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_140 N_A_27_115#_c_170_n N_Y_c_247_n 0.00500271f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_141 N_A_27_115#_c_172_n N_Y_c_247_n 0.00171364f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
