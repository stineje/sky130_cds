* File: sky130_osu_sc_18T_hs__pcgateCKa_new.spice
* Created: Thu Mar 10 17:12:01 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_hs__pcgateCKa_new.pex.spice"
.subckt sky130_osu_sc_18T_hs__pcgateCKa_new  GND VDD SE E CK CKA Q ECK
* 
* ECK	ECK
* Q	Q
* CKA	CKA
* CK	CK
* E	E
* SE	SE
* VDD	VDD
* GND	GND
MM1010 N_A_N233_617#_M1010_d N_SE_M1010_g N_GND_M1010_s N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_GND_M1020_d N_E_M1020_g N_A_N233_617#_M1010_d N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1025 N_GND_M1025_d N_A_86_337#_M1025_g N_A_43_115#_M1025_s N_GND_M1010_b
+ NLOWVT L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1023 A_212_115# N_A_N233_617#_M1023_g N_GND_M1025_d N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1021 N_A_86_337#_M1021_d N_A_254_89#_M1021_g A_212_115# N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1
+ R=6.66667 SA=75001 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1011 A_404_115# N_CK_M1011_g N_A_86_337#_M1021_d N_GND_M1010_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.6 SB=75001 A=0.15 P=2.3 MULT=1
MM1002 N_GND_M1002_d N_A_43_115#_M1002_g A_404_115# N_GND_M1010_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_254_89#_M1003_d N_CK_M1003_g N_GND_M1002_d N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1018 N_GND_M1018_d N_A_43_115#_M1018_g N_A_687_115#_M1018_s N_GND_M1010_b
+ NLOWVT L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_Q_M1005_d N_A_687_115#_M1005_g N_GND_M1018_d N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1015 A_1046_115# N_A_687_115#_M1015_g N_A_963_115#_M1015_s N_GND_M1010_b
+ NLOWVT L=0.15 W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1012 N_GND_M1012_d N_CKA_M1012_g A_1046_115# N_GND_M1010_b NLOWVT L=0.15 W=1
+ AD=0.175 AS=0.105 PD=1.35 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75000.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_ECK_M1009_d N_A_963_115#_M1009_g N_GND_M1012_d N_GND_M1010_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.175 PD=2.53 PS=1.35 NRD=0 NRS=8.388 M=1 R=6.66667
+ SA=75001 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 A_N150_617# N_SE_M1007_g N_A_N233_617#_M1007_s N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20
+ SA=75000.2 SB=75000.5 A=0.45 P=6.3 MULT=1
MM1013 N_VDD_M1013_d N_E_M1013_g A_N150_617# N_VDD_M1007_b PSHORT L=0.15 W=3
+ AD=0.795 AS=0.315 PD=6.53 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75000.5
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1024 N_VDD_M1024_d N_A_86_337#_M1024_g N_A_43_115#_M1024_s N_VDD_M1007_b
+ PSHORT L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20
+ SA=75000.2 SB=75002.4 A=0.45 P=6.3 MULT=1
MM1022 A_212_617# N_A_N233_617#_M1022_g N_VDD_M1024_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20
+ SA=75000.6 SB=75001.9 A=0.45 P=6.3 MULT=1
MM1019 N_A_86_337#_M1019_d N_CK_M1019_g A_212_617# N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20 SA=75001
+ SB=75001.6 A=0.45 P=6.3 MULT=1
MM1008 A_404_617# N_A_254_89#_M1008_g N_A_86_337#_M1019_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75001.6 SB=75001 A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_A_43_115#_M1000_g A_404_617# N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.9
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1001 N_A_254_89#_M1001_d N_CK_M1001_g N_VDD_M1000_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.4
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1016 N_VDD_M1016_d N_A_43_115#_M1016_g N_A_687_115#_M1016_s N_VDD_M1007_b
+ PSHORT L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20
+ SA=75000.2 SB=75000.6 A=0.45 P=6.3 MULT=1
MM1004 N_Q_M1004_d N_A_687_115#_M1004_g N_VDD_M1016_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1014 N_A_963_115#_M1014_d N_A_687_115#_M1014_g N_VDD_M1014_s N_VDD_M1007_b
+ PSHORT L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20
+ SA=75000.2 SB=75001 A=0.45 P=6.3 MULT=1
MM1017 N_VDD_M1017_d N_CKA_M1017_g N_A_963_115#_M1014_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1006 N_ECK_M1006_d N_A_963_115#_M1006_g N_VDD_M1017_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX26_noxref N_GND_M1010_b N_VDD_M1007_b NWDIODE A=30.1404 P=23.47
pX27_noxref noxref_21 N_SE_X27_noxref_CONDUCTOR SE PROBETYPE=1
pX28_noxref noxref_22 E E PROBETYPE=1
pX29_noxref noxref_23 CK CK PROBETYPE=1
pX30_noxref noxref_24 Q Q PROBETYPE=1
pX31_noxref noxref_25 CKA CKA PROBETYPE=1
pX32_noxref noxref_26 ECK ECK PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__pcgateCKa_new.pxi.spice"
*
.ends
*
*
