* File: sky130_osu_sc_18T_ls__dff_1.pxi.spice
* Created: Fri Nov 12 14:15:31 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%GND N_GND_M1004_d N_GND_M1013_d N_GND_M1022_d
+ N_GND_M1006_s N_GND_M1008_d N_GND_M1004_b N_GND_c_2_p N_GND_c_3_p N_GND_c_14_p
+ N_GND_c_59_p N_GND_c_35_p N_GND_c_39_p N_GND_c_40_p N_GND_c_41_p N_GND_c_118_p
+ N_GND_c_119_p GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_LS__DFF_1%GND
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%VDD N_VDD_M1020_d N_VDD_M1016_d N_VDD_M1001_d
+ N_VDD_M1023_s N_VDD_M1011_d N_VDD_M1020_b N_VDD_c_173_p N_VDD_c_174_p
+ N_VDD_c_183_p N_VDD_c_210_p N_VDD_c_194_p N_VDD_c_198_p N_VDD_c_199_p
+ N_VDD_c_200_p N_VDD_c_241_p N_VDD_c_242_p N_VDD_c_257_p VDD N_VDD_c_175_p
+ PM_SKY130_OSU_SC_18T_LS__DFF_1%VDD
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%A_75_344# N_A_75_344#_M1021_d
+ N_A_75_344#_M1009_d N_A_75_344#_M1004_g N_A_75_344#_M1020_g
+ N_A_75_344#_c_275_n N_A_75_344#_c_276_n N_A_75_344#_c_277_n
+ N_A_75_344#_c_293_n N_A_75_344#_c_278_n N_A_75_344#_c_280_n
+ N_A_75_344#_c_294_n N_A_75_344#_c_296_n N_A_75_344#_c_282_n
+ N_A_75_344#_c_283_n N_A_75_344#_c_298_n N_A_75_344#_c_286_n
+ N_A_75_344#_c_287_n N_A_75_344#_c_319_p
+ PM_SKY130_OSU_SC_18T_LS__DFF_1%A_75_344#
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%D N_D_M1003_g N_D_M1007_g N_D_c_362_n
+ N_D_c_363_n D PM_SKY130_OSU_SC_18T_LS__DFF_1%D
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%CK N_CK_M1009_g N_CK_M1018_g N_CK_M1010_g
+ N_CK_M1012_g N_CK_M1024_g N_CK_c_400_n N_CK_M1017_g N_CK_c_401_n N_CK_c_402_n
+ N_CK_c_403_n N_CK_c_404_n N_CK_c_407_n N_CK_c_408_n N_CK_c_411_n N_CK_c_412_n
+ N_CK_c_417_n N_CK_c_418_n N_CK_c_419_n N_CK_c_420_n N_CK_c_421_n N_CK_c_422_n
+ N_CK_c_423_n N_CK_c_424_n N_CK_c_425_n N_CK_c_426_n N_CK_c_427_n N_CK_c_428_n
+ N_CK_c_429_n CK PM_SKY130_OSU_SC_18T_LS__DFF_1%CK
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%A_32_115# N_A_32_115#_M1004_s
+ N_A_32_115#_M1020_s N_A_32_115#_M1013_g N_A_32_115#_M1016_g
+ N_A_32_115#_c_617_n N_A_32_115#_c_619_n N_A_32_115#_c_620_n
+ N_A_32_115#_c_621_n N_A_32_115#_M1015_g N_A_32_115#_M1005_g
+ N_A_32_115#_c_626_n N_A_32_115#_c_627_n N_A_32_115#_c_647_n
+ N_A_32_115#_c_630_n N_A_32_115#_c_631_n N_A_32_115#_c_652_n
+ N_A_32_115#_c_632_n N_A_32_115#_c_634_n N_A_32_115#_c_636_n
+ N_A_32_115#_c_698_n PM_SKY130_OSU_SC_18T_LS__DFF_1%A_32_115#
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%A_243_89# N_A_243_89#_M1024_d
+ N_A_243_89#_M1017_d N_A_243_89#_c_728_n N_A_243_89#_M1021_g
+ N_A_243_89#_c_731_n N_A_243_89#_c_732_n N_A_243_89#_c_733_n
+ N_A_243_89#_M1014_g N_A_243_89#_c_735_n N_A_243_89#_M1019_g
+ N_A_243_89#_c_737_n N_A_243_89#_c_738_n N_A_243_89#_M1000_g
+ N_A_243_89#_c_739_n N_A_243_89#_c_740_n N_A_243_89#_c_741_n
+ N_A_243_89#_c_742_n N_A_243_89#_c_743_n N_A_243_89#_c_746_n
+ N_A_243_89#_c_748_n N_A_243_89#_c_752_n N_A_243_89#_c_762_n
+ N_A_243_89#_c_753_n N_A_243_89#_c_754_n N_A_243_89#_c_755_n
+ N_A_243_89#_c_767_n PM_SKY130_OSU_SC_18T_LS__DFF_1%A_243_89#
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%A_785_89# N_A_785_89#_M1006_d
+ N_A_785_89#_M1023_d N_A_785_89#_M1022_g N_A_785_89#_M1001_g
+ N_A_785_89#_M1008_g N_A_785_89#_M1011_g N_A_785_89#_c_907_n
+ N_A_785_89#_c_908_n N_A_785_89#_c_909_n N_A_785_89#_c_910_n
+ N_A_785_89#_c_914_n N_A_785_89#_c_915_n N_A_785_89#_c_916_n
+ N_A_785_89#_c_917_n N_A_785_89#_c_918_n N_A_785_89#_c_921_n
+ N_A_785_89#_c_922_n N_A_785_89#_c_923_n N_A_785_89#_c_924_n
+ N_A_785_89#_c_925_n N_A_785_89#_c_926_n
+ PM_SKY130_OSU_SC_18T_LS__DFF_1%A_785_89#
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%A_623_115# N_A_623_115#_M1010_d
+ N_A_623_115#_M1019_d N_A_623_115#_c_1033_n N_A_623_115#_M1006_g
+ N_A_623_115#_M1023_g N_A_623_115#_c_1038_n N_A_623_115#_c_1040_n
+ N_A_623_115#_c_1067_n N_A_623_115#_c_1096_n N_A_623_115#_c_1070_n
+ N_A_623_115#_c_1098_n N_A_623_115#_c_1041_n N_A_623_115#_c_1056_n
+ N_A_623_115#_c_1044_n N_A_623_115#_c_1046_n N_A_623_115#_c_1048_n
+ N_A_623_115#_c_1049_n PM_SKY130_OSU_SC_18T_LS__DFF_1%A_623_115#
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%QN N_QN_M1008_s N_QN_M1011_s N_QN_M1025_g
+ N_QN_M1002_g N_QN_c_1152_n N_QN_c_1153_n N_QN_c_1156_n N_QN_c_1157_n
+ N_QN_c_1159_n N_QN_c_1160_n N_QN_c_1161_n N_QN_c_1162_n QN
+ PM_SKY130_OSU_SC_18T_LS__DFF_1%QN
x_PM_SKY130_OSU_SC_18T_LS__DFF_1%Q N_Q_M1025_d N_Q_M1002_d N_Q_c_1227_n
+ N_Q_c_1231_n N_Q_c_1229_n N_Q_c_1230_n N_Q_c_1235_n Q
+ PM_SKY130_OSU_SC_18T_LS__DFF_1%Q
cc_1 N_GND_M1004_b N_A_75_344#_M1004_g 0.0223692f $X=-0.045 $Y=0 $X2=0.5
+ $Y2=1.075
cc_2 N_GND_c_2_p N_A_75_344#_M1004_g 0.00606474f $X=0.63 $Y=0.152 $X2=0.5
+ $Y2=1.075
cc_3 N_GND_c_3_p N_A_75_344#_M1004_g 0.00354579f $X=0.715 $Y=0.825 $X2=0.5
+ $Y2=1.075
cc_4 N_GND_c_4_p N_A_75_344#_M1004_g 0.00468827f $X=6.46 $Y=0.19 $X2=0.5
+ $Y2=1.075
cc_5 N_GND_M1004_b N_A_75_344#_c_275_n 0.0143449f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=1.87
cc_6 N_GND_M1004_b N_A_75_344#_c_276_n 0.0223136f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.765
cc_7 N_GND_M1004_b N_A_75_344#_c_277_n 0.0431517f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.6
cc_8 N_GND_M1004_b N_A_75_344#_c_278_n 0.0183015f $X=-0.045 $Y=0 $X2=1.405
+ $Y2=1.765
cc_9 N_GND_c_3_p N_A_75_344#_c_278_n 0.00456782f $X=0.715 $Y=0.825 $X2=1.405
+ $Y2=1.765
cc_10 N_GND_M1004_b N_A_75_344#_c_280_n 0.00315644f $X=-0.045 $Y=0 $X2=0.71
+ $Y2=1.765
cc_11 N_GND_c_3_p N_A_75_344#_c_280_n 0.00460441f $X=0.715 $Y=0.825 $X2=0.71
+ $Y2=1.765
cc_12 N_GND_M1004_b N_A_75_344#_c_282_n 0.00198494f $X=-0.045 $Y=0 $X2=1.49
+ $Y2=1.68
cc_13 N_GND_M1004_b N_A_75_344#_c_283_n 0.00313975f $X=-0.045 $Y=0 $X2=1.59
+ $Y2=0.825
cc_14 N_GND_c_14_p N_A_75_344#_c_283_n 0.0149076f $X=2.38 $Y=0.152 $X2=1.59
+ $Y2=0.825
cc_15 N_GND_c_4_p N_A_75_344#_c_283_n 0.00958198f $X=6.46 $Y=0.19 $X2=1.59
+ $Y2=0.825
cc_16 N_GND_M1004_b N_A_75_344#_c_286_n 0.00325766f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.765
cc_17 N_GND_M1004_b N_A_75_344#_c_287_n 0.0127034f $X=-0.045 $Y=0 $X2=0.567
+ $Y2=2.6
cc_18 N_GND_M1004_b N_D_M1003_g 0.0334344f $X=-0.045 $Y=0 $X2=0.93 $Y2=1.075
cc_19 N_GND_c_3_p N_D_M1003_g 0.00354579f $X=0.715 $Y=0.825 $X2=0.93 $Y2=1.075
cc_20 N_GND_c_14_p N_D_M1003_g 0.00606474f $X=2.38 $Y=0.152 $X2=0.93 $Y2=1.075
cc_21 N_GND_c_4_p N_D_M1003_g 0.00468827f $X=6.46 $Y=0.19 $X2=0.93 $Y2=1.075
cc_22 N_GND_M1004_b N_D_M1007_g 0.0299924f $X=-0.045 $Y=0 $X2=0.93 $Y2=4.585
cc_23 N_GND_M1004_b N_D_c_362_n 0.0272793f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.22
cc_24 N_GND_M1004_b N_D_c_363_n 0.00311208f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.22
cc_25 N_GND_M1004_b D 0.00874398f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.22
cc_26 N_GND_M1004_b N_CK_c_400_n 0.0311248f $X=-0.045 $Y=0 $X2=4.43 $Y2=2.93
cc_27 N_GND_M1004_b N_CK_c_401_n 0.0438842f $X=-0.045 $Y=0 $X2=4.485 $Y2=2.6
cc_28 N_GND_M1004_b N_CK_c_402_n 0.0244054f $X=-0.045 $Y=0 $X2=1.35 $Y2=2.765
cc_29 N_GND_M1004_b N_CK_c_403_n 0.0254608f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.85
cc_30 N_GND_M1004_b N_CK_c_404_n 0.0173906f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.685
cc_31 N_GND_c_14_p N_CK_c_404_n 0.00606474f $X=2.38 $Y=0.152 $X2=1.83 $Y2=1.685
cc_32 N_GND_c_4_p N_CK_c_404_n 0.00468827f $X=6.46 $Y=0.19 $X2=1.83 $Y2=1.685
cc_33 N_GND_M1004_b N_CK_c_407_n 0.0252285f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.85
cc_34 N_GND_M1004_b N_CK_c_408_n 0.0175305f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.685
cc_35 N_GND_c_35_p N_CK_c_408_n 0.00606474f $X=4.13 $Y=0.152 $X2=3.1 $Y2=1.685
cc_36 N_GND_c_4_p N_CK_c_408_n 0.00468827f $X=6.46 $Y=0.19 $X2=3.1 $Y2=1.685
cc_37 N_GND_M1004_b N_CK_c_411_n 0.0233827f $X=-0.045 $Y=0 $X2=3.58 $Y2=2.765
cc_38 N_GND_M1004_b N_CK_c_412_n 0.0183851f $X=-0.045 $Y=0 $X2=4.457 $Y2=1.685
cc_39 N_GND_c_39_p N_CK_c_412_n 0.00354579f $X=4.215 $Y=0.825 $X2=4.457
+ $Y2=1.685
cc_40 N_GND_c_40_p N_CK_c_412_n 0.00606474f $X=5.08 $Y=0.152 $X2=4.457 $Y2=1.685
cc_41 N_GND_c_41_p N_CK_c_412_n 0.00463923f $X=5.165 $Y=0.825 $X2=4.457
+ $Y2=1.685
cc_42 N_GND_c_4_p N_CK_c_412_n 0.00468827f $X=6.46 $Y=0.19 $X2=4.457 $Y2=1.685
cc_43 N_GND_M1004_b N_CK_c_417_n 0.01373f $X=-0.045 $Y=0 $X2=4.457 $Y2=1.835
cc_44 N_GND_M1004_b N_CK_c_418_n 0.00600607f $X=-0.045 $Y=0 $X2=1.745 $Y2=2.59
cc_45 N_GND_M1004_b N_CK_c_419_n 0.0108248f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.85
cc_46 N_GND_M1004_b N_CK_c_420_n 0.00852144f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.85
cc_47 N_GND_M1004_b N_CK_c_421_n 0.00543853f $X=-0.045 $Y=0 $X2=3.495 $Y2=2.59
cc_48 N_GND_M1004_b N_CK_c_422_n 5.00459e-19 $X=-0.045 $Y=0 $X2=3.185 $Y2=2.59
cc_49 N_GND_M1004_b N_CK_c_423_n 7.61111e-19 $X=-0.045 $Y=0 $X2=4.575 $Y2=2.59
cc_50 N_GND_M1004_b N_CK_c_424_n 0.00235115f $X=-0.045 $Y=0 $X2=1.35 $Y2=2.59
cc_51 N_GND_M1004_b N_CK_c_425_n 0.00265612f $X=-0.045 $Y=0 $X2=3.58 $Y2=2.59
cc_52 N_GND_M1004_b N_CK_c_426_n 0.0341675f $X=-0.045 $Y=0 $X2=3.435 $Y2=2.59
cc_53 N_GND_M1004_b N_CK_c_427_n 0.00614962f $X=-0.045 $Y=0 $X2=1.495 $Y2=2.59
cc_54 N_GND_M1004_b N_CK_c_428_n 0.0181831f $X=-0.045 $Y=0 $X2=4.43 $Y2=2.59
cc_55 N_GND_M1004_b N_CK_c_429_n 0.0041728f $X=-0.045 $Y=0 $X2=3.725 $Y2=2.59
cc_56 N_GND_M1004_b CK 0.00239232f $X=-0.045 $Y=0 $X2=4.575 $Y2=2.59
cc_57 N_GND_M1004_b N_A_32_115#_M1013_g 0.0171814f $X=-0.045 $Y=0 $X2=2.25
+ $Y2=1.075
cc_58 N_GND_c_14_p N_A_32_115#_M1013_g 0.00606474f $X=2.38 $Y=0.152 $X2=2.25
+ $Y2=1.075
cc_59 N_GND_c_59_p N_A_32_115#_M1013_g 0.00354579f $X=2.465 $Y=0.825 $X2=2.25
+ $Y2=1.075
cc_60 N_GND_c_4_p N_A_32_115#_M1013_g 0.00468827f $X=6.46 $Y=0.19 $X2=2.25
+ $Y2=1.075
cc_61 N_GND_M1004_b N_A_32_115#_c_617_n 0.0240953f $X=-0.045 $Y=0 $X2=2.605
+ $Y2=1.85
cc_62 N_GND_c_59_p N_A_32_115#_c_617_n 8.07204e-19 $X=2.465 $Y=0.825 $X2=2.605
+ $Y2=1.85
cc_63 N_GND_M1004_b N_A_32_115#_c_619_n 0.0105855f $X=-0.045 $Y=0 $X2=2.325
+ $Y2=1.85
cc_64 N_GND_M1004_b N_A_32_115#_c_620_n 0.0232417f $X=-0.045 $Y=0 $X2=2.605
+ $Y2=2.765
cc_65 N_GND_M1004_b N_A_32_115#_c_621_n 0.0105265f $X=-0.045 $Y=0 $X2=2.325
+ $Y2=2.765
cc_66 N_GND_M1004_b N_A_32_115#_M1015_g 0.0163216f $X=-0.045 $Y=0 $X2=2.68
+ $Y2=1.075
cc_67 N_GND_c_59_p N_A_32_115#_M1015_g 0.00354579f $X=2.465 $Y=0.825 $X2=2.68
+ $Y2=1.075
cc_68 N_GND_c_35_p N_A_32_115#_M1015_g 0.00606474f $X=4.13 $Y=0.152 $X2=2.68
+ $Y2=1.075
cc_69 N_GND_c_4_p N_A_32_115#_M1015_g 0.00468827f $X=6.46 $Y=0.19 $X2=2.68
+ $Y2=1.075
cc_70 N_GND_M1004_b N_A_32_115#_c_626_n 0.0456538f $X=-0.045 $Y=0 $X2=0.17
+ $Y2=3.14
cc_71 N_GND_M1004_b N_A_32_115#_c_627_n 0.00613464f $X=-0.045 $Y=0 $X2=0.285
+ $Y2=0.825
cc_72 N_GND_c_2_p N_A_32_115#_c_627_n 0.00736239f $X=0.63 $Y=0.152 $X2=0.285
+ $Y2=0.825
cc_73 N_GND_c_4_p N_A_32_115#_c_627_n 0.00476261f $X=6.46 $Y=0.19 $X2=0.285
+ $Y2=0.825
cc_74 N_GND_M1004_b N_A_32_115#_c_630_n 0.00871176f $X=-0.045 $Y=0 $X2=2.42
+ $Y2=2.765
cc_75 N_GND_M1004_b N_A_32_115#_c_631_n 0.0203007f $X=-0.045 $Y=0 $X2=0.285
+ $Y2=1.85
cc_76 N_GND_M1004_b N_A_32_115#_c_632_n 0.00433237f $X=-0.045 $Y=0 $X2=2.42
+ $Y2=1.85
cc_77 N_GND_c_59_p N_A_32_115#_c_632_n 0.00449229f $X=2.465 $Y=0.825 $X2=2.42
+ $Y2=1.85
cc_78 N_GND_M1004_b N_A_32_115#_c_634_n 0.0225319f $X=-0.045 $Y=0 $X2=2.185
+ $Y2=1.85
cc_79 N_GND_c_3_p N_A_32_115#_c_634_n 0.00118122f $X=0.715 $Y=0.825 $X2=2.185
+ $Y2=1.85
cc_80 N_GND_M1004_b N_A_32_115#_c_636_n 0.00468924f $X=-0.045 $Y=0 $X2=0.43
+ $Y2=1.85
cc_81 N_GND_M1004_b N_A_243_89#_c_728_n 0.0173059f $X=-0.045 $Y=0 $X2=1.29
+ $Y2=1.685
cc_82 N_GND_c_14_p N_A_243_89#_c_728_n 0.00606474f $X=2.38 $Y=0.152 $X2=1.29
+ $Y2=1.685
cc_83 N_GND_c_4_p N_A_243_89#_c_728_n 0.00468827f $X=6.46 $Y=0.19 $X2=1.29
+ $Y2=1.685
cc_84 N_GND_M1004_b N_A_243_89#_c_731_n 0.0202867f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.225
cc_85 N_GND_M1004_b N_A_243_89#_c_732_n 0.0187566f $X=-0.045 $Y=0 $X2=1.815
+ $Y2=2.3
cc_86 N_GND_M1004_b N_A_243_89#_c_733_n 0.00755029f $X=-0.045 $Y=0 $X2=1.485
+ $Y2=2.3
cc_87 N_GND_M1004_b N_A_243_89#_M1014_g 0.032457f $X=-0.045 $Y=0 $X2=1.89
+ $Y2=4.585
cc_88 N_GND_M1004_b N_A_243_89#_c_735_n 0.0559794f $X=-0.045 $Y=0 $X2=2.965
+ $Y2=2.3
cc_89 N_GND_M1004_b N_A_243_89#_M1019_g 0.0319667f $X=-0.045 $Y=0 $X2=3.04
+ $Y2=4.585
cc_90 N_GND_M1004_b N_A_243_89#_c_737_n 0.0270462f $X=-0.045 $Y=0 $X2=3.445
+ $Y2=2.3
cc_91 N_GND_M1004_b N_A_243_89#_c_738_n 0.0125754f $X=-0.045 $Y=0 $X2=3.52
+ $Y2=2.225
cc_92 N_GND_M1004_b N_A_243_89#_c_739_n 0.0141451f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.76
cc_93 N_GND_M1004_b N_A_243_89#_c_740_n 0.00426512f $X=-0.045 $Y=0 $X2=1.89
+ $Y2=2.3
cc_94 N_GND_M1004_b N_A_243_89#_c_741_n 0.00426512f $X=-0.045 $Y=0 $X2=3.04
+ $Y2=2.3
cc_95 N_GND_M1004_b N_A_243_89#_c_742_n 0.0265388f $X=-0.045 $Y=0 $X2=3.58
+ $Y2=1.85
cc_96 N_GND_M1004_b N_A_243_89#_c_743_n 0.01755f $X=-0.045 $Y=0 $X2=3.58
+ $Y2=1.685
cc_97 N_GND_c_35_p N_A_243_89#_c_743_n 0.00606474f $X=4.13 $Y=0.152 $X2=3.58
+ $Y2=1.685
cc_98 N_GND_c_4_p N_A_243_89#_c_743_n 0.00468827f $X=6.46 $Y=0.19 $X2=3.58
+ $Y2=1.685
cc_99 N_GND_M1004_b N_A_243_89#_c_746_n 0.0116005f $X=-0.045 $Y=0 $X2=4.56
+ $Y2=1.85
cc_100 N_GND_c_39_p N_A_243_89#_c_746_n 0.00572623f $X=4.215 $Y=0.825 $X2=4.56
+ $Y2=1.85
cc_101 N_GND_M1004_b N_A_243_89#_c_748_n 0.00549177f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=0.825
cc_102 N_GND_c_40_p N_A_243_89#_c_748_n 0.00749582f $X=5.08 $Y=0.152 $X2=4.645
+ $Y2=0.825
cc_103 N_GND_c_41_p N_A_243_89#_c_748_n 0.0358835f $X=5.165 $Y=0.825 $X2=4.645
+ $Y2=0.825
cc_104 N_GND_c_4_p N_A_243_89#_c_748_n 0.00476261f $X=6.46 $Y=0.19 $X2=4.645
+ $Y2=0.825
cc_105 N_GND_M1004_b N_A_243_89#_c_752_n 0.00324634f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=2.105
cc_106 N_GND_M1004_b N_A_243_89#_c_753_n 0.0141454f $X=-0.045 $Y=0 $X2=4.915
+ $Y2=3.1
cc_107 N_GND_M1004_b N_A_243_89#_c_754_n 8.79856e-19 $X=-0.045 $Y=0 $X2=4.645
+ $Y2=1.85
cc_108 N_GND_M1004_b N_A_243_89#_c_755_n 0.0100851f $X=-0.045 $Y=0 $X2=4.915
+ $Y2=2.19
cc_109 N_GND_M1004_b N_A_785_89#_M1022_g 0.0319752f $X=-0.045 $Y=0 $X2=4
+ $Y2=1.075
cc_110 N_GND_c_35_p N_A_785_89#_M1022_g 0.00606474f $X=4.13 $Y=0.152 $X2=4
+ $Y2=1.075
cc_111 N_GND_c_39_p N_A_785_89#_M1022_g 0.00354579f $X=4.215 $Y=0.825 $X2=4
+ $Y2=1.075
cc_112 N_GND_c_4_p N_A_785_89#_M1022_g 0.00468827f $X=6.46 $Y=0.19 $X2=4
+ $Y2=1.075
cc_113 N_GND_M1004_b N_A_785_89#_M1001_g 0.0330331f $X=-0.045 $Y=0 $X2=4
+ $Y2=4.585
cc_114 N_GND_M1004_b N_A_785_89#_c_907_n 0.0263478f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=2.19
cc_115 N_GND_M1004_b N_A_785_89#_c_908_n 0.0291536f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=2.19
cc_116 N_GND_M1004_b N_A_785_89#_c_909_n 0.0138254f $X=-0.045 $Y=0 $X2=6.217
+ $Y2=2.025
cc_117 N_GND_M1004_b N_A_785_89#_c_910_n 0.0186503f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=1.65
cc_118 N_GND_c_118_p N_A_785_89#_c_910_n 0.00606474f $X=6.46 $Y=0.152 $X2=6.305
+ $Y2=1.65
cc_119 N_GND_c_119_p N_A_785_89#_c_910_n 0.00354579f $X=6.545 $Y=0.825 $X2=6.305
+ $Y2=1.65
cc_120 N_GND_c_4_p N_A_785_89#_c_910_n 0.00468827f $X=6.46 $Y=0.19 $X2=6.305
+ $Y2=1.65
cc_121 N_GND_M1004_b N_A_785_89#_c_914_n 0.0135453f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=1.8
cc_122 N_GND_M1004_b N_A_785_89#_c_915_n 0.0305585f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=2.855
cc_123 N_GND_M1004_b N_A_785_89#_c_916_n 0.00495925f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=3.005
cc_124 N_GND_M1004_b N_A_785_89#_c_917_n 0.0039674f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=2.19
cc_125 N_GND_M1004_b N_A_785_89#_c_918_n 0.0136393f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=0.825
cc_126 N_GND_c_118_p N_A_785_89#_c_918_n 0.0074445f $X=6.46 $Y=0.152 $X2=5.595
+ $Y2=0.825
cc_127 N_GND_c_4_p N_A_785_89#_c_918_n 0.00476261f $X=6.46 $Y=0.19 $X2=5.595
+ $Y2=0.825
cc_128 N_GND_M1004_b N_A_785_89#_c_921_n 0.0162343f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=3.455
cc_129 N_GND_M1004_b N_A_785_89#_c_922_n 0.0123965f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=2.19
cc_130 N_GND_M1004_b N_A_785_89#_c_923_n 0.00241536f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=2.19
cc_131 N_GND_M1004_b N_A_785_89#_c_924_n 0.0515942f $X=-0.045 $Y=0 $X2=6.07
+ $Y2=2.19
cc_132 N_GND_M1004_b N_A_785_89#_c_925_n 0.00189525f $X=-0.045 $Y=0 $X2=4.205
+ $Y2=2.19
cc_133 N_GND_M1004_b N_A_785_89#_c_926_n 0.00128332f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=2.19
cc_134 N_GND_M1004_b N_A_623_115#_c_1033_n 0.0221119f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=1.685
cc_135 N_GND_c_41_p N_A_623_115#_c_1033_n 0.00713292f $X=5.165 $Y=0.825 $X2=5.38
+ $Y2=1.685
cc_136 N_GND_c_118_p N_A_623_115#_c_1033_n 0.00606474f $X=6.46 $Y=0.152 $X2=5.38
+ $Y2=1.685
cc_137 N_GND_c_4_p N_A_623_115#_c_1033_n 0.00468827f $X=6.46 $Y=0.19 $X2=5.38
+ $Y2=1.685
cc_138 N_GND_M1004_b N_A_623_115#_M1023_g 0.0594514f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=4.585
cc_139 N_GND_M1004_b N_A_623_115#_c_1038_n 0.0482669f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=1.85
cc_140 N_GND_c_41_p N_A_623_115#_c_1038_n 0.00386381f $X=5.165 $Y=0.825 $X2=5.38
+ $Y2=1.85
cc_141 N_GND_M1004_b N_A_623_115#_c_1040_n 0.0112983f $X=-0.045 $Y=0 $X2=2.76
+ $Y2=1.85
cc_142 N_GND_M1004_b N_A_623_115#_c_1041_n 0.00313975f $X=-0.045 $Y=0 $X2=3.34
+ $Y2=0.825
cc_143 N_GND_c_35_p N_A_623_115#_c_1041_n 0.0151257f $X=4.13 $Y=0.152 $X2=3.34
+ $Y2=0.825
cc_144 N_GND_c_4_p N_A_623_115#_c_1041_n 0.00958198f $X=6.46 $Y=0.19 $X2=3.34
+ $Y2=0.825
cc_145 N_GND_M1004_b N_A_623_115#_c_1044_n 0.00161958f $X=-0.045 $Y=0 $X2=5.175
+ $Y2=1.85
cc_146 N_GND_c_41_p N_A_623_115#_c_1044_n 0.00509685f $X=5.165 $Y=0.825
+ $X2=5.175 $Y2=1.85
cc_147 N_GND_M1004_b N_A_623_115#_c_1046_n 0.0393047f $X=-0.045 $Y=0 $X2=5.03
+ $Y2=1.85
cc_148 N_GND_c_39_p N_A_623_115#_c_1046_n 0.00414959f $X=4.215 $Y=0.825 $X2=5.03
+ $Y2=1.85
cc_149 N_GND_M1004_b N_A_623_115#_c_1048_n 0.00143382f $X=-0.045 $Y=0 $X2=2.905
+ $Y2=1.85
cc_150 N_GND_M1004_b N_A_623_115#_c_1049_n 9.64388e-19 $X=-0.045 $Y=0 $X2=5.175
+ $Y2=1.85
cc_151 N_GND_c_41_p N_A_623_115#_c_1049_n 0.00387325f $X=5.165 $Y=0.825
+ $X2=5.175 $Y2=1.85
cc_152 N_GND_M1004_b N_QN_M1025_g 0.0561449f $X=-0.045 $Y=0 $X2=6.76 $Y2=1.075
cc_153 N_GND_c_119_p N_QN_M1025_g 0.00354579f $X=6.545 $Y=0.825 $X2=6.76
+ $Y2=1.075
cc_154 N_GND_c_4_p N_QN_M1025_g 0.00468827f $X=6.46 $Y=0.19 $X2=6.76 $Y2=1.075
cc_155 N_GND_M1004_b N_QN_M1002_g 0.0186095f $X=-0.045 $Y=0 $X2=6.76 $Y2=4.585
cc_156 N_GND_M1004_b N_QN_c_1152_n 0.0291912f $X=-0.045 $Y=0 $X2=6.7 $Y2=2.395
cc_157 N_GND_M1004_b N_QN_c_1153_n 0.00514553f $X=-0.045 $Y=0 $X2=6.115
+ $Y2=0.825
cc_158 N_GND_c_118_p N_QN_c_1153_n 0.00757793f $X=6.46 $Y=0.152 $X2=6.115
+ $Y2=0.825
cc_159 N_GND_c_4_p N_QN_c_1153_n 0.00476261f $X=6.46 $Y=0.19 $X2=6.115 $Y2=0.825
cc_160 N_GND_M1004_b N_QN_c_1156_n 0.00102655f $X=-0.045 $Y=0 $X2=6.115 $Y2=2.96
cc_161 N_GND_M1004_b N_QN_c_1157_n 0.0133445f $X=-0.045 $Y=0 $X2=6.615 $Y2=1.85
cc_162 N_GND_c_119_p N_QN_c_1157_n 0.00827206f $X=6.545 $Y=0.825 $X2=6.615
+ $Y2=1.85
cc_163 N_GND_M1004_b N_QN_c_1159_n 0.00262941f $X=-0.045 $Y=0 $X2=6.2 $Y2=1.85
cc_164 N_GND_M1004_b N_QN_c_1160_n 0.0138424f $X=-0.045 $Y=0 $X2=6.615 $Y2=2.765
cc_165 N_GND_M1004_b N_QN_c_1161_n 0.00318212f $X=-0.045 $Y=0 $X2=6.2 $Y2=2.765
cc_166 N_GND_M1004_b N_QN_c_1162_n 0.0034889f $X=-0.045 $Y=0 $X2=6.7 $Y2=2.395
cc_167 N_GND_M1004_b QN 0.00252171f $X=-0.045 $Y=0 $X2=6.12 $Y2=2.96
cc_168 N_GND_M1004_b N_Q_c_1227_n 0.00913846f $X=-0.045 $Y=0 $X2=6.975 $Y2=0.825
cc_169 N_GND_c_4_p N_Q_c_1227_n 0.00476261f $X=6.46 $Y=0.19 $X2=6.975 $Y2=0.825
cc_170 N_GND_M1004_b N_Q_c_1229_n 0.0620687f $X=-0.045 $Y=0 $X2=7.09 $Y2=3.16
cc_171 N_GND_M1004_b N_Q_c_1230_n 0.0146196f $X=-0.045 $Y=0 $X2=7.09 $Y2=1.52
cc_172 N_VDD_M1020_b N_A_75_344#_M1020_g 0.0224266f $X=-0.045 $Y=2.905 $X2=0.5
+ $Y2=4.585
cc_173 N_VDD_c_173_p N_A_75_344#_M1020_g 0.00606474f $X=0.63 $Y=6.507 $X2=0.5
+ $Y2=4.585
cc_174 N_VDD_c_174_p N_A_75_344#_M1020_g 0.00354579f $X=0.715 $Y=3.795 $X2=0.5
+ $Y2=4.585
cc_175 N_VDD_c_175_p N_A_75_344#_M1020_g 0.00468827f $X=6.46 $Y=6.47 $X2=0.5
+ $Y2=4.585
cc_176 N_VDD_M1020_b N_A_75_344#_c_276_n 0.00631278f $X=-0.045 $Y=2.905 $X2=0.51
+ $Y2=2.765
cc_177 N_VDD_M1020_b N_A_75_344#_c_293_n 0.00145465f $X=-0.045 $Y=2.905
+ $X2=0.625 $Y2=3.1
cc_178 N_VDD_M1020_d N_A_75_344#_c_294_n 0.00447048f $X=0.575 $Y=3.085 $X2=1.42
+ $Y2=3.185
cc_179 N_VDD_c_174_p N_A_75_344#_c_294_n 0.00499116f $X=0.715 $Y=3.795 $X2=1.42
+ $Y2=3.185
cc_180 N_VDD_M1020_d N_A_75_344#_c_296_n 0.00106276f $X=0.575 $Y=3.085 $X2=0.71
+ $Y2=3.185
cc_181 N_VDD_c_174_p N_A_75_344#_c_296_n 0.00488762f $X=0.715 $Y=3.795 $X2=0.71
+ $Y2=3.185
cc_182 N_VDD_M1020_b N_A_75_344#_c_298_n 0.00313975f $X=-0.045 $Y=2.905 $X2=1.59
+ $Y2=3.455
cc_183 N_VDD_c_183_p N_A_75_344#_c_298_n 0.0149076f $X=2.38 $Y=6.507 $X2=1.59
+ $Y2=3.455
cc_184 N_VDD_c_175_p N_A_75_344#_c_298_n 0.00958198f $X=6.46 $Y=6.47 $X2=1.59
+ $Y2=3.455
cc_185 N_VDD_M1020_b N_A_75_344#_c_286_n 2.30281e-19 $X=-0.045 $Y=2.905 $X2=0.51
+ $Y2=2.765
cc_186 N_VDD_M1020_b N_D_M1007_g 0.0196478f $X=-0.045 $Y=2.905 $X2=0.93
+ $Y2=4.585
cc_187 N_VDD_c_174_p N_D_M1007_g 0.00354579f $X=0.715 $Y=3.795 $X2=0.93
+ $Y2=4.585
cc_188 N_VDD_c_183_p N_D_M1007_g 0.00606474f $X=2.38 $Y=6.507 $X2=0.93 $Y2=4.585
cc_189 N_VDD_c_175_p N_D_M1007_g 0.00468827f $X=6.46 $Y=6.47 $X2=0.93 $Y2=4.585
cc_190 N_VDD_M1020_b N_CK_M1009_g 0.0201249f $X=-0.045 $Y=2.905 $X2=1.29
+ $Y2=4.585
cc_191 N_VDD_c_183_p N_CK_M1009_g 0.00606474f $X=2.38 $Y=6.507 $X2=1.29
+ $Y2=4.585
cc_192 N_VDD_c_175_p N_CK_M1009_g 0.00468827f $X=6.46 $Y=6.47 $X2=1.29 $Y2=4.585
cc_193 N_VDD_M1020_b N_CK_M1012_g 0.020128f $X=-0.045 $Y=2.905 $X2=3.64
+ $Y2=4.585
cc_194 N_VDD_c_194_p N_CK_M1012_g 0.00606474f $X=4.13 $Y=6.507 $X2=3.64
+ $Y2=4.585
cc_195 N_VDD_c_175_p N_CK_M1012_g 0.00468827f $X=6.46 $Y=6.47 $X2=3.64 $Y2=4.585
cc_196 N_VDD_M1020_b N_CK_c_400_n 0.00774555f $X=-0.045 $Y=2.905 $X2=4.43
+ $Y2=2.93
cc_197 N_VDD_M1020_b N_CK_M1017_g 0.0214648f $X=-0.045 $Y=2.905 $X2=4.43
+ $Y2=4.585
cc_198 N_VDD_c_198_p N_CK_M1017_g 0.00354579f $X=4.215 $Y=3.455 $X2=4.43
+ $Y2=4.585
cc_199 N_VDD_c_199_p N_CK_M1017_g 0.00606474f $X=5.08 $Y=6.507 $X2=4.43
+ $Y2=4.585
cc_200 N_VDD_c_200_p N_CK_M1017_g 0.00811856f $X=5.165 $Y=3.795 $X2=4.43
+ $Y2=4.585
cc_201 N_VDD_c_175_p N_CK_M1017_g 0.00468827f $X=6.46 $Y=6.47 $X2=4.43 $Y2=4.585
cc_202 N_VDD_M1020_b N_CK_c_402_n 0.00487085f $X=-0.045 $Y=2.905 $X2=1.35
+ $Y2=2.765
cc_203 N_VDD_M1020_b N_CK_c_411_n 0.00487051f $X=-0.045 $Y=2.905 $X2=3.58
+ $Y2=2.765
cc_204 N_VDD_M1020_b N_CK_c_423_n 0.00302835f $X=-0.045 $Y=2.905 $X2=4.575
+ $Y2=2.59
cc_205 N_VDD_M1020_b N_CK_c_424_n 6.42499e-19 $X=-0.045 $Y=2.905 $X2=1.35
+ $Y2=2.59
cc_206 N_VDD_M1020_b N_CK_c_425_n 0.0022456f $X=-0.045 $Y=2.905 $X2=3.58
+ $Y2=2.59
cc_207 N_VDD_c_198_p N_CK_c_428_n 0.00634153f $X=4.215 $Y=3.455 $X2=4.43
+ $Y2=2.59
cc_208 N_VDD_M1020_b N_A_32_115#_M1016_g 0.0192219f $X=-0.045 $Y=2.905 $X2=2.25
+ $Y2=4.585
cc_209 N_VDD_c_183_p N_A_32_115#_M1016_g 0.00606474f $X=2.38 $Y=6.507 $X2=2.25
+ $Y2=4.585
cc_210 N_VDD_c_210_p N_A_32_115#_M1016_g 0.00354579f $X=2.465 $Y=3.795 $X2=2.25
+ $Y2=4.585
cc_211 N_VDD_c_175_p N_A_32_115#_M1016_g 0.00468827f $X=6.46 $Y=6.47 $X2=2.25
+ $Y2=4.585
cc_212 N_VDD_c_210_p N_A_32_115#_c_620_n 8.24975e-19 $X=2.465 $Y=3.795 $X2=2.605
+ $Y2=2.765
cc_213 N_VDD_M1020_b N_A_32_115#_M1005_g 0.0181098f $X=-0.045 $Y=2.905 $X2=2.68
+ $Y2=4.585
cc_214 N_VDD_c_210_p N_A_32_115#_M1005_g 0.00354579f $X=2.465 $Y=3.795 $X2=2.68
+ $Y2=4.585
cc_215 N_VDD_c_194_p N_A_32_115#_M1005_g 0.00606474f $X=4.13 $Y=6.507 $X2=2.68
+ $Y2=4.585
cc_216 N_VDD_c_175_p N_A_32_115#_M1005_g 0.00468827f $X=6.46 $Y=6.47 $X2=2.68
+ $Y2=4.585
cc_217 N_VDD_M1020_b N_A_32_115#_c_626_n 0.0107523f $X=-0.045 $Y=2.905 $X2=0.17
+ $Y2=3.14
cc_218 N_VDD_M1020_b N_A_32_115#_c_647_n 0.00156053f $X=-0.045 $Y=2.905
+ $X2=0.285 $Y2=3.455
cc_219 N_VDD_c_173_p N_A_32_115#_c_647_n 0.00736239f $X=0.63 $Y=6.507 $X2=0.285
+ $Y2=3.455
cc_220 N_VDD_c_175_p N_A_32_115#_c_647_n 0.00476261f $X=6.46 $Y=6.47 $X2=0.285
+ $Y2=3.455
cc_221 N_VDD_M1020_b N_A_32_115#_c_630_n 0.00424346f $X=-0.045 $Y=2.905 $X2=2.42
+ $Y2=2.765
cc_222 N_VDD_c_210_p N_A_32_115#_c_630_n 0.004428f $X=2.465 $Y=3.795 $X2=2.42
+ $Y2=2.765
cc_223 N_VDD_M1020_b N_A_32_115#_c_652_n 0.010813f $X=-0.045 $Y=2.905 $X2=0.285
+ $Y2=3.242
cc_224 N_VDD_M1020_b N_A_243_89#_M1014_g 0.0215131f $X=-0.045 $Y=2.905 $X2=1.89
+ $Y2=4.585
cc_225 N_VDD_c_183_p N_A_243_89#_M1014_g 0.00606474f $X=2.38 $Y=6.507 $X2=1.89
+ $Y2=4.585
cc_226 N_VDD_c_175_p N_A_243_89#_M1014_g 0.00468827f $X=6.46 $Y=6.47 $X2=1.89
+ $Y2=4.585
cc_227 N_VDD_M1020_b N_A_243_89#_M1019_g 0.0214821f $X=-0.045 $Y=2.905 $X2=3.04
+ $Y2=4.585
cc_228 N_VDD_c_194_p N_A_243_89#_M1019_g 0.00606474f $X=4.13 $Y=6.507 $X2=3.04
+ $Y2=4.585
cc_229 N_VDD_c_175_p N_A_243_89#_M1019_g 0.00468827f $X=6.46 $Y=6.47 $X2=3.04
+ $Y2=4.585
cc_230 N_VDD_M1020_b N_A_243_89#_c_762_n 0.00156053f $X=-0.045 $Y=2.905
+ $X2=4.645 $Y2=3.455
cc_231 N_VDD_c_199_p N_A_243_89#_c_762_n 0.00749582f $X=5.08 $Y=6.507 $X2=4.645
+ $Y2=3.455
cc_232 N_VDD_c_200_p N_A_243_89#_c_762_n 0.108505f $X=5.165 $Y=3.795 $X2=4.645
+ $Y2=3.455
cc_233 N_VDD_c_175_p N_A_243_89#_c_762_n 0.00476261f $X=6.46 $Y=6.47 $X2=4.645
+ $Y2=3.455
cc_234 N_VDD_M1020_b N_A_243_89#_c_753_n 0.00551116f $X=-0.045 $Y=2.905
+ $X2=4.915 $Y2=3.1
cc_235 N_VDD_M1020_b N_A_243_89#_c_767_n 0.013496f $X=-0.045 $Y=2.905 $X2=4.915
+ $Y2=3.185
cc_236 N_VDD_M1020_b N_A_785_89#_M1001_g 0.0197647f $X=-0.045 $Y=2.905 $X2=4
+ $Y2=4.585
cc_237 N_VDD_c_194_p N_A_785_89#_M1001_g 0.00606474f $X=4.13 $Y=6.507 $X2=4
+ $Y2=4.585
cc_238 N_VDD_c_198_p N_A_785_89#_M1001_g 0.00354579f $X=4.215 $Y=3.455 $X2=4
+ $Y2=4.585
cc_239 N_VDD_c_175_p N_A_785_89#_M1001_g 0.00468827f $X=6.46 $Y=6.47 $X2=4
+ $Y2=4.585
cc_240 N_VDD_M1020_b N_A_785_89#_c_916_n 0.0289529f $X=-0.045 $Y=2.905 $X2=6.305
+ $Y2=3.005
cc_241 N_VDD_c_241_p N_A_785_89#_c_916_n 0.00606474f $X=6.46 $Y=6.507 $X2=6.305
+ $Y2=3.005
cc_242 N_VDD_c_242_p N_A_785_89#_c_916_n 0.00354579f $X=6.545 $Y=3.455 $X2=6.305
+ $Y2=3.005
cc_243 N_VDD_c_175_p N_A_785_89#_c_916_n 0.00468827f $X=6.46 $Y=6.47 $X2=6.305
+ $Y2=3.005
cc_244 N_VDD_M1020_b N_A_785_89#_c_921_n 0.00558439f $X=-0.045 $Y=2.905
+ $X2=5.595 $Y2=3.455
cc_245 N_VDD_c_241_p N_A_785_89#_c_921_n 0.0074445f $X=6.46 $Y=6.507 $X2=5.595
+ $Y2=3.455
cc_246 N_VDD_c_175_p N_A_785_89#_c_921_n 0.00476261f $X=6.46 $Y=6.47 $X2=5.595
+ $Y2=3.455
cc_247 N_VDD_M1020_b N_A_623_115#_M1023_g 0.0260072f $X=-0.045 $Y=2.905 $X2=5.38
+ $Y2=4.585
cc_248 N_VDD_c_200_p N_A_623_115#_M1023_g 0.00713292f $X=5.165 $Y=3.795 $X2=5.38
+ $Y2=4.585
cc_249 N_VDD_c_241_p N_A_623_115#_M1023_g 0.00606474f $X=6.46 $Y=6.507 $X2=5.38
+ $Y2=4.585
cc_250 N_VDD_c_175_p N_A_623_115#_M1023_g 0.00468827f $X=6.46 $Y=6.47 $X2=5.38
+ $Y2=4.585
cc_251 N_VDD_M1020_b N_A_623_115#_c_1040_n 0.00168314f $X=-0.045 $Y=2.905
+ $X2=2.76 $Y2=1.85
cc_252 N_VDD_M1020_b N_A_623_115#_c_1056_n 0.00313975f $X=-0.045 $Y=2.905
+ $X2=3.34 $Y2=3.455
cc_253 N_VDD_c_194_p N_A_623_115#_c_1056_n 0.0151257f $X=4.13 $Y=6.507 $X2=3.34
+ $Y2=3.455
cc_254 N_VDD_c_175_p N_A_623_115#_c_1056_n 0.00958198f $X=6.46 $Y=6.47 $X2=3.34
+ $Y2=3.455
cc_255 N_VDD_M1020_b N_QN_M1002_g 0.0248218f $X=-0.045 $Y=2.905 $X2=6.76
+ $Y2=4.585
cc_256 N_VDD_c_242_p N_QN_M1002_g 0.00354579f $X=6.545 $Y=3.455 $X2=6.76
+ $Y2=4.585
cc_257 N_VDD_c_257_p N_QN_M1002_g 0.00606474f $X=6.46 $Y=6.47 $X2=6.76 $Y2=4.585
cc_258 N_VDD_c_175_p N_QN_M1002_g 0.00468827f $X=6.46 $Y=6.47 $X2=6.76 $Y2=4.585
cc_259 N_VDD_M1020_b N_QN_c_1156_n 0.00531805f $X=-0.045 $Y=2.905 $X2=6.115
+ $Y2=2.96
cc_260 N_VDD_c_241_p N_QN_c_1156_n 0.00757793f $X=6.46 $Y=6.507 $X2=6.115
+ $Y2=2.96
cc_261 N_VDD_c_175_p N_QN_c_1156_n 0.00476261f $X=6.46 $Y=6.47 $X2=6.115
+ $Y2=2.96
cc_262 N_VDD_c_242_p N_QN_c_1160_n 0.00818856f $X=6.545 $Y=3.455 $X2=6.615
+ $Y2=2.765
cc_263 N_VDD_M1020_b QN 0.00991454f $X=-0.045 $Y=2.905 $X2=6.12 $Y2=2.96
cc_264 N_VDD_M1020_b N_Q_c_1231_n 0.00156053f $X=-0.045 $Y=2.905 $X2=6.975
+ $Y2=3.455
cc_265 N_VDD_c_257_p N_Q_c_1231_n 0.00757793f $X=6.46 $Y=6.47 $X2=6.975
+ $Y2=3.455
cc_266 N_VDD_c_175_p N_Q_c_1231_n 0.00476261f $X=6.46 $Y=6.47 $X2=6.975
+ $Y2=3.455
cc_267 N_VDD_M1020_b N_Q_c_1229_n 0.0120121f $X=-0.045 $Y=2.905 $X2=7.09
+ $Y2=3.16
cc_268 N_VDD_M1020_b N_Q_c_1235_n 0.00894341f $X=-0.045 $Y=2.905 $X2=7.09
+ $Y2=3.245
cc_269 N_VDD_M1020_b Q 0.0052671f $X=-0.045 $Y=2.905 $X2=6.975 $Y2=3.33
cc_270 N_VDD_c_242_p Q 0.00679667f $X=6.545 $Y=3.455 $X2=6.975 $Y2=3.33
cc_271 N_A_75_344#_M1004_g N_D_M1003_g 0.0292768f $X=0.5 $Y=1.075 $X2=0.93
+ $Y2=1.075
cc_272 N_A_75_344#_c_277_n N_D_M1003_g 0.022942f $X=0.51 $Y=2.6 $X2=0.93
+ $Y2=1.075
cc_273 N_A_75_344#_c_278_n N_D_M1003_g 0.0146235f $X=1.405 $Y=1.765 $X2=0.93
+ $Y2=1.075
cc_274 N_A_75_344#_c_287_n N_D_M1003_g 0.00557207f $X=0.567 $Y=2.6 $X2=0.93
+ $Y2=1.075
cc_275 N_A_75_344#_M1020_g N_D_M1007_g 0.0356418f $X=0.5 $Y=4.585 $X2=0.93
+ $Y2=4.585
cc_276 N_A_75_344#_c_276_n N_D_M1007_g 0.0194268f $X=0.51 $Y=2.765 $X2=0.93
+ $Y2=4.585
cc_277 N_A_75_344#_c_293_n N_D_M1007_g 0.00557207f $X=0.625 $Y=3.1 $X2=0.93
+ $Y2=4.585
cc_278 N_A_75_344#_c_294_n N_D_M1007_g 0.019095f $X=1.42 $Y=3.185 $X2=0.93
+ $Y2=4.585
cc_279 N_A_75_344#_c_278_n N_D_c_362_n 0.00207628f $X=1.405 $Y=1.765 $X2=0.99
+ $Y2=2.22
cc_280 N_A_75_344#_c_286_n N_D_c_362_n 0.00557207f $X=0.51 $Y=2.765 $X2=0.99
+ $Y2=2.22
cc_281 N_A_75_344#_c_278_n N_D_c_363_n 0.0086486f $X=1.405 $Y=1.765 $X2=0.99
+ $Y2=2.22
cc_282 N_A_75_344#_c_287_n N_D_c_363_n 0.0187793f $X=0.567 $Y=2.6 $X2=0.99
+ $Y2=2.22
cc_283 N_A_75_344#_c_278_n D 0.00200799f $X=1.405 $Y=1.765 $X2=0.99 $Y2=2.22
cc_284 N_A_75_344#_c_287_n D 0.007232f $X=0.567 $Y=2.6 $X2=0.99 $Y2=2.22
cc_285 N_A_75_344#_c_294_n N_CK_M1009_g 0.0153724f $X=1.42 $Y=3.185 $X2=1.29
+ $Y2=4.585
cc_286 N_A_75_344#_c_294_n N_CK_c_402_n 0.00150627f $X=1.42 $Y=3.185 $X2=1.35
+ $Y2=2.765
cc_287 N_A_75_344#_c_278_n N_CK_c_403_n 9.45214e-19 $X=1.405 $Y=1.765 $X2=1.83
+ $Y2=1.85
cc_288 N_A_75_344#_c_319_p N_CK_c_403_n 0.00212965f $X=1.582 $Y=1.415 $X2=1.83
+ $Y2=1.85
cc_289 N_A_75_344#_c_282_n N_CK_c_404_n 0.00540119f $X=1.49 $Y=1.68 $X2=1.83
+ $Y2=1.685
cc_290 N_A_75_344#_c_278_n N_CK_c_418_n 0.0019742f $X=1.405 $Y=1.765 $X2=1.745
+ $Y2=2.59
cc_291 N_A_75_344#_c_294_n N_CK_c_418_n 0.00904674f $X=1.42 $Y=3.185 $X2=1.745
+ $Y2=2.59
cc_292 N_A_75_344#_c_278_n N_CK_c_419_n 0.012316f $X=1.405 $Y=1.765 $X2=1.83
+ $Y2=1.85
cc_293 N_A_75_344#_c_319_p N_CK_c_419_n 6.63879e-19 $X=1.582 $Y=1.415 $X2=1.83
+ $Y2=1.85
cc_294 N_A_75_344#_c_278_n N_CK_c_424_n 0.00224444f $X=1.405 $Y=1.765 $X2=1.35
+ $Y2=2.59
cc_295 N_A_75_344#_c_294_n N_CK_c_424_n 0.0101098f $X=1.42 $Y=3.185 $X2=1.35
+ $Y2=2.59
cc_296 N_A_75_344#_c_287_n N_CK_c_424_n 0.0103407f $X=0.567 $Y=2.6 $X2=1.35
+ $Y2=2.59
cc_297 N_A_75_344#_c_294_n N_CK_c_426_n 0.00613532f $X=1.42 $Y=3.185 $X2=3.435
+ $Y2=2.59
cc_298 N_A_75_344#_c_294_n N_CK_c_427_n 0.00409373f $X=1.42 $Y=3.185 $X2=1.495
+ $Y2=2.59
cc_299 N_A_75_344#_c_287_n N_CK_c_427_n 0.00642105f $X=0.567 $Y=2.6 $X2=1.495
+ $Y2=2.59
cc_300 N_A_75_344#_M1020_g N_A_32_115#_c_626_n 0.00426681f $X=0.5 $Y=4.585
+ $X2=0.17 $Y2=3.14
cc_301 N_A_75_344#_c_277_n N_A_32_115#_c_626_n 0.0218335f $X=0.51 $Y=2.6
+ $X2=0.17 $Y2=3.14
cc_302 N_A_75_344#_c_293_n N_A_32_115#_c_626_n 0.00821014f $X=0.625 $Y=3.1
+ $X2=0.17 $Y2=3.14
cc_303 N_A_75_344#_c_296_n N_A_32_115#_c_626_n 0.00210835f $X=0.71 $Y=3.185
+ $X2=0.17 $Y2=3.14
cc_304 N_A_75_344#_c_286_n N_A_32_115#_c_626_n 0.0245251f $X=0.51 $Y=2.765
+ $X2=0.17 $Y2=3.14
cc_305 N_A_75_344#_c_287_n N_A_32_115#_c_626_n 0.0334082f $X=0.567 $Y=2.6
+ $X2=0.17 $Y2=3.14
cc_306 N_A_75_344#_M1004_g N_A_32_115#_c_627_n 0.0084512f $X=0.5 $Y=1.075
+ $X2=0.285 $Y2=0.825
cc_307 N_A_75_344#_M1004_g N_A_32_115#_c_631_n 0.00165831f $X=0.5 $Y=1.075
+ $X2=0.285 $Y2=1.85
cc_308 N_A_75_344#_c_275_n N_A_32_115#_c_631_n 0.00460749f $X=0.475 $Y=1.87
+ $X2=0.285 $Y2=1.85
cc_309 N_A_75_344#_c_280_n N_A_32_115#_c_631_n 0.0125535f $X=0.71 $Y=1.765
+ $X2=0.285 $Y2=1.85
cc_310 N_A_75_344#_c_287_n N_A_32_115#_c_631_n 0.00592135f $X=0.567 $Y=2.6
+ $X2=0.285 $Y2=1.85
cc_311 N_A_75_344#_c_275_n N_A_32_115#_c_634_n 0.0047054f $X=0.475 $Y=1.87
+ $X2=2.185 $Y2=1.85
cc_312 N_A_75_344#_c_277_n N_A_32_115#_c_634_n 0.0043937f $X=0.51 $Y=2.6
+ $X2=2.185 $Y2=1.85
cc_313 N_A_75_344#_c_278_n N_A_32_115#_c_634_n 0.0597111f $X=1.405 $Y=1.765
+ $X2=2.185 $Y2=1.85
cc_314 N_A_75_344#_c_280_n N_A_32_115#_c_634_n 0.00750079f $X=0.71 $Y=1.765
+ $X2=2.185 $Y2=1.85
cc_315 N_A_75_344#_c_287_n N_A_32_115#_c_634_n 0.0143756f $X=0.567 $Y=2.6
+ $X2=2.185 $Y2=1.85
cc_316 N_A_75_344#_c_319_p N_A_32_115#_c_634_n 0.00757997f $X=1.582 $Y=1.415
+ $X2=2.185 $Y2=1.85
cc_317 N_A_75_344#_c_275_n N_A_32_115#_c_636_n 0.00387046f $X=0.475 $Y=1.87
+ $X2=0.43 $Y2=1.85
cc_318 N_A_75_344#_c_277_n N_A_32_115#_c_636_n 0.00369116f $X=0.51 $Y=2.6
+ $X2=0.43 $Y2=1.85
cc_319 N_A_75_344#_c_280_n N_A_32_115#_c_636_n 8.15236e-19 $X=0.71 $Y=1.765
+ $X2=0.43 $Y2=1.85
cc_320 N_A_75_344#_c_287_n N_A_32_115#_c_636_n 8.59347e-19 $X=0.567 $Y=2.6
+ $X2=0.43 $Y2=1.85
cc_321 N_A_75_344#_c_278_n N_A_243_89#_c_728_n 0.0066768f $X=1.405 $Y=1.765
+ $X2=1.29 $Y2=1.685
cc_322 N_A_75_344#_c_282_n N_A_243_89#_c_728_n 0.00488189f $X=1.49 $Y=1.68
+ $X2=1.29 $Y2=1.685
cc_323 N_A_75_344#_c_278_n N_A_243_89#_c_731_n 0.00324141f $X=1.405 $Y=1.765
+ $X2=1.41 $Y2=2.225
cc_324 N_A_75_344#_c_278_n N_A_243_89#_c_739_n 0.00993431f $X=1.405 $Y=1.765
+ $X2=1.41 $Y2=1.76
cc_325 N_A_75_344#_c_294_n A_201_617# 0.00732587f $X=1.42 $Y=3.185 $X2=1.005
+ $Y2=3.085
cc_326 N_D_M1007_g N_CK_c_402_n 0.21477f $X=0.93 $Y=4.585 $X2=1.35 $Y2=2.765
cc_327 N_D_c_362_n N_CK_c_419_n 2.89615e-19 $X=0.99 $Y=2.22 $X2=1.83 $Y2=1.85
cc_328 N_D_c_363_n N_CK_c_419_n 0.00478177f $X=0.99 $Y=2.22 $X2=1.83 $Y2=1.85
cc_329 D N_CK_c_419_n 0.00551577f $X=0.99 $Y=2.22 $X2=1.83 $Y2=1.85
cc_330 N_D_M1007_g N_CK_c_424_n 0.0030898f $X=0.93 $Y=4.585 $X2=1.35 $Y2=2.59
cc_331 N_D_M1007_g N_CK_c_427_n 0.00515433f $X=0.93 $Y=4.585 $X2=1.495 $Y2=2.59
cc_332 D N_CK_c_427_n 0.00375733f $X=0.99 $Y=2.22 $X2=1.495 $Y2=2.59
cc_333 N_D_M1003_g N_A_32_115#_c_634_n 0.00223521f $X=0.93 $Y=1.075 $X2=2.185
+ $Y2=1.85
cc_334 N_D_c_362_n N_A_32_115#_c_634_n 7.9412e-19 $X=0.99 $Y=2.22 $X2=2.185
+ $Y2=1.85
cc_335 N_D_c_363_n N_A_32_115#_c_634_n 0.00111625f $X=0.99 $Y=2.22 $X2=2.185
+ $Y2=1.85
cc_336 D N_A_32_115#_c_634_n 0.0353362f $X=0.99 $Y=2.22 $X2=2.185 $Y2=1.85
cc_337 N_D_M1003_g N_A_243_89#_c_728_n 0.0833388f $X=0.93 $Y=1.075 $X2=1.29
+ $Y2=1.685
cc_338 N_D_M1003_g N_A_243_89#_c_731_n 0.00886317f $X=0.93 $Y=1.075 $X2=1.41
+ $Y2=2.225
cc_339 N_D_c_362_n N_A_243_89#_c_731_n 0.0210215f $X=0.99 $Y=2.22 $X2=1.41
+ $Y2=2.225
cc_340 N_D_c_363_n N_A_243_89#_c_731_n 0.00164409f $X=0.99 $Y=2.22 $X2=1.41
+ $Y2=2.225
cc_341 D N_A_243_89#_c_731_n 0.00342011f $X=0.99 $Y=2.22 $X2=1.41 $Y2=2.225
cc_342 D N_A_243_89#_c_733_n 4.62757e-19 $X=0.99 $Y=2.22 $X2=1.485 $Y2=2.3
cc_343 N_CK_c_404_n N_A_32_115#_M1013_g 0.0479031f $X=1.83 $Y=1.685 $X2=2.25
+ $Y2=1.075
cc_344 N_CK_c_419_n N_A_32_115#_M1013_g 0.00109079f $X=1.83 $Y=1.85 $X2=2.25
+ $Y2=1.075
cc_345 N_CK_c_407_n N_A_32_115#_c_617_n 0.0471402f $X=3.1 $Y=1.85 $X2=2.605
+ $Y2=1.85
cc_346 N_CK_c_403_n N_A_32_115#_c_619_n 0.0479031f $X=1.83 $Y=1.85 $X2=2.325
+ $Y2=1.85
cc_347 N_CK_c_426_n N_A_32_115#_c_620_n 0.00772879f $X=3.435 $Y=2.59 $X2=2.605
+ $Y2=2.765
cc_348 N_CK_c_426_n N_A_32_115#_c_621_n 0.00679967f $X=3.435 $Y=2.59 $X2=2.325
+ $Y2=2.765
cc_349 N_CK_c_408_n N_A_32_115#_M1015_g 0.0471402f $X=3.1 $Y=1.685 $X2=2.68
+ $Y2=1.075
cc_350 N_CK_c_420_n N_A_32_115#_M1015_g 3.67139e-19 $X=3.1 $Y=1.85 $X2=2.68
+ $Y2=1.075
cc_351 N_CK_c_403_n N_A_32_115#_c_630_n 7.30049e-19 $X=1.83 $Y=1.85 $X2=2.42
+ $Y2=2.765
cc_352 N_CK_c_418_n N_A_32_115#_c_630_n 0.00401809f $X=1.745 $Y=2.59 $X2=2.42
+ $Y2=2.765
cc_353 N_CK_c_419_n N_A_32_115#_c_630_n 0.0203851f $X=1.83 $Y=1.85 $X2=2.42
+ $Y2=2.765
cc_354 N_CK_c_426_n N_A_32_115#_c_630_n 0.0206884f $X=3.435 $Y=2.59 $X2=2.42
+ $Y2=2.765
cc_355 N_CK_c_403_n N_A_32_115#_c_632_n 7.18106e-19 $X=1.83 $Y=1.85 $X2=2.42
+ $Y2=1.85
cc_356 N_CK_c_419_n N_A_32_115#_c_632_n 0.00742068f $X=1.83 $Y=1.85 $X2=2.42
+ $Y2=1.85
cc_357 N_CK_c_426_n N_A_32_115#_c_632_n 0.00102309f $X=3.435 $Y=2.59 $X2=2.42
+ $Y2=1.85
cc_358 N_CK_c_403_n N_A_32_115#_c_634_n 0.00576782f $X=1.83 $Y=1.85 $X2=2.185
+ $Y2=1.85
cc_359 N_CK_c_418_n N_A_32_115#_c_634_n 0.00443421f $X=1.745 $Y=2.59 $X2=2.185
+ $Y2=1.85
cc_360 N_CK_c_419_n N_A_32_115#_c_634_n 0.0205082f $X=1.83 $Y=1.85 $X2=2.185
+ $Y2=1.85
cc_361 N_CK_c_424_n N_A_32_115#_c_634_n 7.12046e-19 $X=1.35 $Y=2.59 $X2=2.185
+ $Y2=1.85
cc_362 N_CK_c_427_n N_A_32_115#_c_634_n 0.0126164f $X=1.495 $Y=2.59 $X2=2.185
+ $Y2=1.85
cc_363 N_CK_c_403_n N_A_32_115#_c_698_n 3.3031e-19 $X=1.83 $Y=1.85 $X2=2.33
+ $Y2=1.85
cc_364 N_CK_c_419_n N_A_32_115#_c_698_n 0.00143592f $X=1.83 $Y=1.85 $X2=2.33
+ $Y2=1.85
cc_365 N_CK_c_426_n N_A_32_115#_c_698_n 0.0129652f $X=3.435 $Y=2.59 $X2=2.33
+ $Y2=1.85
cc_366 N_CK_c_404_n N_A_243_89#_c_728_n 0.023382f $X=1.83 $Y=1.685 $X2=1.29
+ $Y2=1.685
cc_367 N_CK_c_419_n N_A_243_89#_c_731_n 0.00613747f $X=1.83 $Y=1.85 $X2=1.41
+ $Y2=2.225
cc_368 N_CK_c_403_n N_A_243_89#_c_732_n 0.0183603f $X=1.83 $Y=1.85 $X2=1.815
+ $Y2=2.3
cc_369 N_CK_c_419_n N_A_243_89#_c_732_n 0.00630484f $X=1.83 $Y=1.85 $X2=1.815
+ $Y2=2.3
cc_370 N_CK_c_426_n N_A_243_89#_c_732_n 0.00613485f $X=3.435 $Y=2.59 $X2=1.815
+ $Y2=2.3
cc_371 N_CK_c_402_n N_A_243_89#_c_733_n 0.00904036f $X=1.35 $Y=2.765 $X2=1.485
+ $Y2=2.3
cc_372 N_CK_c_418_n N_A_243_89#_c_733_n 0.00878348f $X=1.745 $Y=2.59 $X2=1.485
+ $Y2=2.3
cc_373 N_CK_c_424_n N_A_243_89#_c_733_n 0.00109468f $X=1.35 $Y=2.59 $X2=1.485
+ $Y2=2.3
cc_374 N_CK_c_427_n N_A_243_89#_c_733_n 0.00137501f $X=1.495 $Y=2.59 $X2=1.485
+ $Y2=2.3
cc_375 N_CK_M1009_g N_A_243_89#_M1014_g 0.0612157f $X=1.29 $Y=4.585 $X2=1.89
+ $Y2=4.585
cc_376 N_CK_c_402_n N_A_243_89#_M1014_g 0.0128384f $X=1.35 $Y=2.765 $X2=1.89
+ $Y2=4.585
cc_377 N_CK_c_418_n N_A_243_89#_M1014_g 0.0081071f $X=1.745 $Y=2.59 $X2=1.89
+ $Y2=4.585
cc_378 N_CK_c_419_n N_A_243_89#_M1014_g 0.00478024f $X=1.83 $Y=1.85 $X2=1.89
+ $Y2=4.585
cc_379 N_CK_c_424_n N_A_243_89#_M1014_g 0.00184124f $X=1.35 $Y=2.59 $X2=1.89
+ $Y2=4.585
cc_380 N_CK_c_426_n N_A_243_89#_M1014_g 0.00938974f $X=3.435 $Y=2.59 $X2=1.89
+ $Y2=4.585
cc_381 N_CK_c_427_n N_A_243_89#_M1014_g 4.2e-19 $X=1.495 $Y=2.59 $X2=1.89
+ $Y2=4.585
cc_382 N_CK_c_426_n N_A_243_89#_c_735_n 0.00607908f $X=3.435 $Y=2.59 $X2=2.965
+ $Y2=2.3
cc_383 N_CK_M1012_g N_A_243_89#_M1019_g 0.0612221f $X=3.64 $Y=4.585 $X2=3.04
+ $Y2=4.585
cc_384 N_CK_c_411_n N_A_243_89#_M1019_g 0.0118393f $X=3.58 $Y=2.765 $X2=3.04
+ $Y2=4.585
cc_385 N_CK_c_420_n N_A_243_89#_M1019_g 0.00399495f $X=3.1 $Y=1.85 $X2=3.04
+ $Y2=4.585
cc_386 N_CK_c_422_n N_A_243_89#_M1019_g 0.00654233f $X=3.185 $Y=2.59 $X2=3.04
+ $Y2=4.585
cc_387 N_CK_c_425_n N_A_243_89#_M1019_g 0.00128351f $X=3.58 $Y=2.59 $X2=3.04
+ $Y2=4.585
cc_388 N_CK_c_426_n N_A_243_89#_M1019_g 0.00497421f $X=3.435 $Y=2.59 $X2=3.04
+ $Y2=4.585
cc_389 N_CK_c_429_n N_A_243_89#_M1019_g 4.2e-19 $X=3.725 $Y=2.59 $X2=3.04
+ $Y2=4.585
cc_390 N_CK_c_411_n N_A_243_89#_c_737_n 0.00904036f $X=3.58 $Y=2.765 $X2=3.445
+ $Y2=2.3
cc_391 N_CK_c_420_n N_A_243_89#_c_737_n 0.00909647f $X=3.1 $Y=1.85 $X2=3.445
+ $Y2=2.3
cc_392 N_CK_c_421_n N_A_243_89#_c_737_n 0.00924811f $X=3.495 $Y=2.59 $X2=3.445
+ $Y2=2.3
cc_393 N_CK_c_425_n N_A_243_89#_c_737_n 0.00102633f $X=3.58 $Y=2.59 $X2=3.445
+ $Y2=2.3
cc_394 N_CK_c_426_n N_A_243_89#_c_737_n 0.00613485f $X=3.435 $Y=2.59 $X2=3.445
+ $Y2=2.3
cc_395 N_CK_c_429_n N_A_243_89#_c_737_n 0.00137501f $X=3.725 $Y=2.59 $X2=3.445
+ $Y2=2.3
cc_396 N_CK_c_420_n N_A_243_89#_c_738_n 0.00649764f $X=3.1 $Y=1.85 $X2=3.52
+ $Y2=2.225
cc_397 N_CK_c_403_n N_A_243_89#_c_739_n 0.0216263f $X=1.83 $Y=1.85 $X2=1.41
+ $Y2=1.76
cc_398 N_CK_c_424_n N_A_243_89#_c_739_n 2.45465e-19 $X=1.35 $Y=2.59 $X2=1.41
+ $Y2=1.76
cc_399 N_CK_c_419_n N_A_243_89#_c_740_n 0.00568091f $X=1.83 $Y=1.85 $X2=1.89
+ $Y2=2.3
cc_400 N_CK_c_407_n N_A_243_89#_c_741_n 0.0183603f $X=3.1 $Y=1.85 $X2=3.04
+ $Y2=2.3
cc_401 N_CK_c_420_n N_A_243_89#_c_741_n 0.00436024f $X=3.1 $Y=1.85 $X2=3.04
+ $Y2=2.3
cc_402 N_CK_c_407_n N_A_243_89#_c_742_n 0.0220721f $X=3.1 $Y=1.85 $X2=3.58
+ $Y2=1.85
cc_403 N_CK_c_411_n N_A_243_89#_c_742_n 0.00227671f $X=3.58 $Y=2.765 $X2=3.58
+ $Y2=1.85
cc_404 N_CK_c_420_n N_A_243_89#_c_742_n 0.00131283f $X=3.1 $Y=1.85 $X2=3.58
+ $Y2=1.85
cc_405 N_CK_c_425_n N_A_243_89#_c_742_n 5.27321e-19 $X=3.58 $Y=2.59 $X2=3.58
+ $Y2=1.85
cc_406 N_CK_c_429_n N_A_243_89#_c_742_n 8.78837e-19 $X=3.725 $Y=2.59 $X2=3.58
+ $Y2=1.85
cc_407 N_CK_c_408_n N_A_243_89#_c_743_n 0.0263924f $X=3.1 $Y=1.685 $X2=3.58
+ $Y2=1.685
cc_408 N_CK_c_401_n N_A_243_89#_c_746_n 0.00592387f $X=4.485 $Y=2.6 $X2=4.56
+ $Y2=1.85
cc_409 N_CK_c_407_n N_A_243_89#_c_746_n 8.05876e-19 $X=3.1 $Y=1.85 $X2=4.56
+ $Y2=1.85
cc_410 N_CK_c_411_n N_A_243_89#_c_746_n 5.56676e-19 $X=3.58 $Y=2.765 $X2=4.56
+ $Y2=1.85
cc_411 N_CK_c_417_n N_A_243_89#_c_746_n 0.00762848f $X=4.457 $Y=1.835 $X2=4.56
+ $Y2=1.85
cc_412 N_CK_c_420_n N_A_243_89#_c_746_n 0.00853323f $X=3.1 $Y=1.85 $X2=4.56
+ $Y2=1.85
cc_413 N_CK_c_421_n N_A_243_89#_c_746_n 0.00132011f $X=3.495 $Y=2.59 $X2=4.56
+ $Y2=1.85
cc_414 N_CK_c_423_n N_A_243_89#_c_746_n 8.24249e-19 $X=4.575 $Y=2.59 $X2=4.56
+ $Y2=1.85
cc_415 N_CK_c_425_n N_A_243_89#_c_746_n 0.00261697f $X=3.58 $Y=2.59 $X2=4.56
+ $Y2=1.85
cc_416 N_CK_c_426_n N_A_243_89#_c_746_n 3.12599e-19 $X=3.435 $Y=2.59 $X2=4.56
+ $Y2=1.85
cc_417 N_CK_c_428_n N_A_243_89#_c_746_n 0.00341454f $X=4.43 $Y=2.59 $X2=4.56
+ $Y2=1.85
cc_418 N_CK_c_429_n N_A_243_89#_c_746_n 0.00221563f $X=3.725 $Y=2.59 $X2=4.56
+ $Y2=1.85
cc_419 N_CK_c_412_n N_A_243_89#_c_748_n 0.00940234f $X=4.457 $Y=1.685 $X2=4.645
+ $Y2=0.825
cc_420 N_CK_c_417_n N_A_243_89#_c_748_n 0.0022869f $X=4.457 $Y=1.835 $X2=4.645
+ $Y2=0.825
cc_421 N_CK_c_401_n N_A_243_89#_c_752_n 0.00595506f $X=4.485 $Y=2.6 $X2=4.645
+ $Y2=2.105
cc_422 N_CK_c_400_n N_A_243_89#_c_753_n 0.0033284f $X=4.43 $Y=2.93 $X2=4.915
+ $Y2=3.1
cc_423 N_CK_M1017_g N_A_243_89#_c_753_n 0.00491946f $X=4.43 $Y=4.585 $X2=4.915
+ $Y2=3.1
cc_424 N_CK_c_401_n N_A_243_89#_c_753_n 0.00747875f $X=4.485 $Y=2.6 $X2=4.915
+ $Y2=3.1
cc_425 N_CK_c_423_n N_A_243_89#_c_753_n 0.0288018f $X=4.575 $Y=2.59 $X2=4.915
+ $Y2=3.1
cc_426 CK N_A_243_89#_c_753_n 0.00851352f $X=4.575 $Y=2.59 $X2=4.915 $Y2=3.1
cc_427 N_CK_c_401_n N_A_243_89#_c_754_n 0.00114916f $X=4.485 $Y=2.6 $X2=4.645
+ $Y2=1.85
cc_428 N_CK_c_417_n N_A_243_89#_c_754_n 8.09104e-19 $X=4.457 $Y=1.835 $X2=4.645
+ $Y2=1.85
cc_429 N_CK_c_400_n N_A_243_89#_c_755_n 0.00157237f $X=4.43 $Y=2.93 $X2=4.915
+ $Y2=2.19
cc_430 N_CK_c_401_n N_A_243_89#_c_755_n 0.00436926f $X=4.485 $Y=2.6 $X2=4.915
+ $Y2=2.19
cc_431 N_CK_c_423_n N_A_243_89#_c_755_n 0.00529105f $X=4.575 $Y=2.59 $X2=4.915
+ $Y2=2.19
cc_432 CK N_A_243_89#_c_755_n 8.76467e-19 $X=4.575 $Y=2.59 $X2=4.915 $Y2=2.19
cc_433 N_CK_c_400_n N_A_243_89#_c_767_n 0.00260941f $X=4.43 $Y=2.93 $X2=4.915
+ $Y2=3.185
cc_434 N_CK_c_423_n N_A_243_89#_c_767_n 0.00706443f $X=4.575 $Y=2.59 $X2=4.915
+ $Y2=3.185
cc_435 CK N_A_243_89#_c_767_n 0.00259785f $X=4.575 $Y=2.59 $X2=4.915 $Y2=3.185
cc_436 N_CK_c_401_n N_A_785_89#_M1022_g 0.00697006f $X=4.485 $Y=2.6 $X2=4
+ $Y2=1.075
cc_437 N_CK_c_412_n N_A_785_89#_M1022_g 0.0278502f $X=4.457 $Y=1.685 $X2=4
+ $Y2=1.075
cc_438 N_CK_c_400_n N_A_785_89#_M1001_g 0.0287701f $X=4.43 $Y=2.93 $X2=4
+ $Y2=4.585
cc_439 N_CK_c_401_n N_A_785_89#_M1001_g 0.0175925f $X=4.485 $Y=2.6 $X2=4
+ $Y2=4.585
cc_440 N_CK_c_411_n N_A_785_89#_M1001_g 0.214863f $X=3.58 $Y=2.765 $X2=4
+ $Y2=4.585
cc_441 N_CK_c_423_n N_A_785_89#_M1001_g 0.0026346f $X=4.575 $Y=2.59 $X2=4
+ $Y2=4.585
cc_442 N_CK_c_425_n N_A_785_89#_M1001_g 0.00453616f $X=3.58 $Y=2.59 $X2=4
+ $Y2=4.585
cc_443 N_CK_c_428_n N_A_785_89#_M1001_g 0.0114893f $X=4.43 $Y=2.59 $X2=4
+ $Y2=4.585
cc_444 N_CK_c_429_n N_A_785_89#_M1001_g 0.00113587f $X=3.725 $Y=2.59 $X2=4
+ $Y2=4.585
cc_445 CK N_A_785_89#_M1001_g 3.05655e-19 $X=4.575 $Y=2.59 $X2=4 $Y2=4.585
cc_446 N_CK_c_401_n N_A_785_89#_c_907_n 0.0213817f $X=4.485 $Y=2.6 $X2=4.06
+ $Y2=2.19
cc_447 N_CK_c_428_n N_A_785_89#_c_907_n 0.00185875f $X=4.43 $Y=2.59 $X2=4.06
+ $Y2=2.19
cc_448 N_CK_c_401_n N_A_785_89#_c_917_n 8.95026e-19 $X=4.485 $Y=2.6 $X2=4.06
+ $Y2=2.19
cc_449 N_CK_c_428_n N_A_785_89#_c_917_n 0.00488871f $X=4.43 $Y=2.59 $X2=4.06
+ $Y2=2.19
cc_450 N_CK_c_400_n N_A_785_89#_c_924_n 2.34467e-19 $X=4.43 $Y=2.93 $X2=6.07
+ $Y2=2.19
cc_451 N_CK_c_401_n N_A_785_89#_c_924_n 0.0033485f $X=4.485 $Y=2.6 $X2=6.07
+ $Y2=2.19
cc_452 N_CK_c_423_n N_A_785_89#_c_924_n 8.38639e-19 $X=4.575 $Y=2.59 $X2=6.07
+ $Y2=2.19
cc_453 N_CK_c_428_n N_A_785_89#_c_924_n 0.0179446f $X=4.43 $Y=2.59 $X2=6.07
+ $Y2=2.19
cc_454 CK N_A_785_89#_c_924_n 0.0248956f $X=4.575 $Y=2.59 $X2=6.07 $Y2=2.19
cc_455 N_CK_c_401_n N_A_785_89#_c_925_n 8.66236e-19 $X=4.485 $Y=2.6 $X2=4.205
+ $Y2=2.19
cc_456 N_CK_c_428_n N_A_785_89#_c_925_n 0.0247156f $X=4.43 $Y=2.59 $X2=4.205
+ $Y2=2.19
cc_457 N_CK_c_400_n N_A_623_115#_M1023_g 0.00448096f $X=4.43 $Y=2.93 $X2=5.38
+ $Y2=4.585
cc_458 N_CK_c_417_n N_A_623_115#_c_1038_n 0.00662135f $X=4.457 $Y=1.835 $X2=5.38
+ $Y2=1.85
cc_459 N_CK_c_408_n N_A_623_115#_c_1040_n 0.00573412f $X=3.1 $Y=1.685 $X2=2.76
+ $Y2=1.85
cc_460 N_CK_c_420_n N_A_623_115#_c_1040_n 0.057541f $X=3.1 $Y=1.85 $X2=2.76
+ $Y2=1.85
cc_461 N_CK_c_422_n N_A_623_115#_c_1040_n 0.0116326f $X=3.185 $Y=2.59 $X2=2.76
+ $Y2=1.85
cc_462 N_CK_c_425_n N_A_623_115#_c_1040_n 0.00613815f $X=3.58 $Y=2.59 $X2=2.76
+ $Y2=1.85
cc_463 N_CK_c_426_n N_A_623_115#_c_1040_n 0.020361f $X=3.435 $Y=2.59 $X2=2.76
+ $Y2=1.85
cc_464 N_CK_c_429_n N_A_623_115#_c_1040_n 6.61118e-19 $X=3.725 $Y=2.59 $X2=2.76
+ $Y2=1.85
cc_465 N_CK_c_407_n N_A_623_115#_c_1067_n 0.00237125f $X=3.1 $Y=1.85 $X2=3.17
+ $Y2=1.43
cc_466 N_CK_c_408_n N_A_623_115#_c_1067_n 0.0151803f $X=3.1 $Y=1.685 $X2=3.17
+ $Y2=1.43
cc_467 N_CK_c_420_n N_A_623_115#_c_1067_n 0.0103829f $X=3.1 $Y=1.85 $X2=3.17
+ $Y2=1.43
cc_468 N_CK_c_411_n N_A_623_115#_c_1070_n 0.00150627f $X=3.58 $Y=2.765 $X2=3.17
+ $Y2=3.185
cc_469 N_CK_c_421_n N_A_623_115#_c_1070_n 0.00843004f $X=3.495 $Y=2.59 $X2=3.17
+ $Y2=3.185
cc_470 N_CK_c_422_n N_A_623_115#_c_1070_n 0.00323798f $X=3.185 $Y=2.59 $X2=3.17
+ $Y2=3.185
cc_471 N_CK_c_425_n N_A_623_115#_c_1070_n 0.00103871f $X=3.58 $Y=2.59 $X2=3.17
+ $Y2=3.185
cc_472 N_CK_c_426_n N_A_623_115#_c_1070_n 0.012754f $X=3.435 $Y=2.59 $X2=3.17
+ $Y2=3.185
cc_473 N_CK_c_429_n N_A_623_115#_c_1070_n 0.00146098f $X=3.725 $Y=2.59 $X2=3.17
+ $Y2=3.185
cc_474 N_CK_c_417_n N_A_623_115#_c_1044_n 3.50905e-19 $X=4.457 $Y=1.835
+ $X2=5.175 $Y2=1.85
cc_475 N_CK_c_401_n N_A_623_115#_c_1046_n 0.00128484f $X=4.485 $Y=2.6 $X2=5.03
+ $Y2=1.85
cc_476 N_CK_c_407_n N_A_623_115#_c_1046_n 0.00407483f $X=3.1 $Y=1.85 $X2=5.03
+ $Y2=1.85
cc_477 N_CK_c_417_n N_A_623_115#_c_1046_n 0.0082638f $X=4.457 $Y=1.835 $X2=5.03
+ $Y2=1.85
cc_478 N_CK_c_420_n N_A_623_115#_c_1046_n 0.0133835f $X=3.1 $Y=1.85 $X2=5.03
+ $Y2=1.85
cc_479 N_CK_c_421_n N_A_623_115#_c_1046_n 0.00451177f $X=3.495 $Y=2.59 $X2=5.03
+ $Y2=1.85
cc_480 N_CK_c_425_n N_A_623_115#_c_1046_n 6.39375e-19 $X=3.58 $Y=2.59 $X2=5.03
+ $Y2=1.85
cc_481 N_CK_c_429_n N_A_623_115#_c_1046_n 0.0144351f $X=3.725 $Y=2.59 $X2=5.03
+ $Y2=1.85
cc_482 N_CK_c_407_n N_A_623_115#_c_1048_n 9.79344e-19 $X=3.1 $Y=1.85 $X2=2.905
+ $Y2=1.85
cc_483 N_CK_c_420_n N_A_623_115#_c_1048_n 0.00180575f $X=3.1 $Y=1.85 $X2=2.905
+ $Y2=1.85
cc_484 N_CK_c_426_n N_A_623_115#_c_1048_n 0.0128239f $X=3.435 $Y=2.59 $X2=2.905
+ $Y2=1.85
cc_485 N_A_32_115#_c_634_n N_A_243_89#_c_731_n 0.00252532f $X=2.185 $Y=1.85
+ $X2=1.41 $Y2=2.225
cc_486 N_A_32_115#_c_634_n N_A_243_89#_c_732_n 0.00296105f $X=2.185 $Y=1.85
+ $X2=1.815 $Y2=2.3
cc_487 N_A_32_115#_c_621_n N_A_243_89#_M1014_g 0.215294f $X=2.325 $Y=2.765
+ $X2=1.89 $Y2=4.585
cc_488 N_A_32_115#_c_630_n N_A_243_89#_M1014_g 0.00486364f $X=2.42 $Y=2.765
+ $X2=1.89 $Y2=4.585
cc_489 N_A_32_115#_c_619_n N_A_243_89#_c_735_n 0.0342351f $X=2.325 $Y=1.85
+ $X2=2.965 $Y2=2.3
cc_490 N_A_32_115#_c_621_n N_A_243_89#_c_735_n 0.0307748f $X=2.325 $Y=2.765
+ $X2=2.965 $Y2=2.3
cc_491 N_A_32_115#_c_630_n N_A_243_89#_c_735_n 0.0113171f $X=2.42 $Y=2.765
+ $X2=2.965 $Y2=2.3
cc_492 N_A_32_115#_c_632_n N_A_243_89#_c_735_n 8.69982e-19 $X=2.42 $Y=1.85
+ $X2=2.965 $Y2=2.3
cc_493 N_A_32_115#_c_634_n N_A_243_89#_c_735_n 0.00486036f $X=2.185 $Y=1.85
+ $X2=2.965 $Y2=2.3
cc_494 N_A_32_115#_c_698_n N_A_243_89#_c_735_n 4.12801e-19 $X=2.33 $Y=1.85
+ $X2=2.965 $Y2=2.3
cc_495 N_A_32_115#_c_620_n N_A_243_89#_M1019_g 0.211921f $X=2.605 $Y=2.765
+ $X2=3.04 $Y2=4.585
cc_496 N_A_32_115#_M1013_g N_A_623_115#_c_1040_n 9.367e-19 $X=2.25 $Y=1.075
+ $X2=2.76 $Y2=1.85
cc_497 N_A_32_115#_M1016_g N_A_623_115#_c_1040_n 9.36754e-19 $X=2.25 $Y=4.585
+ $X2=2.76 $Y2=1.85
cc_498 N_A_32_115#_c_617_n N_A_623_115#_c_1040_n 0.0061959f $X=2.605 $Y=1.85
+ $X2=2.76 $Y2=1.85
cc_499 N_A_32_115#_c_620_n N_A_623_115#_c_1040_n 0.00738718f $X=2.605 $Y=2.765
+ $X2=2.76 $Y2=1.85
cc_500 N_A_32_115#_M1015_g N_A_623_115#_c_1040_n 0.00481f $X=2.68 $Y=1.075
+ $X2=2.76 $Y2=1.85
cc_501 N_A_32_115#_M1005_g N_A_623_115#_c_1040_n 0.00479454f $X=2.68 $Y=4.585
+ $X2=2.76 $Y2=1.85
cc_502 N_A_32_115#_c_630_n N_A_623_115#_c_1040_n 0.0702347f $X=2.42 $Y=2.765
+ $X2=2.76 $Y2=1.85
cc_503 N_A_32_115#_c_632_n N_A_623_115#_c_1040_n 0.0157315f $X=2.42 $Y=1.85
+ $X2=2.76 $Y2=1.85
cc_504 N_A_32_115#_c_698_n N_A_623_115#_c_1040_n 4.18442e-19 $X=2.33 $Y=1.85
+ $X2=2.76 $Y2=1.85
cc_505 N_A_32_115#_M1013_g N_A_623_115#_c_1096_n 9.13132e-19 $X=2.25 $Y=1.075
+ $X2=2.845 $Y2=1.43
cc_506 N_A_32_115#_M1015_g N_A_623_115#_c_1096_n 0.00974042f $X=2.68 $Y=1.075
+ $X2=2.845 $Y2=1.43
cc_507 N_A_32_115#_M1016_g N_A_623_115#_c_1098_n 9.13132e-19 $X=2.25 $Y=4.585
+ $X2=2.845 $Y2=3.185
cc_508 N_A_32_115#_M1005_g N_A_623_115#_c_1098_n 0.0096885f $X=2.68 $Y=4.585
+ $X2=2.845 $Y2=3.185
cc_509 N_A_32_115#_c_617_n N_A_623_115#_c_1048_n 0.00433812f $X=2.605 $Y=1.85
+ $X2=2.905 $Y2=1.85
cc_510 N_A_32_115#_c_632_n N_A_623_115#_c_1048_n 0.0012094f $X=2.42 $Y=1.85
+ $X2=2.905 $Y2=1.85
cc_511 N_A_32_115#_c_698_n N_A_623_115#_c_1048_n 0.0241863f $X=2.33 $Y=1.85
+ $X2=2.905 $Y2=1.85
cc_512 N_A_243_89#_c_738_n N_A_785_89#_M1022_g 0.0073696f $X=3.52 $Y=2.225 $X2=4
+ $Y2=1.075
cc_513 N_A_243_89#_c_743_n N_A_785_89#_M1022_g 0.0963878f $X=3.58 $Y=1.685 $X2=4
+ $Y2=1.075
cc_514 N_A_243_89#_c_746_n N_A_785_89#_M1022_g 0.0107575f $X=4.56 $Y=1.85 $X2=4
+ $Y2=1.075
cc_515 N_A_243_89#_c_737_n N_A_785_89#_c_907_n 0.0073696f $X=3.445 $Y=2.3
+ $X2=4.06 $Y2=2.19
cc_516 N_A_243_89#_c_746_n N_A_785_89#_c_907_n 0.00290516f $X=4.56 $Y=1.85
+ $X2=4.06 $Y2=2.19
cc_517 N_A_243_89#_c_755_n N_A_785_89#_c_907_n 2.96928e-19 $X=4.915 $Y=2.19
+ $X2=4.06 $Y2=2.19
cc_518 N_A_243_89#_c_738_n N_A_785_89#_c_917_n 0.0035305f $X=3.52 $Y=2.225
+ $X2=4.06 $Y2=2.19
cc_519 N_A_243_89#_c_746_n N_A_785_89#_c_917_n 0.0219931f $X=4.56 $Y=1.85
+ $X2=4.06 $Y2=2.19
cc_520 N_A_243_89#_c_755_n N_A_785_89#_c_917_n 0.00559532f $X=4.915 $Y=2.19
+ $X2=4.06 $Y2=2.19
cc_521 N_A_243_89#_c_753_n N_A_785_89#_c_921_n 0.0285298f $X=4.915 $Y=3.1
+ $X2=5.595 $Y2=3.455
cc_522 N_A_243_89#_c_755_n N_A_785_89#_c_923_n 0.0038132f $X=4.915 $Y=2.19
+ $X2=5.595 $Y2=2.19
cc_523 N_A_243_89#_c_746_n N_A_785_89#_c_924_n 0.00314603f $X=4.56 $Y=1.85
+ $X2=6.07 $Y2=2.19
cc_524 N_A_243_89#_c_752_n N_A_785_89#_c_924_n 6.94255e-19 $X=4.645 $Y=2.105
+ $X2=6.07 $Y2=2.19
cc_525 N_A_243_89#_c_753_n N_A_785_89#_c_924_n 0.00464833f $X=4.915 $Y=3.1
+ $X2=6.07 $Y2=2.19
cc_526 N_A_243_89#_c_755_n N_A_785_89#_c_924_n 0.0225447f $X=4.915 $Y=2.19
+ $X2=6.07 $Y2=2.19
cc_527 N_A_243_89#_c_738_n N_A_785_89#_c_925_n 9.14174e-19 $X=3.52 $Y=2.225
+ $X2=4.205 $Y2=2.19
cc_528 N_A_243_89#_c_746_n N_A_785_89#_c_925_n 0.0010261f $X=4.56 $Y=1.85
+ $X2=4.205 $Y2=2.19
cc_529 N_A_243_89#_c_752_n N_A_785_89#_c_925_n 0.00122156f $X=4.645 $Y=2.105
+ $X2=4.205 $Y2=2.19
cc_530 N_A_243_89#_c_748_n N_A_623_115#_c_1033_n 0.00777279f $X=4.645 $Y=0.825
+ $X2=5.38 $Y2=1.685
cc_531 N_A_243_89#_c_752_n N_A_623_115#_M1023_g 0.00201047f $X=4.645 $Y=2.105
+ $X2=5.38 $Y2=4.585
cc_532 N_A_243_89#_c_762_n N_A_623_115#_M1023_g 0.0113755f $X=4.645 $Y=3.455
+ $X2=5.38 $Y2=4.585
cc_533 N_A_243_89#_c_753_n N_A_623_115#_M1023_g 0.012583f $X=4.915 $Y=3.1
+ $X2=5.38 $Y2=4.585
cc_534 N_A_243_89#_c_755_n N_A_623_115#_M1023_g 0.0023936f $X=4.915 $Y=2.19
+ $X2=5.38 $Y2=4.585
cc_535 N_A_243_89#_c_767_n N_A_623_115#_M1023_g 0.00340068f $X=4.915 $Y=3.185
+ $X2=5.38 $Y2=4.585
cc_536 N_A_243_89#_c_748_n N_A_623_115#_c_1038_n 0.00153999f $X=4.645 $Y=0.825
+ $X2=5.38 $Y2=1.85
cc_537 N_A_243_89#_c_752_n N_A_623_115#_c_1038_n 0.00153999f $X=4.645 $Y=2.105
+ $X2=5.38 $Y2=1.85
cc_538 N_A_243_89#_c_754_n N_A_623_115#_c_1038_n 5.35151e-19 $X=4.645 $Y=1.85
+ $X2=5.38 $Y2=1.85
cc_539 N_A_243_89#_c_735_n N_A_623_115#_c_1040_n 0.0124213f $X=2.965 $Y=2.3
+ $X2=2.76 $Y2=1.85
cc_540 N_A_243_89#_M1019_g N_A_623_115#_c_1040_n 0.0111407f $X=3.04 $Y=4.585
+ $X2=2.76 $Y2=1.85
cc_541 N_A_243_89#_c_742_n N_A_623_115#_c_1067_n 0.00183061f $X=3.58 $Y=1.85
+ $X2=3.17 $Y2=1.43
cc_542 N_A_243_89#_c_746_n N_A_623_115#_c_1067_n 0.00435378f $X=4.56 $Y=1.85
+ $X2=3.17 $Y2=1.43
cc_543 N_A_243_89#_M1019_g N_A_623_115#_c_1070_n 0.0162544f $X=3.04 $Y=4.585
+ $X2=3.17 $Y2=3.185
cc_544 N_A_243_89#_c_754_n N_A_623_115#_c_1044_n 0.00755683f $X=4.645 $Y=1.85
+ $X2=5.175 $Y2=1.85
cc_545 N_A_243_89#_c_735_n N_A_623_115#_c_1046_n 0.00156696f $X=2.965 $Y=2.3
+ $X2=5.03 $Y2=1.85
cc_546 N_A_243_89#_c_737_n N_A_623_115#_c_1046_n 0.00244106f $X=3.445 $Y=2.3
+ $X2=5.03 $Y2=1.85
cc_547 N_A_243_89#_c_741_n N_A_623_115#_c_1046_n 5.19983e-19 $X=3.04 $Y=2.3
+ $X2=5.03 $Y2=1.85
cc_548 N_A_243_89#_c_742_n N_A_623_115#_c_1046_n 0.0113766f $X=3.58 $Y=1.85
+ $X2=5.03 $Y2=1.85
cc_549 N_A_243_89#_c_746_n N_A_623_115#_c_1046_n 0.0492477f $X=4.56 $Y=1.85
+ $X2=5.03 $Y2=1.85
cc_550 N_A_243_89#_c_754_n N_A_623_115#_c_1046_n 0.0171747f $X=4.645 $Y=1.85
+ $X2=5.03 $Y2=1.85
cc_551 N_A_243_89#_c_755_n N_A_623_115#_c_1046_n 0.00219678f $X=4.915 $Y=2.19
+ $X2=5.03 $Y2=1.85
cc_552 N_A_243_89#_c_735_n N_A_623_115#_c_1048_n 0.00120486f $X=2.965 $Y=2.3
+ $X2=2.905 $Y2=1.85
cc_553 N_A_243_89#_c_748_n N_A_623_115#_c_1049_n 0.00126742f $X=4.645 $Y=0.825
+ $X2=5.175 $Y2=1.85
cc_554 N_A_243_89#_c_752_n N_A_623_115#_c_1049_n 0.00126742f $X=4.645 $Y=2.105
+ $X2=5.175 $Y2=1.85
cc_555 N_A_785_89#_c_918_n N_A_623_115#_c_1033_n 0.0235974f $X=5.595 $Y=0.825
+ $X2=5.38 $Y2=1.685
cc_556 N_A_785_89#_c_908_n N_A_623_115#_M1023_g 0.0046172f $X=6.215 $Y=2.19
+ $X2=5.38 $Y2=4.585
cc_557 N_A_785_89#_c_921_n N_A_623_115#_M1023_g 0.0248329f $X=5.595 $Y=3.455
+ $X2=5.38 $Y2=4.585
cc_558 N_A_785_89#_c_923_n N_A_623_115#_M1023_g 0.00245806f $X=5.595 $Y=2.19
+ $X2=5.38 $Y2=4.585
cc_559 N_A_785_89#_c_924_n N_A_623_115#_M1023_g 0.0167433f $X=6.07 $Y=2.19
+ $X2=5.38 $Y2=4.585
cc_560 N_A_785_89#_c_924_n N_A_623_115#_c_1038_n 0.0041429f $X=6.07 $Y=2.19
+ $X2=5.38 $Y2=1.85
cc_561 N_A_785_89#_c_918_n N_A_623_115#_c_1044_n 0.0115453f $X=5.595 $Y=0.825
+ $X2=5.175 $Y2=1.85
cc_562 N_A_785_89#_c_924_n N_A_623_115#_c_1044_n 0.00508416f $X=6.07 $Y=2.19
+ $X2=5.175 $Y2=1.85
cc_563 N_A_785_89#_M1022_g N_A_623_115#_c_1046_n 0.00707887f $X=4 $Y=1.075
+ $X2=5.03 $Y2=1.85
cc_564 N_A_785_89#_c_907_n N_A_623_115#_c_1046_n 0.00187603f $X=4.06 $Y=2.19
+ $X2=5.03 $Y2=1.85
cc_565 N_A_785_89#_c_917_n N_A_623_115#_c_1046_n 0.00166223f $X=4.06 $Y=2.19
+ $X2=5.03 $Y2=1.85
cc_566 N_A_785_89#_c_924_n N_A_623_115#_c_1046_n 0.0735565f $X=6.07 $Y=2.19
+ $X2=5.03 $Y2=1.85
cc_567 N_A_785_89#_c_925_n N_A_623_115#_c_1046_n 0.0289631f $X=4.205 $Y=2.19
+ $X2=5.03 $Y2=1.85
cc_568 N_A_785_89#_c_918_n N_A_623_115#_c_1049_n 0.00389142f $X=5.595 $Y=0.825
+ $X2=5.175 $Y2=1.85
cc_569 N_A_785_89#_c_924_n N_A_623_115#_c_1049_n 0.0291144f $X=6.07 $Y=2.19
+ $X2=5.175 $Y2=1.85
cc_570 N_A_785_89#_c_909_n N_QN_M1025_g 0.0153129f $X=6.217 $Y=2.025 $X2=6.76
+ $Y2=1.075
cc_571 N_A_785_89#_c_910_n N_QN_M1025_g 0.0248825f $X=6.305 $Y=1.65 $X2=6.76
+ $Y2=1.075
cc_572 N_A_785_89#_c_922_n N_QN_M1025_g 4.79563e-19 $X=6.215 $Y=2.19 $X2=6.76
+ $Y2=1.075
cc_573 N_A_785_89#_c_915_n N_QN_M1002_g 0.0102953f $X=6.305 $Y=2.855 $X2=6.76
+ $Y2=4.585
cc_574 N_A_785_89#_c_916_n N_QN_M1002_g 0.0234784f $X=6.305 $Y=3.005 $X2=6.76
+ $Y2=4.585
cc_575 N_A_785_89#_c_908_n N_QN_c_1152_n 0.021196f $X=6.215 $Y=2.19 $X2=6.7
+ $Y2=2.395
cc_576 N_A_785_89#_c_922_n N_QN_c_1152_n 3.0115e-19 $X=6.215 $Y=2.19 $X2=6.7
+ $Y2=2.395
cc_577 N_A_785_89#_c_926_n N_QN_c_1152_n 4.60229e-19 $X=6.215 $Y=2.19 $X2=6.7
+ $Y2=2.395
cc_578 N_A_785_89#_c_910_n N_QN_c_1153_n 0.00804393f $X=6.305 $Y=1.65 $X2=6.115
+ $Y2=0.825
cc_579 N_A_785_89#_c_914_n N_QN_c_1153_n 0.00485394f $X=6.305 $Y=1.8 $X2=6.115
+ $Y2=0.825
cc_580 N_A_785_89#_c_918_n N_QN_c_1153_n 0.0513779f $X=5.595 $Y=0.825 $X2=6.115
+ $Y2=0.825
cc_581 N_A_785_89#_c_915_n N_QN_c_1156_n 0.00567875f $X=6.305 $Y=2.855 $X2=6.115
+ $Y2=2.96
cc_582 N_A_785_89#_c_916_n N_QN_c_1156_n 0.00708078f $X=6.305 $Y=3.005 $X2=6.115
+ $Y2=2.96
cc_583 N_A_785_89#_c_921_n N_QN_c_1156_n 0.135407f $X=5.595 $Y=3.455 $X2=6.115
+ $Y2=2.96
cc_584 N_A_785_89#_c_909_n N_QN_c_1157_n 0.00799433f $X=6.217 $Y=2.025 $X2=6.615
+ $Y2=1.85
cc_585 N_A_785_89#_c_914_n N_QN_c_1157_n 0.011031f $X=6.305 $Y=1.8 $X2=6.615
+ $Y2=1.85
cc_586 N_A_785_89#_c_922_n N_QN_c_1157_n 0.0110498f $X=6.215 $Y=2.19 $X2=6.615
+ $Y2=1.85
cc_587 N_A_785_89#_c_926_n N_QN_c_1157_n 0.00387586f $X=6.215 $Y=2.19 $X2=6.615
+ $Y2=1.85
cc_588 N_A_785_89#_c_908_n N_QN_c_1159_n 0.00308111f $X=6.215 $Y=2.19 $X2=6.2
+ $Y2=1.85
cc_589 N_A_785_89#_c_918_n N_QN_c_1159_n 0.00869401f $X=5.595 $Y=0.825 $X2=6.2
+ $Y2=1.85
cc_590 N_A_785_89#_c_922_n N_QN_c_1159_n 0.0120703f $X=6.215 $Y=2.19 $X2=6.2
+ $Y2=1.85
cc_591 N_A_785_89#_c_924_n N_QN_c_1159_n 0.0010572f $X=6.07 $Y=2.19 $X2=6.2
+ $Y2=1.85
cc_592 N_A_785_89#_c_926_n N_QN_c_1159_n 0.00336135f $X=6.215 $Y=2.19 $X2=6.2
+ $Y2=1.85
cc_593 N_A_785_89#_c_915_n N_QN_c_1160_n 0.016126f $X=6.305 $Y=2.855 $X2=6.615
+ $Y2=2.765
cc_594 N_A_785_89#_c_916_n N_QN_c_1160_n 0.00248624f $X=6.305 $Y=3.005 $X2=6.615
+ $Y2=2.765
cc_595 N_A_785_89#_c_922_n N_QN_c_1160_n 0.00426371f $X=6.215 $Y=2.19 $X2=6.615
+ $Y2=2.765
cc_596 N_A_785_89#_c_926_n N_QN_c_1160_n 0.00253233f $X=6.215 $Y=2.19 $X2=6.615
+ $Y2=2.765
cc_597 N_A_785_89#_c_908_n N_QN_c_1161_n 0.00265611f $X=6.215 $Y=2.19 $X2=6.2
+ $Y2=2.765
cc_598 N_A_785_89#_c_921_n N_QN_c_1161_n 0.00859877f $X=5.595 $Y=3.455 $X2=6.2
+ $Y2=2.765
cc_599 N_A_785_89#_c_922_n N_QN_c_1161_n 0.00471962f $X=6.215 $Y=2.19 $X2=6.2
+ $Y2=2.765
cc_600 N_A_785_89#_c_924_n N_QN_c_1161_n 9.40773e-19 $X=6.07 $Y=2.19 $X2=6.2
+ $Y2=2.765
cc_601 N_A_785_89#_c_926_n N_QN_c_1161_n 0.00140341f $X=6.215 $Y=2.19 $X2=6.2
+ $Y2=2.765
cc_602 N_A_785_89#_c_908_n N_QN_c_1162_n 0.00216137f $X=6.215 $Y=2.19 $X2=6.7
+ $Y2=2.395
cc_603 N_A_785_89#_c_909_n N_QN_c_1162_n 0.00323473f $X=6.217 $Y=2.025 $X2=6.7
+ $Y2=2.395
cc_604 N_A_785_89#_c_915_n N_QN_c_1162_n 0.00226435f $X=6.305 $Y=2.855 $X2=6.7
+ $Y2=2.395
cc_605 N_A_785_89#_c_922_n N_QN_c_1162_n 0.00987106f $X=6.215 $Y=2.19 $X2=6.7
+ $Y2=2.395
cc_606 N_A_785_89#_c_926_n N_QN_c_1162_n 0.00377439f $X=6.215 $Y=2.19 $X2=6.7
+ $Y2=2.395
cc_607 N_A_785_89#_c_916_n QN 0.00740862f $X=6.305 $Y=3.005 $X2=6.12 $Y2=2.96
cc_608 N_A_785_89#_c_921_n QN 0.00717604f $X=5.595 $Y=3.455 $X2=6.12 $Y2=2.96
cc_609 N_A_785_89#_c_922_n QN 0.00350993f $X=6.215 $Y=2.19 $X2=6.12 $Y2=2.96
cc_610 N_A_785_89#_c_926_n QN 0.00842298f $X=6.215 $Y=2.19 $X2=6.12 $Y2=2.96
cc_611 N_A_623_115#_c_1070_n A_551_617# 0.00342591f $X=3.17 $Y=3.185 $X2=2.755
+ $Y2=3.085
cc_612 N_A_623_115#_c_1098_n A_551_617# 0.00144354f $X=2.845 $Y=3.185 $X2=2.755
+ $Y2=3.085
cc_613 N_A_623_115#_c_1040_n A_551_115# 6.64472e-19 $X=2.76 $Y=1.85 $X2=2.755
+ $Y2=0.575
cc_614 N_A_623_115#_c_1067_n A_551_115# 0.00317038f $X=3.17 $Y=1.43 $X2=2.755
+ $Y2=0.575
cc_615 N_A_623_115#_c_1096_n A_551_115# 0.00148865f $X=2.845 $Y=1.43 $X2=2.755
+ $Y2=0.575
cc_616 N_QN_M1002_g N_Q_c_1231_n 0.00125257f $X=6.76 $Y=4.585 $X2=6.975
+ $Y2=3.455
cc_617 N_QN_M1025_g N_Q_c_1229_n 0.0380298f $X=6.76 $Y=1.075 $X2=7.09 $Y2=3.16
cc_618 N_QN_c_1157_n N_Q_c_1229_n 0.0111776f $X=6.615 $Y=1.85 $X2=7.09 $Y2=3.16
cc_619 N_QN_c_1160_n N_Q_c_1229_n 0.0111776f $X=6.615 $Y=2.765 $X2=7.09 $Y2=3.16
cc_620 N_QN_c_1162_n N_Q_c_1229_n 0.0438362f $X=6.7 $Y=2.395 $X2=7.09 $Y2=3.16
cc_621 N_QN_M1025_g N_Q_c_1230_n 0.00414595f $X=6.76 $Y=1.075 $X2=7.09 $Y2=1.52
cc_622 N_QN_M1002_g N_Q_c_1235_n 0.00198876f $X=6.76 $Y=4.585 $X2=7.09 $Y2=3.245
cc_623 N_QN_M1002_g Q 0.010705f $X=6.76 $Y=4.585 $X2=6.975 $Y2=3.33
cc_624 N_QN_c_1160_n Q 0.00245821f $X=6.615 $Y=2.765 $X2=6.975 $Y2=3.33
