* File: sky130_osu_sc_18T_ls__dffsr_1.pex.spice
* Created: Fri Nov 12 14:16:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%GND 1 2 3 4 5 6 7 8 9 127 131 133 140
+ 142 152 158 160 170 172 182 184 191 193 203 205 212 238 240
c248 191 0 1.63226e-19 $X=7.47 $Y=0.825
c249 182 0 1.67294e-19 $X=6.52 $Y=0.825
c250 158 0 3.07193e-19 $X=3.02 $Y=0.825
c251 152 0 2.98797e-19 $X=2.5 $Y=0.825
c252 140 0 1.90798e-19 $X=1.22 $Y=0.825
c253 127 0 1.91032e-19 $X=-0.05 $Y=0
r254 238 240 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.855 $Y2=0.152
r255 214 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=0.152
+ $X2=9.71 $Y2=0.152
r256 210 234 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.152
r257 210 212 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.825
r258 206 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.152
+ $X2=8.75 $Y2=0.152
r259 205 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=0.152
+ $X2=9.71 $Y2=0.152
r260 201 233 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.152
r261 201 203 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.825
r262 194 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.152
+ $X2=7.47 $Y2=0.152
r263 193 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.152
+ $X2=8.75 $Y2=0.152
r264 189 232 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.152
r265 189 191 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.825
r266 184 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=0.152
+ $X2=7.47 $Y2=0.152
r267 180 182 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.52 $Y=0.305
+ $X2=6.52 $Y2=0.825
r268 173 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.152
+ $X2=4.77 $Y2=0.152
r269 168 228 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.152
r270 168 170 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.825
r271 160 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.152
+ $X2=4.77 $Y2=0.152
r272 156 158 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.02 $Y=0.305
+ $X2=3.02 $Y2=0.825
r273 155 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.152
+ $X2=2.5 $Y2=0.152
r274 154 155 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=2.935 $Y=0.152
+ $X2=2.585 $Y2=0.152
r275 150 224 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.152
r276 150 152 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.825
r277 143 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0.152
+ $X2=1.22 $Y2=0.152
r278 142 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.152
+ $X2=2.5 $Y2=0.152
r279 138 223 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.152
r280 138 140 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.825
r281 133 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.152
+ $X2=1.22 $Y2=0.152
r282 129 131 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r283 127 240 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=0.19
+ $X2=9.855 $Y2=0.19
r284 127 238 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r285 127 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.52 $Y2=0.305
r286 127 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.435 $Y2=0.152
r287 127 185 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.605 $Y2=0.152
r288 127 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.02 $Y2=0.305
r289 127 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=2.935 $Y2=0.152
r290 127 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.105 $Y2=0.152
r291 127 129 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r292 127 134 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r293 127 214 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.855 $Y=0.152
+ $X2=9.795 $Y2=0.152
r294 127 205 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=9.625 $Y2=0.152
r295 127 206 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.835 $Y2=0.152
r296 127 193 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.665 $Y2=0.152
r297 127 194 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=7.815 $Y=0.152
+ $X2=7.555 $Y2=0.152
r298 127 184 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.385 $Y2=0.152
r299 127 185 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.605 $Y2=0.152
r300 127 172 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.435 $Y2=0.152
r301 127 173 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.855 $Y2=0.152
r302 127 160 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=4.685 $Y2=0.152
r303 127 161 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.105 $Y2=0.152
r304 127 142 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.415 $Y2=0.152
r305 127 143 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.305 $Y2=0.152
r306 127 133 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.135 $Y2=0.152
r307 127 134 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r308 9 212 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=9.57
+ $Y=0.575 $X2=9.71 $Y2=0.825
r309 8 203 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.61
+ $Y=0.575 $X2=8.75 $Y2=0.825
r310 7 191 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.825
r311 6 182 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.825
r312 5 170 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.575 $X2=4.77 $Y2=0.825
r313 4 158 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.575 $X2=3.02 $Y2=0.825
r314 3 152 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.5 $Y2=0.825
r315 2 140 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.575 $X2=1.22 $Y2=0.825
r316 1 131 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%VDD 1 2 3 4 5 6 7 89 93 97 105 109 115
+ 119 127 131 139 143 149 153 161 167 182 186
c145 161 0 1.98165e-19 $X=9.71 $Y=3.455
r146 182 186 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=6.507
+ $X2=9.855 $Y2=6.507
r147 170 182 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=6.47
+ $X2=0.335 $Y2=6.47
r148 167 186 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=6.47
+ $X2=9.855 $Y2=6.47
r149 165 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=6.507
+ $X2=9.71 $Y2=6.507
r150 165 167 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.795 $Y=6.507
+ $X2=9.855 $Y2=6.507
r151 161 164 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=9.71 $Y=3.455
+ $X2=9.71 $Y2=5.835
r152 159 180 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.71 $Y=6.355
+ $X2=9.71 $Y2=6.507
r153 159 164 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.71 $Y=6.355
+ $X2=9.71 $Y2=5.835
r154 156 158 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=8.495 $Y=6.507
+ $X2=9.175 $Y2=6.507
r155 154 179 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=6.507
+ $X2=7.9 $Y2=6.507
r156 154 156 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=7.985 $Y=6.507
+ $X2=8.495 $Y2=6.507
r157 153 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=6.507
+ $X2=9.71 $Y2=6.507
r158 153 158 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.625 $Y=6.507
+ $X2=9.175 $Y2=6.507
r159 149 152 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=5.835
r160 147 179 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=6.507
r161 147 152 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=5.835
r162 144 177 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=6.507
+ $X2=6.52 $Y2=6.507
r163 144 146 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=6.605 $Y=6.507
+ $X2=7.135 $Y2=6.507
r164 143 179 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.9 $Y2=6.507
r165 143 146 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.135 $Y2=6.507
r166 139 142 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.52 $Y=3.455
+ $X2=6.52 $Y2=5.835
r167 137 177 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.52 $Y=6.355
+ $X2=6.52 $Y2=6.507
r168 137 142 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.52 $Y=6.355
+ $X2=6.52 $Y2=5.835
r169 134 136 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=6.507
+ $X2=5.775 $Y2=6.507
r170 132 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=6.507
+ $X2=4.77 $Y2=6.507
r171 132 134 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=4.855 $Y=6.507
+ $X2=5.095 $Y2=6.507
r172 131 177 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=6.507
+ $X2=6.52 $Y2=6.507
r173 131 136 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=6.435 $Y=6.507
+ $X2=5.775 $Y2=6.507
r174 127 130 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.77 $Y=3.795
+ $X2=4.77 $Y2=5.835
r175 125 175 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.77 $Y=6.355
+ $X2=4.77 $Y2=6.507
r176 125 130 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.77 $Y=6.355
+ $X2=4.77 $Y2=5.835
r177 122 124 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=6.507
+ $X2=4.415 $Y2=6.507
r178 120 174 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=6.507
+ $X2=3.02 $Y2=6.507
r179 120 122 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.105 $Y=6.507
+ $X2=3.735 $Y2=6.507
r180 119 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=6.507
+ $X2=4.77 $Y2=6.507
r181 119 124 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.685 $Y=6.507
+ $X2=4.415 $Y2=6.507
r182 115 118 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=3.02 $Y=3.795
+ $X2=3.02 $Y2=5.835
r183 113 174 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.02 $Y=6.355
+ $X2=3.02 $Y2=6.507
r184 113 118 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.02 $Y=6.355
+ $X2=3.02 $Y2=5.835
r185 110 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=6.507
+ $X2=2.07 $Y2=6.507
r186 110 112 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.155 $Y=6.507
+ $X2=2.375 $Y2=6.507
r187 109 174 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=6.507
+ $X2=3.02 $Y2=6.507
r188 109 112 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=2.935 $Y=6.507
+ $X2=2.375 $Y2=6.507
r189 105 108 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.07 $Y=4.135
+ $X2=2.07 $Y2=5.835
r190 103 172 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.07 $Y=6.355
+ $X2=2.07 $Y2=6.507
r191 103 108 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.07 $Y=6.355
+ $X2=2.07 $Y2=5.835
r192 100 102 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=6.507
+ $X2=1.695 $Y2=6.507
r193 98 170 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r194 98 100 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.015 $Y2=6.507
r195 97 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=6.507
+ $X2=2.07 $Y2=6.507
r196 97 102 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.985 $Y=6.507
+ $X2=1.695 $Y2=6.507
r197 93 96 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r198 91 170 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r199 91 96 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r200 89 167 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=9.65 $Y=6.355 $X2=9.855 $Y2=6.44
r201 89 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=6.355 $X2=9.175 $Y2=6.44
r202 89 156 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=6.355 $X2=8.495 $Y2=6.44
r203 89 179 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=6.355 $X2=7.815 $Y2=6.44
r204 89 146 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=6.355 $X2=7.135 $Y2=6.44
r205 89 177 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=6.355 $X2=6.455 $Y2=6.44
r206 89 136 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=6.355 $X2=5.775 $Y2=6.44
r207 89 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=6.355 $X2=5.095 $Y2=6.44
r208 89 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=6.355 $X2=4.415 $Y2=6.44
r209 89 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=6.355 $X2=3.735 $Y2=6.44
r210 89 174 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=6.355 $X2=3.055 $Y2=6.44
r211 89 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=6.355 $X2=2.375 $Y2=6.44
r212 89 102 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=6.355 $X2=1.695 $Y2=6.44
r213 89 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=6.355 $X2=1.015 $Y2=6.44
r214 89 170 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=6.355 $X2=0.335 $Y2=6.44
r215 7 164 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=9.57
+ $Y=3.085 $X2=9.71 $Y2=5.835
r216 7 161 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=9.57
+ $Y=3.085 $X2=9.71 $Y2=3.455
r217 6 152 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=7.76
+ $Y=3.085 $X2=7.9 $Y2=5.835
r218 6 149 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=7.76
+ $Y=3.085 $X2=7.9 $Y2=4.135
r219 5 142 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=5.835
r220 5 139 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=3.455
r221 4 130 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=4.63 $Y=3.085 $X2=4.77 $Y2=5.835
r222 4 127 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=4.63 $Y=3.085 $X2=4.77 $Y2=3.795
r223 3 118 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=2.895 $Y=3.085 $X2=3.02 $Y2=5.835
r224 3 115 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=2.895 $Y=3.085 $X2=3.02 $Y2=3.795
r225 2 108 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=5.835
r226 2 105 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=1.93
+ $Y=3.085 $X2=2.07 $Y2=4.135
r227 1 96 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r228 1 93 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%RN 3 5 7 13 15 21
c40 21 0 7.48684e-20 $X=0.325 $Y=3.33
c41 3 0 1.63751e-20 $X=0.475 $Y=1.075
r42 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=3.33
+ $X2=0.325 $Y2=3.33
r43 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=2.305
+ $X2=0.53 $Y2=2.305
r44 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r45 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.47
+ $X2=0.32 $Y2=2.305
r46 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=2.47 $X2=0.32
+ $Y2=3.33
r47 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=2.305 $X2=0.53 $Y2=2.305
r48 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.53 $Y2=2.305
r49 5 7 1084.5 $w=1.5e-07 $l=2.115e-06 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=4.585
r50 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.53 $Y2=2.305
r51 1 3 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_110_115# 1 3 10 13 15 17 18 20 23 26
+ 29 33 36 39 43 47 52 53 54 60 65 67 70 71 76
c207 71 0 1.63751e-20 $X=1.375 $Y=1.48
c208 60 0 7.48684e-20 $X=0.87 $Y=2.74
c209 53 0 1.90798e-19 $X=1.145 $Y=1.59
c210 39 0 1.09867e-19 $X=8.545 $Y=2.75
c211 26 0 1.70295e-19 $X=8.8 $Y=2.605
r212 71 73 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.375 $Y=1.48
+ $X2=1.23 $Y2=1.48
r213 70 76 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.715 $Y=1.48
+ $X2=8.86 $Y2=1.48
r214 70 71 7.06756 $w=1.7e-07 $l=7.34e-06 $layer=MET1_cond $X=8.715 $Y=1.48
+ $X2=1.375 $Y2=1.48
r215 67 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.86 $Y=1.48
+ $X2=8.86 $Y2=1.48
r216 67 69 5.02622 $w=2.67e-07 $l=1.1e-07 $layer=LI1_cond $X=8.86 $Y=1.48
+ $X2=8.86 $Y2=1.59
r217 63 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.48
+ $X2=1.23 $Y2=1.48
r218 63 65 6.15596 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=1.27 $Y=1.48
+ $X2=1.27 $Y2=1.59
r219 58 60 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.74
+ $X2=0.87 $Y2=2.74
r220 55 57 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.87 $Y2=1.59
r221 54 57 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.59
+ $X2=0.87 $Y2=1.59
r222 53 65 2.19618 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=1.27 $Y2=1.59
r223 53 54 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=0.955 $Y2=1.59
r224 52 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.655
+ $X2=0.87 $Y2=2.74
r225 51 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=1.59
r226 51 52 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=2.655
r227 47 49 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r228 45 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=2.74
r229 45 47 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=3.455
r230 41 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=1.59
r231 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=0.825
r232 39 40 60.25 $w=2.04e-07 $l=2.55e-07 $layer=POLY_cond $X=8.545 $Y=2.75
+ $X2=8.8 $Y2=2.75
r233 38 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.86
+ $Y=1.59 $X2=8.86 $Y2=1.59
r234 36 38 12.05 $w=2.4e-07 $l=6e-08 $layer=POLY_cond $X=8.8 $Y=1.59 $X2=8.86
+ $Y2=1.59
r235 32 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.59 $X2=1.23 $Y2=1.59
r236 32 33 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.23 $Y=1.59 $X2=1.29
+ $Y2=1.59
r237 27 29 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.29 $Y=2.82
+ $X2=1.425 $Y2=2.82
r238 26 40 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.8 $Y=2.605
+ $X2=8.8 $Y2=2.75
r239 25 36 13.7767 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=1.755
+ $X2=8.8 $Y2=1.59
r240 25 26 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=8.8 $Y=1.755
+ $X2=8.8 $Y2=2.605
r241 21 39 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.545 $Y=2.895
+ $X2=8.545 $Y2=2.75
r242 21 23 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=8.545 $Y=2.895
+ $X2=8.545 $Y2=4.585
r243 18 36 53.2208 $w=2.4e-07 $l=3.37565e-07 $layer=POLY_cond $X=8.535 $Y=1.425
+ $X2=8.8 $Y2=1.59
r244 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.535 $Y=1.425
+ $X2=8.535 $Y2=0.945
r245 15 33 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.435 $Y=1.425
+ $X2=1.29 $Y2=1.59
r246 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.435 $Y=1.425
+ $X2=1.435 $Y2=0.945
r247 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=2.895
+ $X2=1.425 $Y2=2.82
r248 11 13 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=1.425 $Y=2.895
+ $X2=1.425 $Y2=4.585
r249 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=2.745
+ $X2=1.29 $Y2=2.82
r250 9 33 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.755
+ $X2=1.29 $Y2=1.59
r251 9 10 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=1.29 $Y=1.755
+ $X2=1.29 $Y2=2.745
r252 3 49 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r253 3 47 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r254 1 43 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%SN 1 2 5 9 13 17 22 25 30 34 37 42 44
+ 45 50
c172 45 0 2.97185e-19 $X=1.855 $Y=2.96
r173 45 47 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=2.96
+ $X2=1.71 $Y2=2.96
r174 44 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.79 $Y=2.96
+ $X2=7.935 $Y2=2.96
r175 44 45 5.71471 $w=1.7e-07 $l=5.935e-06 $layer=MET1_cond $X=7.79 $Y=2.96
+ $X2=1.855 $Y2=2.96
r176 39 42 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=8.025 $Y2=2.295
r177 34 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.935 $Y=2.96
+ $X2=7.935 $Y2=2.96
r178 32 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=2.42
+ $X2=7.935 $Y2=2.295
r179 32 34 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.935 $Y=2.42
+ $X2=7.935 $Y2=2.96
r180 30 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=2.96
+ $X2=1.71 $Y2=2.96
r181 28 37 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.455
+ $X2=1.71 $Y2=2.37
r182 28 30 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.71 $Y=2.455
+ $X2=1.71 $Y2=2.96
r183 25 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.025
+ $Y=2.255 $X2=8.025 $Y2=2.255
r184 25 27 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=2.255
+ $X2=8.035 $Y2=2.42
r185 25 26 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=2.255
+ $X2=8.035 $Y2=2.09
r186 22 23 5.53115 $w=3.05e-07 $l=3.5e-08 $layer=POLY_cond $X=1.855 $Y=2.37
+ $X2=1.89 $Y2=2.37
r187 21 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=2.37 $X2=1.71 $Y2=2.37
r188 21 22 22.9148 $w=3.05e-07 $l=1.45e-07 $layer=POLY_cond $X=1.71 $Y=2.37
+ $X2=1.855 $Y2=2.37
r189 17 27 1110.14 $w=1.5e-07 $l=2.165e-06 $layer=POLY_cond $X=8.115 $Y=4.585
+ $X2=8.115 $Y2=2.42
r190 13 26 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=8.045 $Y=1.075
+ $X2=8.045 $Y2=2.09
r191 9 19 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=1.925 $Y=1.075
+ $X2=1.925 $Y2=1.775
r192 3 22 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=2.535
+ $X2=1.855 $Y2=2.37
r193 3 5 1051.17 $w=1.5e-07 $l=2.05e-06 $layer=POLY_cond $X=1.855 $Y=2.535
+ $X2=1.855 $Y2=4.585
r194 2 23 10.4756 $w=2.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=2.205
+ $X2=1.89 $Y2=2.37
r195 1 19 38.6248 $w=2.2e-07 $l=1.1e-07 $layer=POLY_cond $X=1.89 $Y=1.885
+ $X2=1.89 $Y2=1.775
r196 1 2 93.3405 $w=2.2e-07 $l=3.2e-07 $layer=POLY_cond $X=1.89 $Y=1.885
+ $X2=1.89 $Y2=2.205
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_432_520# 1 3 11 15 18 24 25 26 27 28
+ 30 33 37 42
c90 42 0 1.71621e-19 $X=3.887 $Y=1.415
c91 25 0 1.29912e-19 $X=3.71 $Y=1.765
c92 18 0 1.52962e-19 $X=2.295 $Y=2.765
c93 15 0 1.44224e-19 $X=2.285 $Y=4.585
c94 11 0 1.32807e-19 $X=2.285 $Y=1.075
r95 41 42 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.887 $Y=1.245
+ $X2=3.887 $Y2=1.415
r96 37 39 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=3.895 $Y=3.455
+ $X2=3.895 $Y2=5.835
r97 35 37 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=3.895 $Y=3.375
+ $X2=3.895 $Y2=3.455
r98 33 41 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=3.895 $Y=0.825
+ $X2=3.895 $Y2=1.245
r99 30 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.795 $Y=1.68
+ $X2=3.795 $Y2=1.415
r100 27 35 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=3.725 $Y=3.185
+ $X2=3.895 $Y2=3.375
r101 27 28 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=3.725 $Y=3.185
+ $X2=2.38 $Y2=3.185
r102 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=1.765
+ $X2=3.795 $Y2=1.68
r103 25 26 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.71 $Y=1.765
+ $X2=2.38 $Y2=1.765
r104 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=3.1
+ $X2=2.38 $Y2=3.185
r105 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.295 $Y=3.1
+ $X2=2.295 $Y2=2.765
r106 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=1.85
+ $X2=2.38 $Y2=1.765
r107 21 24 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.295 $Y=1.85
+ $X2=2.295 $Y2=2.765
r108 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=2.765 $X2=2.295 $Y2=2.765
r109 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.765
+ $X2=2.295 $Y2=2.93
r110 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.765
+ $X2=2.295 $Y2=2.6
r111 15 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.285 $Y=4.585
+ $X2=2.285 $Y2=2.93
r112 11 19 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=2.285 $Y=1.075
+ $X2=2.285 $Y2=2.6
r113 3 39 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=3.67
+ $Y=3.085 $X2=3.895 $Y2=5.835
r114 3 37 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=3.67
+ $Y=3.085 $X2=3.895 $Y2=3.455
r115 1 33 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=3.67
+ $Y=0.575 $X2=3.895 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%D 3 7 10 14 19
c39 19 0 1.41836e-19 $X=3.295 $Y=2.22
c40 10 0 1.12321e-19 $X=3.295 $Y=2.22
r41 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.295 $Y=2.22
+ $X2=3.295 $Y2=2.22
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=2.22 $X2=3.295 $Y2=2.22
r43 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=2.22
+ $X2=3.295 $Y2=2.385
r44 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=2.22
+ $X2=3.295 $Y2=2.055
r45 7 12 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=3.235 $Y=4.585
+ $X2=3.235 $Y2=2.385
r46 3 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.235 $Y=1.075
+ $X2=3.235 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c233 55 0 6.79641e-20 $X=5.49 $Y=2.59
c234 48 0 1.98654e-19 $X=4.135 $Y=1.85
c235 44 0 1.86602e-19 $X=4.05 $Y=2.59
c236 30 0 1.29912e-19 $X=4.135 $Y=1.685
c237 25 0 1.41836e-19 $X=3.655 $Y=2.765
r238 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.03 $Y=2.59
+ $X2=5.885 $Y2=2.59
r239 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.735 $Y=2.59
+ $X2=6.88 $Y2=2.59
r240 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.735 $Y=2.59
+ $X2=6.03 $Y2=2.59
r241 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.8 $Y=2.59
+ $X2=3.655 $Y2=2.59
r242 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.74 $Y=2.59
+ $X2=5.885 $Y2=2.59
r243 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.74 $Y=2.59
+ $X2=3.8 $Y2=2.59
r244 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=2.59
+ $X2=5.885 $Y2=2.59
r245 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.885 $Y=2.59
+ $X2=5.885 $Y2=2.765
r246 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.655 $Y=2.59
+ $X2=3.655 $Y2=2.59
r247 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.655 $Y=2.59
+ $X2=3.655 $Y2=2.765
r248 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.88 $Y=2.59
+ $X2=6.88 $Y2=2.59
r249 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.88 $Y=2.59
+ $X2=6.88 $Y2=2.765
r250 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.59
+ $X2=5.885 $Y2=2.59
r251 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.8 $Y=2.59
+ $X2=5.49 $Y2=2.59
r252 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.405 $Y=2.505
+ $X2=5.49 $Y2=2.59
r253 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.405 $Y=2.505
+ $X2=5.405 $Y2=1.85
r254 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.135 $Y=2.505
+ $X2=4.135 $Y2=1.85
r255 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=2.59
+ $X2=3.655 $Y2=2.59
r256 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.05 $Y=2.59
+ $X2=4.135 $Y2=2.505
r257 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.05 $Y=2.59
+ $X2=3.74 $Y2=2.59
r258 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=2.765 $X2=6.88 $Y2=2.765
r259 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.762 $Y=1.685
+ $X2=6.762 $Y2=1.835
r260 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=2.765 $X2=5.885 $Y2=2.765
r261 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=2.765
+ $X2=5.885 $Y2=2.93
r262 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.85 $X2=5.405 $Y2=1.85
r263 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.85
+ $X2=5.405 $Y2=1.685
r264 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.85 $X2=4.135 $Y2=1.85
r265 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.85
+ $X2=4.135 $Y2=1.685
r266 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=2.765 $X2=3.655 $Y2=2.765
r267 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=2.765
+ $X2=3.655 $Y2=2.93
r268 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.79 $Y=2.6
+ $X2=6.837 $Y2=2.765
r269 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.79 $Y=2.6
+ $X2=6.79 $Y2=1.835
r270 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.735 $Y=2.93
+ $X2=6.837 $Y2=2.765
r271 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=6.735 $Y=2.93
+ $X2=6.735 $Y2=4.585
r272 17 40 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.735 $Y=1.075
+ $X2=6.735 $Y2=1.685
r273 13 39 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.945 $Y=4.585
+ $X2=5.945 $Y2=2.93
r274 10 34 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.345 $Y=1.075
+ $X2=5.345 $Y2=1.685
r275 7 30 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.195 $Y=1.075
+ $X2=4.195 $Y2=1.685
r276 3 27 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.595 $Y=4.585
+ $X2=3.595 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_217_617# 1 3 11 15 17 18 21 22 27 31
+ 35 39 40 43 49 54 55 56 61
c165 56 0 1.32807e-19 $X=1.855 $Y=1.85
c166 55 0 2.71143e-19 $X=4.49 $Y=1.85
c167 49 0 1.5821e-19 $X=4.725 $Y=2.765
c168 43 0 1.63226e-19 $X=1.71 $Y=0.825
c169 31 0 6.36774e-20 $X=4.985 $Y=4.585
c170 22 0 1.86602e-19 $X=4.63 $Y=2.765
c171 21 0 6.79641e-20 $X=4.91 $Y=2.765
c172 15 0 6.36774e-20 $X=4.555 $Y=4.585
r173 56 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.85
+ $X2=1.71 $Y2=1.85
r174 55 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.49 $Y=1.85
+ $X2=4.635 $Y2=1.85
r175 55 56 2.53719 $w=1.7e-07 $l=2.635e-06 $layer=MET1_cond $X=4.49 $Y=1.85
+ $X2=1.855 $Y2=1.85
r176 52 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.85
+ $X2=4.635 $Y2=1.85
r177 52 54 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=4.635 $Y=1.81
+ $X2=4.725 $Y2=1.81
r178 47 54 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.725 $Y=1.935
+ $X2=4.725 $Y2=1.81
r179 47 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.725 $Y=1.935
+ $X2=4.725 $Y2=2.765
r180 46 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.85
+ $X2=1.71 $Y2=1.85
r181 43 46 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=1.71 $Y=0.825
+ $X2=1.71 $Y2=1.85
r182 41 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.935
+ $X2=1.71 $Y2=1.85
r183 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=2.02
+ $X2=1.71 $Y2=1.935
r184 39 40 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.625 $Y=2.02
+ $X2=1.295 $Y2=2.02
r185 35 37 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.21 $Y=3.795
+ $X2=1.21 $Y2=5.835
r186 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.295 $Y2=2.02
r187 33 35 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.21 $Y2=3.795
r188 29 31 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.985 $Y=2.9
+ $X2=4.985 $Y2=4.585
r189 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.985 $Y=1.715
+ $X2=4.985 $Y2=1.075
r190 24 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=2.765 $X2=4.725 $Y2=2.765
r191 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=2.765
+ $X2=4.725 $Y2=2.765
r192 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=2.765
+ $X2=4.985 $Y2=2.9
r193 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=2.765
+ $X2=4.725 $Y2=2.765
r194 20 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=1.85 $X2=4.725 $Y2=1.85
r195 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=1.85
+ $X2=4.725 $Y2=1.85
r196 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=1.85
+ $X2=4.985 $Y2=1.715
r197 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=1.85
+ $X2=4.725 $Y2=1.85
r198 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.63 $Y2=2.765
r199 13 15 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.555 $Y2=4.585
r200 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.63 $Y2=1.85
r201 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.555 $Y2=1.075
r202 3 37 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=1.085 $Y=3.085 $X2=1.21 $Y2=5.835
r203 3 35 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=1.085 $Y=3.085 $X2=1.21 $Y2=3.795
r204 1 43 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.575 $X2=1.71 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_704_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c191 35 0 1.98654e-19 $X=3.715 $Y=1.76
c192 18 0 1.12321e-19 $X=4.195 $Y=4.585
r193 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=3.185
+ $X2=7.22 $Y2=3.185
r194 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=2.19
+ $X2=7.22 $Y2=2.19
r195 60 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=3.1
+ $X2=7.22 $Y2=3.185
r196 59 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.275
+ $X2=7.22 $Y2=2.19
r197 59 60 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=7.22 $Y=2.275
+ $X2=7.22 $Y2=3.1
r198 55 57 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.95 $Y=3.455
+ $X2=6.95 $Y2=5.835
r199 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=3.27
+ $X2=6.95 $Y2=3.185
r200 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.95 $Y=3.27
+ $X2=6.95 $Y2=3.455
r201 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=2.105
+ $X2=6.95 $Y2=2.19
r202 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.935
+ $X2=6.95 $Y2=1.85
r203 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.95 $Y=1.935
+ $X2=6.95 $Y2=2.105
r204 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.765
+ $X2=6.95 $Y2=1.85
r205 47 49 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.95 $Y=1.765
+ $X2=6.95 $Y2=0.825
r206 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=1.85
+ $X2=6.95 $Y2=1.85
r207 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.865 $Y=1.85
+ $X2=5.885 $Y2=1.85
r208 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=1.85 $X2=5.885 $Y2=1.85
r209 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.85
+ $X2=5.885 $Y2=2.015
r210 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.85
+ $X2=5.885 $Y2=1.685
r211 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.595 $Y=1.76
+ $X2=3.715 $Y2=1.76
r212 32 41 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.945 $Y=1.075
+ $X2=5.945 $Y2=1.685
r213 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.825 $Y=2.225
+ $X2=5.825 $Y2=2.015
r214 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=2.3
+ $X2=5.345 $Y2=2.3
r215 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.75 $Y=2.3
+ $X2=5.825 $Y2=2.225
r216 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.75 $Y=2.3
+ $X2=5.42 $Y2=2.3
r217 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.345 $Y=2.375
+ $X2=5.345 $Y2=2.3
r218 22 24 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=5.345 $Y=2.375
+ $X2=5.345 $Y2=4.585
r219 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=2.3
+ $X2=4.195 $Y2=2.3
r220 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=2.3
+ $X2=5.345 $Y2=2.3
r221 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.27 $Y=2.3 $X2=4.27
+ $Y2=2.3
r222 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=2.375
+ $X2=4.195 $Y2=2.3
r223 16 18 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=4.195 $Y=2.375
+ $X2=4.195 $Y2=4.585
r224 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=2.3
+ $X2=4.195 $Y2=2.3
r225 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.12 $Y=2.3
+ $X2=3.79 $Y2=2.3
r226 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=2.225
+ $X2=3.79 $Y2=2.3
r227 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.715 $Y=1.835
+ $X2=3.715 $Y2=1.76
r228 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.715 $Y=1.835
+ $X2=3.715 $Y2=2.225
r229 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.685
+ $X2=3.595 $Y2=1.76
r230 9 11 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.595 $Y=1.685
+ $X2=3.595 $Y2=1.075
r231 3 57 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.81
+ $Y=3.085 $X2=6.95 $Y2=5.835
r232 3 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.81
+ $Y=3.085 $X2=6.95 $Y2=3.455
r233 1 49 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.81
+ $Y=0.575 $X2=6.95 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_1246_89# 1 3 11 15 23 26 28 32 33 35
+ 36 37 38 40 46 50 54 56 61 62 67
c173 46 0 1.63226e-19 $X=8.26 $Y=0.825
c174 37 0 8.77106e-20 $X=9.47 $Y=2.855
c175 32 0 2.20654e-19 $X=9.38 $Y=2.19
r176 62 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.51 $Y=2.19
+ $X2=6.365 $Y2=2.19
r177 61 67 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.235 $Y=2.19
+ $X2=9.38 $Y2=2.19
r178 61 62 2.62385 $w=1.7e-07 $l=2.725e-06 $layer=MET1_cond $X=9.235 $Y=2.19
+ $X2=6.51 $Y2=2.19
r179 56 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.38 $Y=2.19
+ $X2=9.38 $Y2=2.19
r180 54 56 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.845 $Y=2.19
+ $X2=9.38 $Y2=2.19
r181 50 52 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=8.76 $Y=3.795
+ $X2=8.76 $Y2=5.835
r182 48 54 5.37722 $w=2.41e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=2.275
+ $X2=8.845 $Y2=2.19
r183 48 50 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=8.76 $Y=2.275
+ $X2=8.76 $Y2=3.795
r184 44 48 25.3112 $w=2.41e-07 $l=6.89202e-07 $layer=LI1_cond $X=8.26 $Y=1.825
+ $X2=8.76 $Y2=2.275
r185 44 46 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=8.26 $Y=1.825
+ $X2=8.26 $Y2=0.825
r186 40 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.365 $Y=2.19
+ $X2=6.365 $Y2=2.19
r187 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=2.855
+ $X2=9.47 $Y2=3.005
r188 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=1.65 $X2=9.47
+ $Y2=1.8
r189 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.445 $Y=2.355
+ $X2=9.445 $Y2=2.855
r190 33 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.445 $Y=2.025
+ $X2=9.445 $Y2=1.8
r191 32 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.38
+ $Y=2.19 $X2=9.38 $Y2=2.19
r192 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=2.19
+ $X2=9.382 $Y2=2.355
r193 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=2.19
+ $X2=9.382 $Y2=2.025
r194 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=2.19 $X2=6.365 $Y2=2.19
r195 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=2.19
+ $X2=6.365 $Y2=2.355
r196 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=2.19
+ $X2=6.365 $Y2=2.025
r197 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=9.495 $Y=4.585
+ $X2=9.495 $Y2=3.005
r198 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.495 $Y=1.075
+ $X2=9.495 $Y2=1.65
r199 15 30 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=6.305 $Y=4.585
+ $X2=6.305 $Y2=2.355
r200 11 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.305 $Y=1.075
+ $X2=6.305 $Y2=2.025
r201 3 52 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=8.62
+ $Y=3.085 $X2=8.76 $Y2=5.835
r202 3 50 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=8.62
+ $Y=3.085 $X2=8.76 $Y2=3.795
r203 1 46 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=8.12
+ $Y=0.575 $X2=8.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_1084_115# 1 3 10 11 13 16 20 26 31 32
+ 33 34 35 38 42 47 52 53 58
c157 53 0 1.5821e-19 $X=5.21 $Y=1.85
c158 32 0 1.67294e-19 $X=5.475 $Y=1.43
c159 31 0 1.57671e-19 $X=5.065 $Y=1.85
c160 16 0 6.36774e-20 $X=7.685 $Y=4.585
r161 53 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.21 $Y=1.85
+ $X2=5.065 $Y2=1.85
r162 52 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=1.85
+ $X2=7.595 $Y2=1.85
r163 52 53 2.15686 $w=1.7e-07 $l=2.24e-06 $layer=MET1_cond $X=7.45 $Y=1.85
+ $X2=5.21 $Y2=1.85
r164 47 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=1.85
+ $X2=7.595 $Y2=1.85
r165 47 50 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.595 $Y=1.85
+ $X2=7.595 $Y2=2.765
r166 42 44 69.1466 $w=3.38e-07 $l=2.04e-06 $layer=LI1_cond $X=5.645 $Y=3.795
+ $X2=5.645 $Y2=5.835
r167 40 42 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=5.645 $Y=3.27
+ $X2=5.645 $Y2=3.795
r168 36 38 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=5.645 $Y=1.345
+ $X2=5.645 $Y2=0.825
r169 34 40 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=3.185
+ $X2=5.645 $Y2=3.27
r170 34 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=3.185
+ $X2=5.15 $Y2=3.185
r171 32 36 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=1.43
+ $X2=5.645 $Y2=1.345
r172 32 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=1.43
+ $X2=5.15 $Y2=1.43
r173 31 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.065 $Y=1.85
+ $X2=5.065 $Y2=1.85
r174 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=3.1
+ $X2=5.15 $Y2=3.185
r175 29 31 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.065 $Y=3.1
+ $X2=5.065 $Y2=1.85
r176 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=1.515
+ $X2=5.15 $Y2=1.43
r177 28 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.065 $Y=1.515
+ $X2=5.065 $Y2=1.85
r178 25 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=2.765 $X2=7.595 $Y2=2.765
r179 25 26 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=2.765
+ $X2=7.685 $Y2=2.765
r180 22 25 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=2.765
+ $X2=7.595 $Y2=2.765
r181 18 20 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=7.505 $Y=1.77
+ $X2=7.685 $Y2=1.77
r182 14 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.685 $Y=2.9
+ $X2=7.685 $Y2=2.765
r183 14 16 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=7.685 $Y=2.9
+ $X2=7.685 $Y2=4.585
r184 11 20 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.685 $Y=1.69
+ $X2=7.685 $Y2=1.77
r185 11 13 197.62 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=7.685 $Y=1.69
+ $X2=7.685 $Y2=1.075
r186 10 22 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.505 $Y=2.63
+ $X2=7.505 $Y2=2.765
r187 9 18 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.505 $Y=1.85
+ $X2=7.505 $Y2=1.77
r188 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.505 $Y=1.85
+ $X2=7.505 $Y2=2.63
r189 3 44 171.429 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=3 $X=5.42
+ $Y=3.085 $X2=5.645 $Y2=5.835
r190 3 42 171.429 $w=1.7e-07 $l=8.1477e-07 $layer=licon1_PDIFF $count=3 $X=5.42
+ $Y=3.085 $X2=5.645 $Y2=3.795
r191 1 38 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=5.42
+ $Y=0.575 $X2=5.645 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c81 44 0 8.77106e-20 $X=9.285 $Y=2.96
c82 35 0 9.99996e-20 $X=9.78 $Y=2.765
c83 33 0 1.20654e-19 $X=9.78 $Y=1.85
c84 27 0 1.09867e-19 $X=9.28 $Y=2.96
c85 23 0 1.70295e-19 $X=9.28 $Y=0.825
c86 18 0 1.98165e-19 $X=9.865 $Y=2.395
r87 42 44 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=9.28 $Y=2.96
+ $X2=9.285 $Y2=2.96
r88 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.865 $Y=2.68
+ $X2=9.865 $Y2=2.395
r89 37 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.865 $Y=1.935
+ $X2=9.865 $Y2=2.395
r90 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=2.765
+ $X2=9.865 $Y2=2.68
r91 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=2.765
+ $X2=9.365 $Y2=2.765
r92 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.85
+ $X2=9.865 $Y2=1.935
r93 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=1.85
+ $X2=9.365 $Y2=1.85
r94 29 31 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=9.28 $Y=3.455
+ $X2=9.28 $Y2=5.835
r95 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=2.96
+ $X2=9.28 $Y2=2.96
r96 27 29 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.28 $Y=2.96
+ $X2=9.28 $Y2=3.455
r97 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=2.85
+ $X2=9.365 $Y2=2.765
r98 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.28 $Y=2.85
+ $X2=9.28 $Y2=2.96
r99 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=1.765
+ $X2=9.365 $Y2=1.85
r100 21 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.28 $Y=1.765
+ $X2=9.28 $Y2=0.825
r101 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.865
+ $Y=2.395 $X2=9.865 $Y2=2.395
r102 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=2.395
+ $X2=9.865 $Y2=2.56
r103 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=2.395
+ $X2=9.865 $Y2=2.23
r104 15 20 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=9.925 $Y=4.585
+ $X2=9.925 $Y2=2.56
r105 11 19 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.925 $Y=1.075
+ $X2=9.925 $Y2=2.23
r106 3 31 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=9.155
+ $Y=3.085 $X2=9.28 $Y2=5.835
r107 3 29 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=9.155
+ $Y=3.085 $X2=9.28 $Y2=3.455
r108 1 23 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=9.155
+ $Y=0.575 $X2=9.28 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_300_617# 1 2 11 15 16 19
r20 19 21 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.5 $Y=3.795
+ $X2=2.5 $Y2=5.835
r21 17 19 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.5 $Y=3.715 $X2=2.5
+ $Y2=3.795
r22 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=3.63
+ $X2=2.5 $Y2=3.715
r23 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.415 $Y=3.63
+ $X2=1.725 $Y2=3.63
r24 11 13 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.64 $Y=3.795
+ $X2=1.64 $Y2=5.835
r25 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.715
+ $X2=1.725 $Y2=3.63
r26 9 11 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.64 $Y=3.715 $X2=1.64
+ $Y2=3.795
r27 2 21 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.36
+ $Y=3.085 $X2=2.5 $Y2=5.835
r28 2 19 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=2.36
+ $Y=3.085 $X2=2.5 $Y2=3.795
r29 1 13 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=5.835
r30 1 11 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=3.085 $X2=1.64 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%A_1469_617# 1 2 11 15 16 19
r19 19 21 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=8.33 $Y=3.795
+ $X2=8.33 $Y2=5.835
r20 17 19 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=8.33 $Y=3.715 $X2=8.33
+ $Y2=3.795
r21 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.245 $Y=3.63
+ $X2=8.33 $Y2=3.715
r22 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.245 $Y=3.63
+ $X2=7.555 $Y2=3.63
r23 11 13 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=7.47 $Y=3.795
+ $X2=7.47 $Y2=5.835
r24 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=3.715
+ $X2=7.555 $Y2=3.63
r25 9 11 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.47 $Y=3.715 $X2=7.47
+ $Y2=3.795
r26 2 21 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=8.19
+ $Y=3.085 $X2=8.33 $Y2=5.835
r27 2 19 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=8.19
+ $Y=3.085 $X2=8.33 $Y2=3.795
r28 1 13 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=7.345
+ $Y=3.085 $X2=7.47 $Y2=5.835
r29 1 11 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=7.345
+ $Y=3.085 $X2=7.47 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFSR_1%Q 1 3 11 15 22 25 29 32
r20 27 29 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=3.09
+ $X2=10.255 $Y2=3.09
r21 23 25 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=1.515
+ $X2=10.255 $Y2=1.515
r22 22 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=3.005
+ $X2=10.255 $Y2=3.09
r23 21 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=1.6
+ $X2=10.255 $Y2=1.515
r24 21 22 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=10.255 $Y=1.6
+ $X2=10.255 $Y2=3.005
r25 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=10.14 $Y=3.455
+ $X2=10.14 $Y2=5.835
r26 15 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.14 $Y=3.33
+ $X2=10.14 $Y2=3.33
r27 15 17 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.14 $Y2=3.455
r28 13 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=3.175
+ $X2=10.14 $Y2=3.09
r29 13 15 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.14 $Y=3.175
+ $X2=10.14 $Y2=3.33
r30 9 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=1.43
+ $X2=10.14 $Y2=1.515
r31 9 11 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=10.14 $Y=1.43
+ $X2=10.14 $Y2=0.825
r32 3 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=10
+ $Y=3.085 $X2=10.14 $Y2=5.835
r33 3 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=10
+ $Y=3.085 $X2=10.14 $Y2=3.455
r34 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=10 $Y=0.575
+ $X2=10.14 $Y2=0.825
.ends

