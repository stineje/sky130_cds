* File: sky130_osu_sc_12T_ls__tnbufi_l.pex.spice
* Created: Fri Nov 12 15:40:57 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_L%GND 1 17 19 26 35 38
r31 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r32 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r33 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r34 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r35 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r36 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r37 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r38 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r39 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_L%VDD 1 13 15 21 25 29 32
r17 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r18 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r19 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r20 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287 $X2=1.02
+ $Y2=4.287
r21 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r22 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.275
r23 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r24 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r25 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r26 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r27 1 21 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.025 $X2=0.69 $Y2=3.275
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_L%A_27_115# 1 3 11 16 20 24 26 28 30
c41 30 0 2.92524e-19 $X=0.69 $Y=2.06
r42 30 32 0.130481 $w=1.68e-07 $l=2e-09 $layer=LI1_cond $X=0.69 $Y=2.06 $X2=0.69
+ $Y2=2.062
r43 27 28 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.062
+ $X2=0.26 $Y2=2.062
r44 26 32 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=2.062
+ $X2=0.69 $Y2=2.062
r45 26 27 16.4779 $w=1.73e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=2.062
+ $X2=0.345 $Y2=2.062
r46 22 28 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.26 $Y=2.15 $X2=0.26
+ $Y2=2.062
r47 22 24 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=0.26 $Y=2.15
+ $X2=0.26 $Y2=3.275
r48 18 28 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=0.26 $Y=1.975
+ $X2=0.26 $Y2=2.062
r49 18 20 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=0.26 $Y=1.975
+ $X2=0.26 $Y2=0.74
r50 14 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.06 $X2=0.69 $Y2=2.06
r51 14 16 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=2.06
+ $X2=0.905 $Y2=2.06
r52 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.895
+ $X2=0.905 $Y2=2.06
r53 9 11 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=0.905 $Y=1.895
+ $X2=0.905 $Y2=0.755
r54 3 24 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.275
r55 1 20 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_L%OE 5 7 9 12 13 18 26
c42 7 0 1.78563e-19 $X=0.475 $Y=2.9
r43 24 26 0.00168464 $w=3.71e-07 $l=5e-09 $layer=MET1_cond $X=0.745 $Y=2.48
+ $X2=0.745 $Y2=2.485
r44 18 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r45 18 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.655
r46 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.655 $X2=0.69 $Y2=2.655
r47 13 14 66.3154 $w=1.49e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.61
+ $X2=0.475 $Y2=1.61
r48 7 16 49.2914 $w=4.58e-07 $l=4.23124e-07 $layer=POLY_cond $X=0.905 $Y=2.9
+ $X2=0.587 $Y2=2.655
r49 7 12 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.905 $Y=2.9
+ $X2=0.905 $Y2=3.445
r50 7 9 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=3.445
r51 3 14 2.66937 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.535
+ $X2=0.475 $Y2=1.61
r52 3 5 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.475 $Y=1.535
+ $X2=0.475 $Y2=0.755
r53 1 13 2.66937 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=1.685
+ $X2=0.27 $Y2=1.61
r54 1 7 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=0.27 $Y=1.685
+ $X2=0.27 $Y2=2.75
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_L%A 3 7 10 14 20
c36 7 0 1.13961e-19 $X=1.265 $Y=3.445
r37 18 20 0.00168464 $w=3.71e-07 $l=5e-09 $layer=MET1_cond $X=1.085 $Y=2.11
+ $X2=1.085 $Y2=2.115
r38 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=2.11
+ $X2=1.14 $Y2=2.11
r39 14 16 10.2591 $w=2.2e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=2.045
+ $X2=1.325 $Y2=2.045
r40 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.98 $X2=1.325 $Y2=1.98
r41 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.98
+ $X2=1.325 $Y2=2.145
r42 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.98
+ $X2=1.325 $Y2=1.815
r43 7 12 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=1.265 $Y=3.445
+ $X2=1.265 $Y2=2.145
r44 3 11 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.265 $Y=0.755
+ $X2=1.265 $Y2=1.815
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_L%Y 1 3 10 16 24 27 31
r31 31 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.37
+ $X2=1.48 $Y2=1.485
r32 27 28 0.0806629 $w=2.95e-07 $l=1.15e-07 $layer=MET1_cond $X=1.477 $Y=2.85
+ $X2=1.477 $Y2=2.735
r33 24 28 0.986954 $w=1.7e-07 $l=1.025e-06 $layer=MET1_cond $X=1.51 $Y=1.71
+ $X2=1.51 $Y2=2.735
r34 24 33 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.51 $Y=1.71
+ $X2=1.51 $Y2=1.485
r35 16 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.85
+ $X2=1.48 $Y2=2.85
r36 16 19 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.48 $Y=2.85
+ $X2=1.48 $Y2=3.275
r37 13 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.37
+ $X2=1.48 $Y2=1.37
r38 10 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.48 $Y=0.74
+ $X2=1.48 $Y2=1.37
r39 3 19 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=3.025 $X2=1.48 $Y2=3.275
r40 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.74
.ends

