* File: sky130_osu_sc_12T_ls__buf_4.spice
* Created: Fri Nov 12 15:35:14 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__buf_4.pex.spice"
.subckt sky130_osu_sc_12T_ls__buf_4  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1005 N_GND_M1005_d N_A_M1005_g N_A_27_115#_M1005_s N_GND_M1005_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1005_d N_GND_M1005_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001.5 A=0.078 P=1.34 MULT=1
MM1001 N_Y_M1000_d N_A_27_115#_M1001_g N_GND_M1001_s N_GND_M1005_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1007 N_Y_M1007_d N_A_27_115#_M1007_g N_GND_M1001_s N_GND_M1005_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.5
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1008 N_Y_M1007_d N_A_27_115#_M1008_g N_GND_M1008_s N_GND_M1005_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.9
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g N_A_27_115#_M1003_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A_27_115#_M1002_g N_VDD_M1003_d N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1002_d N_A_27_115#_M1004_g N_VDD_M1004_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A_27_115#_M1006_g N_VDD_M1004_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1006_d N_A_27_115#_M1009_g N_VDD_M1009_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref N_GND_M1005_b N_VDD_M1003_b NWDIODE A=5.7783 P=9.73
pX11_noxref noxref_6 A A PROBETYPE=1
pX12_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__buf_4.pxi.spice"
*
.ends
*
*
