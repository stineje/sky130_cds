* File: sky130_osu_sc_18T_hs__tnbufi_1.pxi.spice
* Created: Fri Nov 12 13:53:50 2021
* 
x_PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%GND N_GND_M1003_d N_GND_M1003_b N_GND_c_7_p
+ N_GND_c_2_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%GND
x_PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%VDD N_VDD_M1002_d N_VDD_M1002_b N_VDD_c_36_p
+ N_VDD_c_40_p N_VDD_c_41_p VDD N_VDD_c_37_p
+ PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%VDD
x_PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1002_s N_A_27_115#_M1001_g N_A_27_115#_c_57_n N_A_27_115#_c_59_n
+ N_A_27_115#_c_62_n N_A_27_115#_c_63_n N_A_27_115#_c_64_n N_A_27_115#_c_65_n
+ PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%OE N_OE_c_98_n N_OE_M1003_g N_OE_c_102_n
+ N_OE_M1002_g N_OE_M1000_g N_OE_c_103_n N_OE_c_104_n OE
+ PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%OE
x_PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%A N_A_M1005_g N_A_M1004_g N_A_c_143_n
+ N_A_c_144_n N_A_c_145_n A PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%A
x_PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%Y N_Y_M1005_d N_Y_M1004_d N_Y_c_189_n
+ N_Y_c_191_n Y N_Y_c_193_n N_Y_c_195_n PM_SKY130_OSU_SC_18T_HS__TNBUFI_1%Y
cc_1 N_GND_M1003_b N_A_27_115#_M1001_g 0.040426f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=1.075
cc_2 N_GND_c_2_p N_A_27_115#_M1001_g 0.00354579f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=1.075
cc_3 N_GND_c_3_p N_A_27_115#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=1.075
cc_4 N_GND_M1003_b N_A_27_115#_c_57_n 0.0434193f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=2.175
cc_5 N_GND_c_2_p N_A_27_115#_c_57_n 0.00105454f $X=0.69 $Y=0.825 $X2=0.905
+ $Y2=2.175
cc_6 N_GND_M1003_b N_A_27_115#_c_59_n 0.0198903f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_7 N_GND_c_7_p N_A_27_115#_c_59_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_8 N_GND_c_3_p N_A_27_115#_c_59_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_9 N_GND_M1003_b N_A_27_115#_c_62_n 0.0221237f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.455
cc_10 N_GND_M1003_b N_A_27_115#_c_63_n 0.00872418f $X=-0.045 $Y=0 $X2=0.605
+ $Y2=2.175
cc_11 N_GND_M1003_b N_A_27_115#_c_64_n 0.00647094f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.175
cc_12 N_GND_M1003_b N_A_27_115#_c_65_n 0.00382188f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=2.175
cc_13 N_GND_c_2_p N_A_27_115#_c_65_n 0.00516381f $X=0.69 $Y=0.825 $X2=0.69
+ $Y2=2.175
cc_14 N_GND_M1003_b N_OE_c_98_n 0.0186719f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.65
cc_15 N_GND_c_7_p N_OE_c_98_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.65
cc_16 N_GND_c_2_p N_OE_c_98_n 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.65
cc_17 N_GND_c_3_p N_OE_c_98_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.65
cc_18 N_GND_M1003_b N_OE_c_102_n 0.102331f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.01
cc_19 N_GND_M1003_b N_OE_c_103_n 0.0253119f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.725
cc_20 N_GND_M1003_b N_OE_c_104_n 0.00123196f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.765
cc_21 N_GND_M1003_b OE 5.10551e-19 $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_22 N_GND_M1003_b N_A_M1005_g 0.0430503f $X=-0.045 $Y=0 $X2=1.265 $Y2=1.075
cc_23 N_GND_c_3_p N_A_M1005_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.265 $Y2=1.075
cc_24 N_GND_M1003_b N_A_M1004_g 0.0426097f $X=-0.045 $Y=0 $X2=1.265 $Y2=4.585
cc_25 N_GND_M1003_b N_A_c_143_n 0.031953f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.09
cc_26 N_GND_M1003_b N_A_c_144_n 0.0125638f $X=-0.045 $Y=0 $X2=1.14 $Y2=3.33
cc_27 N_GND_M1003_b N_A_c_145_n 0.00872469f $X=-0.045 $Y=0 $X2=1.325 $Y2=2.09
cc_28 N_GND_M1003_b N_Y_c_189_n 0.00913846f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.825
cc_29 N_GND_c_3_p N_Y_c_189_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.48 $Y2=0.825
cc_30 N_GND_M1003_b N_Y_c_191_n 0.0151339f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.59
cc_31 N_GND_M1003_b Y 0.0395158f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.82
cc_32 N_GND_M1003_b N_Y_c_193_n 0.0122638f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.48
cc_33 N_GND_c_2_p N_Y_c_193_n 9.45275e-19 $X=0.69 $Y=0.825 $X2=1.48 $Y2=1.48
cc_34 N_GND_M1003_b N_Y_c_195_n 0.0157299f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.59
cc_35 N_VDD_M1002_b N_A_27_115#_c_62_n 0.0081036f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.455
cc_36 N_VDD_c_36_p N_A_27_115#_c_62_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=3.455
cc_37 N_VDD_c_37_p N_A_27_115#_c_62_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26
+ $Y2=3.455
cc_38 N_VDD_M1002_b N_OE_c_102_n 0.0554912f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=3.01
cc_39 N_VDD_c_36_p N_OE_c_102_n 0.00606474f $X=0.605 $Y=6.507 $X2=0.475 $Y2=3.01
cc_40 N_VDD_c_40_p N_OE_c_102_n 0.00772129f $X=0.69 $Y=3.795 $X2=0.475 $Y2=3.01
cc_41 N_VDD_c_41_p N_OE_c_102_n 0.00606474f $X=1.02 $Y=6.44 $X2=0.475 $Y2=3.01
cc_42 N_VDD_c_37_p N_OE_c_102_n 0.00937653f $X=1.02 $Y=6.47 $X2=0.475 $Y2=3.01
cc_43 N_VDD_M1002_b N_OE_c_104_n 0.0016861f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.765
cc_44 N_VDD_c_40_p N_OE_c_104_n 0.0038942f $X=0.69 $Y=3.795 $X2=0.69 $Y2=2.765
cc_45 N_VDD_M1002_b OE 0.00591461f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_46 N_VDD_c_40_p OE 0.00408652f $X=0.69 $Y=3.795 $X2=0.69 $Y2=2.96
cc_47 N_VDD_M1002_b N_A_M1004_g 0.0226933f $X=-0.045 $Y=2.905 $X2=1.265
+ $Y2=4.585
cc_48 N_VDD_c_41_p N_A_M1004_g 0.00606474f $X=1.02 $Y=6.44 $X2=1.265 $Y2=4.585
cc_49 N_VDD_c_37_p N_A_M1004_g 0.00468827f $X=1.02 $Y=6.47 $X2=1.265 $Y2=4.585
cc_50 N_VDD_M1002_b N_A_c_144_n 9.23313e-19 $X=-0.045 $Y=2.905 $X2=1.14 $Y2=3.33
cc_51 N_VDD_M1002_b N_Y_c_191_n 0.00976763f $X=-0.045 $Y=2.905 $X2=1.48 $Y2=2.59
cc_52 N_VDD_c_41_p N_Y_c_191_n 0.00757793f $X=1.02 $Y=6.44 $X2=1.48 $Y2=2.59
cc_53 N_VDD_c_37_p N_Y_c_191_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.48 $Y2=2.59
cc_54 N_A_27_115#_M1001_g N_OE_c_98_n 0.0267414f $X=0.905 $Y=1.075 $X2=0.475
+ $Y2=1.65
cc_55 N_A_27_115#_c_59_n N_OE_c_98_n 0.00804393f $X=0.26 $Y=0.825 $X2=0.475
+ $Y2=1.65
cc_56 N_A_27_115#_M1001_g N_OE_c_102_n 0.00301188f $X=0.905 $Y=1.075 $X2=0.475
+ $Y2=3.01
cc_57 N_A_27_115#_c_57_n N_OE_c_102_n 0.0400875f $X=0.905 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_58 N_A_27_115#_c_59_n N_OE_c_102_n 0.0121188f $X=0.26 $Y=0.825 $X2=0.475
+ $Y2=3.01
cc_59 N_A_27_115#_c_62_n N_OE_c_102_n 0.0486822f $X=0.26 $Y=3.455 $X2=0.475
+ $Y2=3.01
cc_60 N_A_27_115#_c_63_n N_OE_c_102_n 0.00111679f $X=0.605 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_61 N_A_27_115#_c_64_n N_OE_c_102_n 0.00632922f $X=0.26 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_62 N_A_27_115#_c_65_n N_OE_c_102_n 7.56328e-19 $X=0.69 $Y=2.175 $X2=0.475
+ $Y2=3.01
cc_63 N_A_27_115#_c_59_n N_OE_c_103_n 0.0104429f $X=0.26 $Y=0.825 $X2=0.475
+ $Y2=1.725
cc_64 N_A_27_115#_c_63_n N_OE_c_103_n 0.00711711f $X=0.605 $Y=2.175 $X2=0.475
+ $Y2=1.725
cc_65 N_A_27_115#_c_57_n N_OE_c_104_n 2.15234e-19 $X=0.905 $Y=2.175 $X2=0.69
+ $Y2=2.765
cc_66 N_A_27_115#_c_62_n N_OE_c_104_n 0.0193056f $X=0.26 $Y=3.455 $X2=0.69
+ $Y2=2.765
cc_67 N_A_27_115#_c_65_n N_OE_c_104_n 0.00847614f $X=0.69 $Y=2.175 $X2=0.69
+ $Y2=2.765
cc_68 N_A_27_115#_c_57_n OE 0.00125736f $X=0.905 $Y=2.175 $X2=0.69 $Y2=2.96
cc_69 N_A_27_115#_c_62_n OE 0.00651113f $X=0.26 $Y=3.455 $X2=0.69 $Y2=2.96
cc_70 N_A_27_115#_c_63_n OE 0.00158904f $X=0.605 $Y=2.175 $X2=0.69 $Y2=2.96
cc_71 N_A_27_115#_c_65_n OE 7.36678e-19 $X=0.69 $Y=2.175 $X2=0.69 $Y2=2.96
cc_72 N_A_27_115#_M1001_g N_A_M1005_g 0.0580253f $X=0.905 $Y=1.075 $X2=1.265
+ $Y2=1.075
cc_73 N_A_27_115#_c_57_n N_A_c_143_n 0.0580253f $X=0.905 $Y=2.175 $X2=1.325
+ $Y2=2.09
cc_74 N_A_27_115#_c_65_n N_A_c_143_n 2.55709e-19 $X=0.69 $Y=2.175 $X2=1.325
+ $Y2=2.09
cc_75 N_A_27_115#_c_57_n N_A_c_144_n 0.00134082f $X=0.905 $Y=2.175 $X2=1.14
+ $Y2=3.33
cc_76 N_A_27_115#_c_65_n N_A_c_144_n 0.00813625f $X=0.69 $Y=2.175 $X2=1.14
+ $Y2=3.33
cc_77 N_A_27_115#_M1001_g N_A_c_145_n 0.00160395f $X=0.905 $Y=1.075 $X2=1.325
+ $Y2=2.09
cc_78 N_A_27_115#_c_65_n N_A_c_145_n 0.00878007f $X=0.69 $Y=2.175 $X2=1.325
+ $Y2=2.09
cc_79 N_A_27_115#_c_62_n A 0.00539687f $X=0.26 $Y=3.455 $X2=1.14 $Y2=3.33
cc_80 N_A_27_115#_M1001_g Y 3.32545e-19 $X=0.905 $Y=1.075 $X2=1.525 $Y2=1.82
cc_81 N_A_27_115#_M1001_g N_Y_c_193_n 0.00101819f $X=0.905 $Y=1.075 $X2=1.48
+ $Y2=1.48
cc_82 N_OE_c_102_n N_A_M1004_g 0.206659f $X=0.475 $Y=3.01 $X2=1.265 $Y2=4.585
cc_83 N_OE_c_104_n N_A_M1004_g 4.61952e-19 $X=0.69 $Y=2.765 $X2=1.265 $Y2=4.585
cc_84 N_OE_c_102_n N_A_c_144_n 0.0110152f $X=0.475 $Y=3.01 $X2=1.14 $Y2=3.33
cc_85 N_OE_c_104_n N_A_c_144_n 0.0187675f $X=0.69 $Y=2.765 $X2=1.14 $Y2=3.33
cc_86 OE N_A_c_144_n 0.007197f $X=0.69 $Y=2.96 $X2=1.14 $Y2=3.33
cc_87 N_OE_c_102_n A 0.0113129f $X=0.475 $Y=3.01 $X2=1.14 $Y2=3.33
cc_88 OE A 0.004991f $X=0.69 $Y=2.96 $X2=1.14 $Y2=3.33
cc_89 N_A_c_144_n A_196_617# 0.00616226f $X=1.14 $Y=3.33 $X2=0.98 $Y2=3.085
cc_90 A A_196_617# 0.0123769f $X=1.14 $Y=3.33 $X2=0.98 $Y2=3.085
cc_91 N_A_M1005_g N_Y_c_189_n 0.00587516f $X=1.265 $Y=1.075 $X2=1.48 $Y2=0.825
cc_92 N_A_c_143_n N_Y_c_189_n 8.70049e-19 $X=1.325 $Y=2.09 $X2=1.48 $Y2=0.825
cc_93 N_A_c_145_n N_Y_c_189_n 0.00216439f $X=1.325 $Y=2.09 $X2=1.48 $Y2=0.825
cc_94 N_A_M1004_g N_Y_c_191_n 0.0165057f $X=1.265 $Y=4.585 $X2=1.48 $Y2=2.59
cc_95 N_A_c_143_n N_Y_c_191_n 0.00102058f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_96 N_A_c_144_n N_Y_c_191_n 0.049778f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_97 N_A_c_145_n N_Y_c_191_n 0.00330615f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_98 A N_Y_c_191_n 0.00706656f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_99 N_A_M1005_g Y 0.00768908f $X=1.265 $Y=1.075 $X2=1.525 $Y2=1.82
cc_100 N_A_M1004_g Y 0.00511826f $X=1.265 $Y=4.585 $X2=1.525 $Y2=1.82
cc_101 N_A_c_143_n Y 0.00539093f $X=1.325 $Y=2.09 $X2=1.525 $Y2=1.82
cc_102 N_A_c_144_n Y 0.012418f $X=1.14 $Y=3.33 $X2=1.525 $Y2=1.82
cc_103 N_A_c_145_n Y 0.0130872f $X=1.325 $Y=2.09 $X2=1.525 $Y2=1.82
cc_104 N_A_M1005_g N_Y_c_193_n 0.00686905f $X=1.265 $Y=1.075 $X2=1.48 $Y2=1.48
cc_105 N_A_c_143_n N_Y_c_193_n 0.00129509f $X=1.325 $Y=2.09 $X2=1.48 $Y2=1.48
cc_106 N_A_c_145_n N_Y_c_193_n 0.00203451f $X=1.325 $Y=2.09 $X2=1.48 $Y2=1.48
cc_107 N_A_M1004_g N_Y_c_195_n 0.00489736f $X=1.265 $Y=4.585 $X2=1.48 $Y2=2.59
cc_108 N_A_c_143_n N_Y_c_195_n 0.00138163f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
cc_109 N_A_c_144_n N_Y_c_195_n 0.00656407f $X=1.14 $Y=3.33 $X2=1.48 $Y2=2.59
cc_110 N_A_c_145_n N_Y_c_195_n 0.00227834f $X=1.325 $Y=2.09 $X2=1.48 $Y2=2.59
