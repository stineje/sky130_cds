* File: sky130_osu_sc_12T_ms__dffr_1.pex.spice
* Created: Fri Nov 12 15:22:38 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%GND 1 2 3 4 5 6 7 8 9 121 125 127 134
+ 136 143 145 152 154 164 166 176 178 185 187 194 196 203 230 232
c245 194 0 5.73867e-20 $X=7.9 $Y=0.74
c246 176 0 1.71621e-19 $X=6.09 $Y=0.755
c247 152 0 3.07651e-19 $X=2.59 $Y=0.755
c248 134 0 5.44281e-20 $X=1.21 $Y=0.74
c249 121 0 1.61973e-19 $X=-0.05 $Y=0
r250 230 232 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.175 $Y2=0.152
r251 205 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.152
+ $X2=8.85 $Y2=0.152
r252 201 226 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.152
r253 201 203 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.74
r254 196 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.152
+ $X2=8.85 $Y2=0.152
r255 192 194 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.74
r256 188 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.152
+ $X2=7.04 $Y2=0.152
r257 183 222 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.152
r258 183 185 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.74
r259 179 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.152
+ $X2=6.09 $Y2=0.152
r260 178 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.152
+ $X2=7.04 $Y2=0.152
r261 174 221 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.152
r262 174 176 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.755
r263 166 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.152
+ $X2=6.09 $Y2=0.152
r264 162 164 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.34 $Y=0.305
+ $X2=4.34 $Y2=0.74
r265 155 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.152
+ $X2=2.59 $Y2=0.152
r266 150 217 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.152
r267 150 152 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.755
r268 146 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.152
+ $X2=2.07 $Y2=0.152
r269 145 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.152
+ $X2=2.59 $Y2=0.152
r270 141 216 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.152
r271 141 143 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.74
r272 137 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.152
+ $X2=1.21 $Y2=0.152
r273 136 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.152
+ $X2=2.07 $Y2=0.152
r274 132 215 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.152
r275 132 134 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.74
r276 127 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.152
+ $X2=1.21 $Y2=0.152
r277 123 125 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r278 121 232 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=0.19 $X2=9.175 $Y2=0.19
r279 121 230 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=0.19 $X2=0.335 $Y2=0.19
r280 121 192 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r281 121 187 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r282 121 197 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.985 $Y2=0.152
r283 121 162 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.34 $Y2=0.305
r284 121 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.255 $Y2=0.152
r285 121 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.425 $Y2=0.152
r286 121 123 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r287 121 128 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r288 121 205 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.935 $Y2=0.152
r289 121 196 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.765 $Y2=0.152
r290 121 197 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=7.985 $Y2=0.152
r291 121 187 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r292 121 188 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.125 $Y2=0.152
r293 121 178 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.955 $Y2=0.152
r294 121 179 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.175 $Y2=0.152
r295 121 166 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.005 $Y2=0.152
r296 121 167 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.425 $Y2=0.152
r297 121 154 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=4.255 $Y2=0.152
r298 121 155 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=2.675 $Y2=0.152
r299 121 145 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.505 $Y2=0.152
r300 121 146 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.155 $Y2=0.152
r301 121 136 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.985 $Y2=0.152
r302 121 137 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.295 $Y2=0.152
r303 121 127 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.125 $Y2=0.152
r304 121 128 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r305 9 203 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.575 $X2=8.85 $Y2=0.74
r306 8 194 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.74
r307 7 185 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.575 $X2=7.04 $Y2=0.74
r308 6 176 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.575 $X2=6.09 $Y2=0.755
r309 5 164 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.575 $X2=4.34 $Y2=0.74
r310 4 152 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.575 $X2=2.59 $Y2=0.755
r311 3 143 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.74
r312 2 134 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.74
r313 1 125 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%VDD 1 2 3 4 5 6 7 85 89 91 99 107 109
+ 117 119 127 129 137 139 145 149 164 168
c124 145 0 1.98165e-19 $X=8.85 $Y=3.265
r125 164 168 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=4.287
+ $X2=9.175 $Y2=4.287
r126 153 164 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=4.25 $X2=0.335 $Y2=4.25
r127 149 168 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=4.25 $X2=9.175 $Y2=4.25
r128 147 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=4.287
+ $X2=8.85 $Y2=4.287
r129 147 149 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=8.935 $Y=4.287
+ $X2=9.175 $Y2=4.287
r130 143 162 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.85 $Y=4.135
+ $X2=8.85 $Y2=4.287
r131 143 145 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.85 $Y=4.135
+ $X2=8.85 $Y2=3.265
r132 140 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=4.287
+ $X2=7.83 $Y2=4.287
r133 140 142 21.9153 $w=3.03e-07 $l=5.8e-07 $layer=LI1_cond $X=7.915 $Y=4.287
+ $X2=8.495 $Y2=4.287
r134 139 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=4.287
+ $X2=8.85 $Y2=4.287
r135 139 142 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.765 $Y=4.287
+ $X2=8.495 $Y2=4.287
r136 135 161 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.83 $Y=4.135
+ $X2=7.83 $Y2=4.287
r137 135 137 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=7.83 $Y=4.135
+ $X2=7.83 $Y2=3.275
r138 132 134 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.455 $Y=4.287
+ $X2=7.135 $Y2=4.287
r139 130 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.09 $Y2=4.287
r140 130 132 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.455 $Y2=4.287
r141 129 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=4.287
+ $X2=7.83 $Y2=4.287
r142 129 134 23.0489 $w=3.03e-07 $l=6.1e-07 $layer=LI1_cond $X=7.745 $Y=4.287
+ $X2=7.135 $Y2=4.287
r143 125 159 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=4.287
r144 125 127 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=3.21
r145 122 124 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=4.287
+ $X2=5.775 $Y2=4.287
r146 120 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=4.287
+ $X2=4.34 $Y2=4.287
r147 120 122 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.425 $Y=4.287
+ $X2=5.095 $Y2=4.287
r148 119 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=6.09 $Y2=4.287
r149 119 124 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=5.775 $Y2=4.287
r150 115 158 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.34 $Y=4.135
+ $X2=4.34 $Y2=4.287
r151 115 117 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.34 $Y=4.135
+ $X2=4.34 $Y2=3.295
r152 112 114 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=4.287
+ $X2=3.735 $Y2=4.287
r153 110 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=4.287
+ $X2=2.59 $Y2=4.287
r154 110 112 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.675 $Y=4.287
+ $X2=3.055 $Y2=4.287
r155 109 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=4.287
+ $X2=4.34 $Y2=4.287
r156 109 114 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=4.255 $Y=4.287
+ $X2=3.735 $Y2=4.287
r157 105 156 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.59 $Y=4.135
+ $X2=2.59 $Y2=4.287
r158 105 107 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.59 $Y=4.135
+ $X2=2.59 $Y2=3.295
r159 102 155 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=4.287
+ $X2=2 $Y2=4.287
r160 102 104 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=2.085 $Y=4.287
+ $X2=2.375 $Y2=4.287
r161 101 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=4.287
+ $X2=2.59 $Y2=4.287
r162 101 104 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=4.287
+ $X2=2.375 $Y2=4.287
r163 97 155 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2 $Y=4.135 $X2=2
+ $Y2=4.287
r164 97 99 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2 $Y=4.135 $X2=2
+ $Y2=3.275
r165 94 96 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=4.287
+ $X2=1.695 $Y2=4.287
r166 92 153 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r167 92 94 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.015 $Y2=4.287
r168 91 155 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=4.287
+ $X2=2 $Y2=4.287
r169 91 96 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.915 $Y=4.287
+ $X2=1.695 $Y2=4.287
r170 87 153 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r171 87 89 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r172 85 149 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=4.135 $X2=9.175 $Y2=4.22
r173 85 142 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=4.135 $X2=8.495 $Y2=4.22
r174 85 161 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=4.135 $X2=7.815 $Y2=4.22
r175 85 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=4.135 $X2=7.135 $Y2=4.22
r176 85 132 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=4.135 $X2=6.455 $Y2=4.22
r177 85 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=4.135 $X2=5.775 $Y2=4.22
r178 85 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=4.135 $X2=5.095 $Y2=4.22
r179 85 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=4.135 $X2=4.415 $Y2=4.22
r180 85 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=4.135 $X2=3.735 $Y2=4.22
r181 85 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=4.135 $X2=3.055 $Y2=4.22
r182 85 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=4.135 $X2=2.375 $Y2=4.22
r183 85 96 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=4.135 $X2=1.695 $Y2=4.22
r184 85 94 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=4.135 $X2=1.015 $Y2=4.22
r185 85 153 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=4.135 $X2=0.335 $Y2=4.22
r186 7 145 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=2.605 $X2=8.85 $Y2=3.265
r187 6 137 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=3.025 $X2=7.83 $Y2=3.275
r188 5 127 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=5.95
+ $Y=2.605 $X2=6.09 $Y2=3.21
r189 4 117 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=2.605 $X2=4.34 $Y2=3.295
r190 3 107 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.605 $X2=2.59 $Y2=3.295
r191 2 99 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=3.025 $X2=2 $Y2=3.275
r192 1 89 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%RN 3 5 7 13 15 21
c38 21 0 7.50258e-20 $X=0.325 $Y=2.85
r39 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=2.85
+ $X2=0.325 $Y2=2.85
r40 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.53 $Y2=1.825
r41 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r42 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=1.99
+ $X2=0.32 $Y2=1.825
r43 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=1.99 $X2=0.32
+ $Y2=2.85
r44 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.825 $X2=0.53 $Y2=1.825
r45 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.53 $Y2=1.825
r46 5 7 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=3.235
r47 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.53 $Y2=1.825
r48 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%A_110_115# 1 3 9 11 14 16 18 20 22 26 32
+ 36 41 42 43 46 51 55 59 60 61 63 65 68
c197 68 0 5.73867e-20 $X=7.89 $Y=1.37
c198 65 0 5.44281e-20 $X=1.22 $Y=1.37
c199 46 0 7.50258e-20 $X=0.87 $Y=2.26
c200 16 0 1.70108e-19 $X=7.615 $Y=1.52
r201 63 68 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=7.89 $Y=1.255
+ $X2=7.89 $Y2=1.37
r202 62 63 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=7.89 $Y=1.085
+ $X2=7.89 $Y2=1.255
r203 60 62 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=7.805 $Y=1
+ $X2=7.89 $Y2=1.085
r204 60 61 6.25874 $w=1.7e-07 $l=6.5e-06 $layer=MET1_cond $X=7.805 $Y=1
+ $X2=1.305 $Y2=1
r205 59 65 0.0829981 $w=2.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.22 $Y=1.255
+ $X2=1.22 $Y2=1.37
r206 58 61 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.22 $Y=1.085
+ $X2=1.305 $Y2=1
r207 58 59 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.22 $Y=1.085
+ $X2=1.22 $Y2=1.255
r208 57 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.89 $Y=1.37
+ $X2=7.89 $Y2=1.37
r209 55 57 7.74603 $w=2.52e-07 $l=1.6e-07 $layer=LI1_cond $X=7.89 $Y=1.21
+ $X2=7.89 $Y2=1.37
r210 53 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.22 $Y=1.37
+ $X2=1.22 $Y2=1.37
r211 51 53 9.25118 $w=2.11e-07 $l=1.6e-07 $layer=LI1_cond $X=1.26 $Y=1.21
+ $X2=1.26 $Y2=1.37
r212 48 49 10.0734 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.87 $Y2=1.16
r213 44 46 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.26
+ $X2=0.87 $Y2=2.26
r214 43 49 5.3812 $w=2.18e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.955 $Y=1.21
+ $X2=0.87 $Y2=1.16
r215 42 51 2.00497 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.135 $Y=1.21
+ $X2=1.26 $Y2=1.21
r216 42 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.135 $Y=1.21
+ $X2=0.955 $Y2=1.21
r217 41 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=2.26
r218 40 49 2.19618 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.16
r219 40 41 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=2.175
r220 36 38 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.95
+ $X2=0.69 $Y2=3.63
r221 34 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.26
r222 34 36 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.95
r223 30 48 2.19618 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=1.16
r224 30 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=0.755
r225 29 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.21 $X2=7.89 $Y2=1.21
r226 24 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.21 $X2=1.22 $Y2=1.21
r227 24 26 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.22 $Y=1.21
+ $X2=1.425 $Y2=1.21
r228 20 29 38.8445 $w=3.55e-07 $l=2.07918e-07 $layer=POLY_cond $X=7.685 $Y=1.045
+ $X2=7.782 $Y2=1.21
r229 20 22 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.685 $Y=1.045
+ $X2=7.685 $Y2=0.755
r230 16 29 58.5319 $w=3.55e-07 $l=3.84539e-07 $layer=POLY_cond $X=7.615 $Y=1.52
+ $X2=7.782 $Y2=1.21
r231 16 18 987.074 $w=1.5e-07 $l=1.925e-06 $layer=POLY_cond $X=7.615 $Y=1.52
+ $X2=7.615 $Y2=3.445
r232 12 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.375
+ $X2=1.425 $Y2=1.21
r233 12 14 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=1.425 $Y=1.375
+ $X2=1.425 $Y2=3.445
r234 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.045
+ $X2=1.425 $Y2=1.21
r235 9 11 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.425 $Y=1.045
+ $X2=1.425 $Y2=0.755
r236 3 38 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.63
r237 3 36 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.95
r238 1 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%A_342_442# 1 3 11 15 18 22 23 25 26 28
+ 31 36 38
c83 38 0 1.72079e-19 $X=3.365 $Y=0.755
c84 25 0 1.29912e-19 $X=3.28 $Y=1.285
r85 38 40 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=3.365 $Y=0.755
+ $X2=3.465 $Y2=0.755
r86 36 37 15.1353 $w=2.66e-07 $l=3.3e-07 $layer=LI1_cond $X=2.025 $Y=2.375
+ $X2=2.025 $Y2=2.705
r87 31 33 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=3.465 $Y=2.955
+ $X2=3.465 $Y2=3.635
r88 29 31 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=2.79
+ $X2=3.465 $Y2=2.955
r89 27 38 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.365 $Y=0.935
+ $X2=3.365 $Y2=0.755
r90 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=0.935
+ $X2=3.365 $Y2=1.2
r91 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=1.285
+ $X2=3.365 $Y2=1.2
r92 25 26 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.28 $Y=1.285
+ $X2=2.2 $Y2=1.285
r93 24 37 3.35683 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.195 $Y=2.705
+ $X2=2.025 $Y2=2.705
r94 23 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.295 $Y=2.705
+ $X2=3.465 $Y2=2.79
r95 23 24 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.295 $Y=2.705
+ $X2=2.195 $Y2=2.705
r96 22 36 9.15133 $w=2.66e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.11 $Y=2.21
+ $X2=2.025 $Y2=2.375
r97 21 26 6.81649 $w=1.7e-07 $l=2.25555e-07 $layer=LI1_cond $X=2.11 $Y=1.47
+ $X2=2.2 $Y2=1.285
r98 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.11 $Y=1.47
+ $X2=2.11 $Y2=2.21
r99 18 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.375 $X2=1.94 $Y2=2.375
r100 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.375
+ $X2=1.892 $Y2=2.54
r101 18 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.375
+ $X2=1.892 $Y2=2.21
r102 15 19 746.074 $w=1.5e-07 $l=1.455e-06 $layer=POLY_cond $X=1.855 $Y=0.755
+ $X2=1.855 $Y2=2.21
r103 11 20 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.785 $Y=3.445
+ $X2=1.785 $Y2=2.54
r104 3 33 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.605 $X2=3.465 $Y2=3.635
r105 3 31 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.605 $X2=3.465 $Y2=2.955
r106 1 40 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.575 $X2=3.465 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%D 3 7 10 14 19
c42 19 0 1.41836e-19 $X=2.865 $Y=1.74
c43 10 0 1.12321e-19 $X=2.865 $Y=1.74
r44 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.74
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.74 $X2=2.865 $Y2=1.74
r46 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.905
r47 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.575
r48 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=2.805 $Y=3.235
+ $X2=2.805 $Y2=1.905
r49 3 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.805 $Y=0.835
+ $X2=2.805 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%CK 3 7 10 13 15 17 18 20 23 25 29 30 33
+ 34 37 42 46 50 54 56 57 59 65 72 76 77 78 79 86
c251 76 0 1.89675e-19 $X=5.31 $Y=2.11
c252 59 0 3.12771e-20 $X=6.45 $Y=2.11
c253 57 0 6.79641e-20 $X=5.06 $Y=2.11
c254 56 0 1.70195e-19 $X=5.37 $Y=2.11
c255 50 0 1.98654e-19 $X=3.705 $Y=1.37
c256 46 0 1.86602e-19 $X=3.62 $Y=2.11
c257 37 0 4.72879e-20 $X=5.455 $Y=2.285
c258 30 0 1.29912e-19 $X=3.705 $Y=1.205
c259 25 0 1.41836e-19 $X=3.225 $Y=2.285
c260 18 0 1.37092e-19 $X=6.305 $Y=2.45
r261 79 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=2.11
+ $X2=5.455 $Y2=2.11
r262 78 86 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.305 $Y=2.11
+ $X2=6.45 $Y2=2.11
r263 78 79 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.305 $Y=2.11
+ $X2=5.6 $Y2=2.11
r264 77 81 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.37 $Y=2.11
+ $X2=3.225 $Y2=2.11
r265 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.31 $Y=2.11
+ $X2=5.455 $Y2=2.11
r266 76 77 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.31 $Y=2.11
+ $X2=3.37 $Y2=2.11
r267 72 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=2.11
+ $X2=5.455 $Y2=2.11
r268 72 74 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.455 $Y=2.11
+ $X2=5.455 $Y2=2.285
r269 65 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.225 $Y=2.11
+ $X2=3.225 $Y2=2.11
r270 65 68 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.225 $Y=2.11
+ $X2=3.225 $Y2=2.285
r271 59 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.45 $Y=2.11
+ $X2=6.45 $Y2=2.11
r272 59 62 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.45 $Y=2.11
+ $X2=6.45 $Y2=2.285
r273 56 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.11
+ $X2=5.455 $Y2=2.11
r274 56 57 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.37 $Y=2.11
+ $X2=5.06 $Y2=2.11
r275 52 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=2.025
+ $X2=5.06 $Y2=2.11
r276 52 54 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.975 $Y=2.025
+ $X2=4.975 $Y2=1.37
r277 48 50 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.705 $Y=2.025
+ $X2=3.705 $Y2=1.37
r278 47 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.11
+ $X2=3.225 $Y2=2.11
r279 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.11
+ $X2=3.705 $Y2=2.025
r280 46 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.62 $Y=2.11
+ $X2=3.31 $Y2=2.11
r281 45 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=2.285 $X2=6.45 $Y2=2.285
r282 40 42 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=6.305 $Y=1.28
+ $X2=6.385 $Y2=1.28
r283 37 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=2.285 $X2=5.455 $Y2=2.285
r284 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=2.285
+ $X2=5.455 $Y2=2.45
r285 33 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.37 $X2=4.975 $Y2=1.37
r286 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.37
+ $X2=4.975 $Y2=1.205
r287 29 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.37 $X2=3.705 $Y2=1.37
r288 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.37
+ $X2=3.705 $Y2=1.205
r289 25 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=2.285 $X2=3.225 $Y2=2.285
r290 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.285
+ $X2=3.225 $Y2=2.45
r291 23 45 38.571 $w=3.25e-07 $l=1.75656e-07 $layer=POLY_cond $X=6.385 $Y=2.12
+ $X2=6.407 $Y2=2.285
r292 22 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.385 $Y=1.355
+ $X2=6.385 $Y2=1.28
r293 22 23 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.385 $Y=1.355
+ $X2=6.385 $Y2=2.12
r294 18 45 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.305 $Y=2.45
+ $X2=6.407 $Y2=2.285
r295 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.305 $Y=2.45
+ $X2=6.305 $Y2=3.235
r296 15 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=1.28
r297 15 17 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=0.835
r298 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.515 $Y=3.235
+ $X2=5.515 $Y2=2.45
r299 10 34 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.915 $Y=0.835
+ $X2=4.915 $Y2=1.205
r300 7 30 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.765 $Y=0.835
+ $X2=3.765 $Y2=1.205
r301 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.165 $Y=3.235
+ $X2=3.165 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%A_217_605# 1 3 11 15 17 18 21 22 27 31
+ 35 37 38 41 47 52 53 58 60
c138 53 0 1.35571e-19 $X=4.06 $Y=1.37
c139 47 0 1.5821e-19 $X=4.295 $Y=2.285
c140 31 0 6.36774e-20 $X=4.555 $Y=3.235
c141 22 0 1.86602e-19 $X=4.2 $Y=2.285
c142 21 0 6.79641e-20 $X=4.48 $Y=2.285
c143 15 0 6.36774e-20 $X=4.125 $Y=3.235
r144 56 58 0.0982977 $w=2.45e-07 $l=1.4e-07 $layer=MET1_cond $X=1.64 $Y=1.372
+ $X2=1.78 $Y2=1.372
r145 53 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.37
+ $X2=4.205 $Y2=1.37
r146 53 58 2.19537 $w=1.7e-07 $l=2.28e-06 $layer=MET1_cond $X=4.06 $Y=1.37
+ $X2=1.78 $Y2=1.37
r147 50 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=1.37
+ $X2=4.205 $Y2=1.37
r148 50 52 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=1.33
+ $X2=4.295 $Y2=1.33
r149 45 52 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.295 $Y=1.455
+ $X2=4.295 $Y2=1.33
r150 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.295 $Y=1.455
+ $X2=4.295 $Y2=2.285
r151 44 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.37
+ $X2=1.64 $Y2=1.37
r152 41 44 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.64 $Y=0.74
+ $X2=1.64 $Y2=1.37
r153 39 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.64 $Y=1.725
+ $X2=1.64 $Y2=1.37
r154 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.64 $Y2=1.725
r155 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.295 $Y2=1.81
r156 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.895
+ $X2=1.295 $Y2=1.81
r157 33 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.21 $Y=1.895
+ $X2=1.21 $Y2=3.275
r158 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.555 $Y2=3.235
r159 25 27 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.555 $Y=1.235
+ $X2=4.555 $Y2=0.835
r160 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=2.285 $X2=4.295 $Y2=2.285
r161 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=2.285
+ $X2=4.295 $Y2=2.285
r162 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=2.285
+ $X2=4.555 $Y2=2.42
r163 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=2.285
+ $X2=4.295 $Y2=2.285
r164 20 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.37 $X2=4.295 $Y2=1.37
r165 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=1.37
+ $X2=4.295 $Y2=1.37
r166 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=1.37
+ $X2=4.555 $Y2=1.235
r167 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=1.37
+ $X2=4.295 $Y2=1.37
r168 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=2.42
+ $X2=4.2 $Y2=2.285
r169 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.125 $Y=2.42
+ $X2=4.125 $Y2=3.235
r170 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=1.235
+ $X2=4.2 $Y2=1.37
r171 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.125 $Y=1.235
+ $X2=4.125 $Y2=0.835
r172 3 35 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=3.025 $X2=1.21 $Y2=3.275
r173 1 41 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%A_618_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 51 55 60 63 67 69 70 75
c196 75 0 1.37092e-19 $X=6.36 $Y=1.74
c197 70 0 5.08695e-19 $X=5.6 $Y=1.74
c198 69 0 2.9867e-19 $X=6.215 $Y=1.74
c199 51 0 5.69161e-20 $X=6.52 $Y=0.755
c200 44 0 1.89675e-19 $X=5.455 $Y=1.725
c201 34 0 1.98654e-19 $X=3.285 $Y=1.28
c202 18 0 1.12321e-19 $X=3.765 $Y=3.235
r203 70 72 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=1.74
+ $X2=5.455 $Y2=1.74
r204 69 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.215 $Y=1.74
+ $X2=6.36 $Y2=1.74
r205 69 70 0.592173 $w=1.7e-07 $l=6.15e-07 $layer=MET1_cond $X=6.215 $Y=1.74
+ $X2=5.6 $Y2=1.74
r206 65 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=2.705
+ $X2=6.795 $Y2=2.705
r207 63 64 17.474 $w=1.92e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=1.725
+ $X2=6.795 $Y2=1.725
r208 62 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.36 $Y=1.74
+ $X2=6.36 $Y2=1.74
r209 62 63 10.1667 $w=1.92e-07 $l=1.6e-07 $layer=LI1_cond $X=6.36 $Y=1.725
+ $X2=6.52 $Y2=1.725
r210 60 67 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.62
+ $X2=6.795 $Y2=2.705
r211 59 64 1.10697 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=6.795 $Y=1.825
+ $X2=6.795 $Y2=1.725
r212 59 60 48.9848 $w=1.78e-07 $l=7.95e-07 $layer=LI1_cond $X=6.795 $Y=1.825
+ $X2=6.795 $Y2=2.62
r213 55 57 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.52 $Y=2.955
+ $X2=6.52 $Y2=3.635
r214 53 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.79
+ $X2=6.52 $Y2=2.705
r215 53 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=2.79
+ $X2=6.52 $Y2=2.955
r216 49 63 1.44825 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.52 $Y=1.625 $X2=6.52
+ $Y2=1.725
r217 49 51 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.52 $Y=1.625
+ $X2=6.52 $Y2=0.755
r218 47 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=1.74
+ $X2=5.455 $Y2=1.74
r219 44 47 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.455 $Y=1.725
+ $X2=5.455 $Y2=1.74
r220 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.725 $X2=5.455 $Y2=1.725
r221 39 41 18.9959 $w=3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.47 $Y=1.725
+ $X2=5.47 $Y2=1.82
r222 39 40 55.9777 $w=3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.47 $Y=1.725
+ $X2=5.47 $Y2=1.52
r223 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.165 $Y=1.28
+ $X2=3.285 $Y2=1.28
r224 30 40 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=5.515 $Y=0.835
+ $X2=5.515 $Y2=1.52
r225 27 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.99 $Y=1.82
+ $X2=4.915 $Y2=1.82
r226 26 41 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.32 $Y=1.82
+ $X2=5.47 $Y2=1.82
r227 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.32 $Y=1.82
+ $X2=4.99 $Y2=1.82
r228 22 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.915 $Y=1.895
+ $X2=4.915 $Y2=1.82
r229 22 24 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=4.915 $Y=1.895
+ $X2=4.915 $Y2=3.235
r230 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.82
+ $X2=3.765 $Y2=1.82
r231 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=1.82
+ $X2=4.915 $Y2=1.82
r232 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.84 $Y=1.82 $X2=3.84
+ $Y2=1.82
r233 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.895
+ $X2=3.765 $Y2=1.82
r234 16 18 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=3.765 $Y=1.895
+ $X2=3.765 $Y2=3.235
r235 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=1.82
+ $X2=3.765 $Y2=1.82
r236 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.69 $Y=1.82
+ $X2=3.36 $Y2=1.82
r237 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.285 $Y=1.745
+ $X2=3.36 $Y2=1.82
r238 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.355
+ $X2=3.285 $Y2=1.28
r239 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.285 $Y=1.355
+ $X2=3.285 $Y2=1.745
r240 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.205
+ $X2=3.165 $Y2=1.28
r241 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.165 $Y=1.205
+ $X2=3.165 $Y2=0.835
r242 3 57 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=3.635
r243 3 55 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=2.955
r244 1 51 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%A_1160_89# 1 3 11 14 26 29 30 31 32 33
+ 35 36 39 40 42 43 44 45 46 48 52 54 55 58 61 64 69 70 71 73 75 80 81
c211 44 0 8.77106e-20 $X=8.61 $Y=2.375
c212 39 0 2.20611e-19 $X=8.52 $Y=1.74
c213 36 0 1.31857e-19 $X=5.965 $Y=1.605
c214 35 0 2.19969e-19 $X=5.965 $Y=1.77
c215 33 0 1.50225e-19 $X=5.89 $Y=2.255
c216 31 0 2.82071e-19 $X=5.89 $Y=1.365
r217 80 81 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.52 $Y=1.74
+ $X2=8.375 $Y2=1.74
r218 75 81 1.32143 $w=1.75e-07 $l=1.46e-06 $layer=MET1_cond $X=6.915 $Y=1.737
+ $X2=8.375 $Y2=1.737
r219 72 75 0.0698591 $w=1.75e-07 $l=1.2657e-07 $layer=MET1_cond $X=6.825
+ $Y=1.825 $X2=6.915 $Y2=1.737
r220 72 73 0.501568 $w=1.8e-07 $l=5.7e-07 $layer=MET1_cond $X=6.825 $Y=1.825
+ $X2=6.825 $Y2=2.395
r221 71 77 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=2.48
+ $X2=5.935 $Y2=2.48
r222 70 73 0.0699153 $w=1.7e-07 $l=1.25499e-07 $layer=MET1_cond $X=6.735 $Y=2.48
+ $X2=6.825 $Y2=2.395
r223 70 71 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=6.735 $Y=2.48
+ $X2=6.08 $Y2=2.48
r224 64 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.52 $Y=1.74
+ $X2=8.52 $Y2=1.74
r225 62 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=1.74
+ $X2=7.47 $Y2=1.74
r226 62 64 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.555 $Y=1.74
+ $X2=8.52 $Y2=1.74
r227 60 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.825
+ $X2=7.47 $Y2=1.74
r228 60 61 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=7.47 $Y=1.825
+ $X2=7.47 $Y2=2.96
r229 56 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.655
+ $X2=7.47 $Y2=1.74
r230 56 58 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.47 $Y=1.655
+ $X2=7.47 $Y2=0.74
r231 54 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=3.045
+ $X2=7.47 $Y2=2.96
r232 54 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.385 $Y=3.045
+ $X2=7.125 $Y2=3.045
r233 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=3.13
+ $X2=7.125 $Y2=3.045
r234 50 52 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.04 $Y=3.13
+ $X2=7.04 $Y2=3.275
r235 48 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.935 $Y=2.48
+ $X2=5.935 $Y2=2.48
r236 46 68 17.1635 $w=1.82e-07 $l=2.62393e-07 $layer=LI1_cond $X=5.935 $Y=2.025
+ $X2=5.95 $Y2=1.77
r237 46 48 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.935 $Y=2.025
+ $X2=5.935 $Y2=2.48
r238 44 45 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=2.375
+ $X2=8.61 $Y2=2.525
r239 42 43 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=1.17 $X2=8.61
+ $Y2=1.32
r240 41 44 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=8.585 $Y=1.905
+ $X2=8.585 $Y2=2.375
r241 40 43 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.585 $Y=1.575
+ $X2=8.585 $Y2=1.32
r242 39 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.52
+ $Y=1.74 $X2=8.52 $Y2=1.74
r243 39 41 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.74
+ $X2=8.522 $Y2=1.905
r244 39 40 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.74
+ $X2=8.522 $Y2=1.575
r245 35 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.965
+ $Y=1.77 $X2=5.965 $Y2=1.77
r246 35 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=1.77
+ $X2=5.965 $Y2=1.935
r247 35 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=1.77
+ $X2=5.965 $Y2=1.605
r248 32 33 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.89 $Y=2.105
+ $X2=5.89 $Y2=2.255
r249 32 37 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.905 $Y=2.105
+ $X2=5.905 $Y2=1.935
r250 31 36 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.905 $Y=1.365
+ $X2=5.905 $Y2=1.605
r251 30 31 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=5.89 $Y=1.205
+ $X2=5.89 $Y2=1.365
r252 29 45 228.147 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=8.635 $Y=3.235
+ $X2=8.635 $Y2=2.525
r253 26 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.635 $Y=0.835
+ $X2=8.635 $Y2=1.17
r254 14 33 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=5.875 $Y=3.235
+ $X2=5.875 $Y2=2.255
r255 11 30 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.875 $Y=0.835
+ $X2=5.875 $Y2=1.205
r256 3 52 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=3.025 $X2=7.04 $Y2=3.275
r257 1 58 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.575 $X2=7.47 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%A_998_115# 1 3 11 15 18 23 25 26 29 33
+ 36 41 44 45 46 47 54
c143 47 0 2.65484e-19 $X=5.44 $Y=1.37
c144 46 0 3.12771e-20 $X=6.985 $Y=1.37
c145 45 0 1.5821e-19 $X=4.78 $Y=1.37
c146 41 0 1.71621e-19 $X=5.215 $Y=0.755
c147 36 0 1.70108e-19 $X=7.13 $Y=1.37
c148 33 0 9.35412e-20 $X=5.315 $Y=1.37
c149 23 0 1.57671e-19 $X=4.635 $Y=1.37
r150 47 52 0.0905432 $w=2.3e-07 $l=1.25e-07 $layer=MET1_cond $X=5.44 $Y=1.37
+ $X2=5.315 $Y2=1.37
r151 46 54 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=1.37
+ $X2=7.13 $Y2=1.37
r152 46 47 1.48765 $w=1.7e-07 $l=1.545e-06 $layer=MET1_cond $X=6.985 $Y=1.37
+ $X2=5.44 $Y2=1.37
r153 45 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.78 $Y=1.37
+ $X2=4.635 $Y2=1.37
r154 44 52 0.0969593 $w=2.3e-07 $l=1.35e-07 $layer=MET1_cond $X=5.18 $Y=1.37
+ $X2=5.315 $Y2=1.37
r155 44 45 0.385153 $w=1.7e-07 $l=4e-07 $layer=MET1_cond $X=5.18 $Y=1.37
+ $X2=4.78 $Y2=1.37
r156 41 43 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=5.222 $Y=0.755
+ $X2=5.222 $Y2=1.035
r157 36 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=1.37
+ $X2=7.13 $Y2=1.37
r158 33 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=1.37
+ $X2=5.315 $Y2=1.37
r159 33 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.315 $Y=1.37
+ $X2=5.315 $Y2=1.035
r160 27 29 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=5.215 $Y=2.79
+ $X2=5.215 $Y2=3.295
r161 25 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=2.705
+ $X2=5.215 $Y2=2.79
r162 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=2.705
+ $X2=4.72 $Y2=2.705
r163 23 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.37
+ $X2=4.635 $Y2=1.37
r164 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=2.62
+ $X2=4.72 $Y2=2.705
r165 21 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.635 $Y=2.62
+ $X2=4.635 $Y2=1.37
r166 18 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.37 $X2=7.13 $Y2=1.37
r167 18 20 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=7.162 $Y=1.37
+ $X2=7.162 $Y2=1.535
r168 18 19 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=7.162 $Y=1.37
+ $X2=7.162 $Y2=1.205
r169 15 20 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=7.255 $Y=3.445
+ $X2=7.255 $Y2=1.535
r170 11 19 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.255 $Y=0.755
+ $X2=7.255 $Y2=1.205
r171 3 29 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.605 $X2=5.215 $Y2=3.295
r172 1 41 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.575 $X2=5.215 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c86 42 0 8.77106e-20 $X=8.425 $Y=2.48
c87 33 0 1.02575e-19 $X=8.92 $Y=2.285
c88 31 0 1.18035e-19 $X=8.92 $Y=1.37
c89 18 0 1.98165e-19 $X=9.005 $Y=1.915
r90 40 42 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=8.42 $Y=2.48
+ $X2=8.425 $Y2=2.48
r91 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.005 $Y=2.2
+ $X2=9.005 $Y2=1.915
r92 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.005 $Y=1.455
+ $X2=9.005 $Y2=1.915
r93 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=2.285
+ $X2=9.005 $Y2=2.2
r94 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=2.285
+ $X2=8.505 $Y2=2.285
r95 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=1.37
+ $X2=9.005 $Y2=1.455
r96 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=1.37
+ $X2=8.505 $Y2=1.37
r97 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.48
r98 27 29 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=3.265
r99 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=2.37
+ $X2=8.505 $Y2=2.285
r100 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.42 $Y=2.37
+ $X2=8.42 $Y2=2.48
r101 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=1.285
+ $X2=8.505 $Y2=1.37
r102 21 23 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.42 $Y=1.285
+ $X2=8.42 $Y2=0.74
r103 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=1.915 $X2=9.005 $Y2=1.915
r104 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.915
+ $X2=9.005 $Y2=2.08
r105 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.915
+ $X2=9.005 $Y2=1.75
r106 15 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.065 $Y=3.235
+ $X2=9.065 $Y2=2.08
r107 11 19 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=9.065 $Y=0.835
+ $X2=9.065 $Y2=1.75
r108 3 29 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=2.605 $X2=8.42 $Y2=3.265
r109 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.575 $X2=8.42 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFR_1%Q 1 3 11 15 18 21 25 28
r20 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=2.807
+ $X2=9.395 $Y2=2.807
r21 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=2.85
+ $X2=9.275 $Y2=2.85
r22 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=9.275 $Y=2.807
+ $X2=9.28 $Y2=2.807
r23 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=1.035
+ $X2=9.395 $Y2=1.035
r24 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.395 $Y=2.68
+ $X2=9.395 $Y2=2.807
r25 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.12
+ $X2=9.395 $Y2=1.035
r26 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=9.395 $Y=1.12
+ $X2=9.395 $Y2=2.68
r27 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.28 $Y=2.935
+ $X2=9.28 $Y2=2.807
r28 13 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.28 $Y=2.935
+ $X2=9.28 $Y2=3.265
r29 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=0.95 $X2=9.28
+ $Y2=1.035
r30 9 11 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.28 $Y=0.95 $X2=9.28
+ $Y2=0.74
r31 3 15 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=2.605 $X2=9.28 $Y2=3.265
r32 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.575 $X2=9.28 $Y2=0.74
.ends

