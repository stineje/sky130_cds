* File: sky130_osu_sc_12T_ls__and2_8.spice
* Created: Fri Nov 12 15:34:11 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__and2_8.pex.spice"
.subckt sky130_osu_sc_12T_ls__and2_8  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1007 A_110_115# N_A_M1007_g N_A_27_115#_M1007_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75004.1 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1007_b NSHORT L=0.15 W=0.52
+ AD=0.091 AS=0.0546 PD=0.87 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75000.5
+ SB=75003.7 A=0.078 P=1.34 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1001_d N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.091 PD=0.8 PS=0.87 NRD=0 NRS=16.152 M=1 R=3.46667
+ SA=75001 SB=75003.2 A=0.078 P=1.34 MULT=1
MM1008 N_Y_M1000_d N_A_27_115#_M1008_g N_GND_M1008_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.5
+ SB=75002.8 A=0.078 P=1.34 MULT=1
MM1010 N_Y_M1010_d N_A_27_115#_M1010_g N_GND_M1008_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.9
+ SB=75002.3 A=0.078 P=1.34 MULT=1
MM1012 N_Y_M1010_d N_A_27_115#_M1012_g N_GND_M1012_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75002.3
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1014 N_Y_M1014_d N_A_27_115#_M1014_g N_GND_M1012_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75002.8
+ SB=75001.5 A=0.078 P=1.34 MULT=1
MM1015 N_Y_M1014_d N_A_27_115#_M1015_g N_GND_M1015_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75003.2
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1016 N_Y_M1016_d N_A_27_115#_M1016_g N_GND_M1015_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75003.6
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1019 N_Y_M1016_d N_A_27_115#_M1019_g N_GND_M1019_s N_GND_M1007_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75004.1
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1005 N_A_27_115#_M1005_d N_A_M1005_g N_VDD_M1005_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1017 N_VDD_M1017_d N_B_M1017_g N_A_27_115#_M1005_d N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75003.6 A=0.189 P=2.82 MULT=1
MM1002 N_VDD_M1017_d N_A_27_115#_M1002_g N_Y_M1002_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_27_115#_M1003_g N_Y_M1002_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1003_d N_A_27_115#_M1004_g N_Y_M1004_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_27_115#_M1006_g N_Y_M1004_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_VDD_M1006_d N_A_27_115#_M1009_g N_Y_M1009_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_VDD_M1011_d N_A_27_115#_M1011_g N_Y_M1009_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_VDD_M1011_d N_A_27_115#_M1013_g N_Y_M1013_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_VDD_M1018_d N_A_27_115#_M1018_g N_Y_M1013_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref N_GND_M1007_b N_VDD_M1005_b NWDIODE A=10.2897 P=14.11
pX21_noxref noxref_8 A A PROBETYPE=1
pX22_noxref noxref_9 B B PROBETYPE=1
pX23_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__and2_8.pxi.spice"
*
.ends
*
*
