* File: sky130_osu_sc_15T_hs__inv_4.spice
* Created: Fri Nov 12 14:30:59 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__inv_4.pex.spice"
.subckt sky130_osu_sc_15T_hs__inv_4  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_GND_M1002_d N_A_M1005_g N_Y_M1005_s N_GND_M1001_b NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_GND_M1007_d N_A_M1007_g N_Y_M1005_s N_GND_M1001_b NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001.5 A=0.3 P=4.3 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6 SB=75001
+ A=0.3 P=4.3 MULT=1
MM1004 N_VDD_M1003_d N_A_M1004_g N_Y_M1004_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001 SB=75000.6
+ A=0.3 P=4.3 MULT=1
MM1006 N_VDD_M1006_d N_A_M1006_g N_Y_M1004_s N_VDD_M1000_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001.5
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX8_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=6.962 P=10.62
pX9_noxref noxref_5 A A PROBETYPE=1
pX10_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__inv_4.pxi.spice"
*
.ends
*
*
