* File: sky130_osu_sc_12T_ms__oai21_l.pex.spice
* Created: Fri Nov 12 15:25:46 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%GND 1 17 19 26 35 38
r39 35 38 0.321969 $w=3e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.15 $X2=1.02
+ $Y2=0.15
r40 28 33 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.15 $X2=0.69
+ $Y2=0.15
r41 24 33 3.44808 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=0.3 $X2=0.69
+ $Y2=0.15
r42 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.3
+ $X2=0.69 $Y2=0.735
r43 19 33 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.15 $X2=0.69
+ $Y2=0.15
r44 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.185
+ $X2=1.02 $Y2=0.185
r45 17 28 9.96333 $w=3e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.15 $X2=0.775
+ $Y2=0.15
r46 17 19 10.1799 $w=2.98e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.15
+ $X2=0.605 $Y2=0.15
r47 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.57 $X2=0.69 $Y2=0.735
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%VDD 1 13 15 21 26 29 32
r25 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r26 26 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r27 19 26 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.05 $Y=4.135
+ $X2=1.05 $Y2=4.287
r28 19 21 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.05 $Y=4.135
+ $X2=1.05 $Y2=3.655
r29 15 26 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=4.287
+ $X2=1.05 $Y2=4.287
r30 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=4.287
+ $X2=0.34 $Y2=4.287
r31 13 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r32 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r33 1 21 600 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.605 $X2=1.05 $Y2=3.655
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%A0 3 5 8 12 15 16 19 25
r38 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.415 $Y=2.85
+ $X2=0.415 $Y2=2.85
r39 19 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.415 $Y=2.28
+ $X2=0.415 $Y2=2.85
r40 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=2.28 $X2=0.415 $Y2=2.28
r41 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.28
+ $X2=0.415 $Y2=2.445
r42 15 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.28
+ $X2=0.415 $Y2=2.115
r43 10 12 57.4094 $w=1.55e-07 $l=1.2e-07 $layer=POLY_cond $X=0.355 $Y=1.292
+ $X2=0.475 $Y2=1.292
r44 8 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=2.445
r45 3 12 3.61756 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=0.475 $Y=1.215
+ $X2=0.475 $Y2=1.292
r46 3 5 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=1.215
+ $X2=0.475 $Y2=0.83
r47 1 10 3.61756 $w=1.5e-07 $l=7.8e-08 $layer=POLY_cond $X=0.355 $Y=1.37
+ $X2=0.355 $Y2=1.292
r48 1 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.355 $Y=1.37
+ $X2=0.355 $Y2=2.115
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%A1 3 7 10 15 18 22
c57 15 0 1.60731e-19 $X=0.845 $Y=1.74
c58 7 0 1.14151e-19 $X=0.905 $Y=0.83
c59 3 0 3.26014e-20 $X=0.835 $Y=3.235
r60 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.895 $Y=2.48
+ $X2=0.895 $Y2=2.48
r61 18 19 5.0779 $w=2.18e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.48 $X2=0.87
+ $Y2=2.395
r62 15 19 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.845 $Y=1.74
+ $X2=0.845 $Y2=2.395
r63 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.74 $X2=0.845 $Y2=1.74
r64 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.845 $Y=1.74
+ $X2=0.845 $Y2=1.875
r65 10 11 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.845 $Y=1.74
+ $X2=0.845 $Y2=1.605
r66 7 11 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=0.905 $Y=0.83
+ $X2=0.905 $Y2=1.605
r67 3 12 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.835 $Y=3.235
+ $X2=0.835 $Y2=1.875
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%B0 1 3 7 13 15 17 20
c47 13 0 1.14151e-19 $X=1.2 $Y=2.11
r48 15 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.285 $Y=1.5
+ $X2=1.395 $Y2=1.5
r49 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.11 $X2=1.2
+ $Y2=2.11
r50 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=1.585
+ $X2=1.285 $Y2=1.5
r51 11 13 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.2 $Y=1.585
+ $X2=1.2 $Y2=2.11
r52 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.5 $X2=1.395 $Y2=1.5
r53 5 10 38.8629 $w=2.72e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.335 $Y=1.335
+ $X2=1.39 $Y2=1.5
r54 5 7 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.335 $Y=1.335
+ $X2=1.335 $Y2=0.83
r55 1 10 38.8629 $w=2.72e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.325 $Y=1.665
+ $X2=1.39 $Y2=1.5
r56 1 3 912.723 $w=1.5e-07 $l=1.78e-06 $layer=POLY_cond $X=1.325 $Y=1.665
+ $X2=1.325 $Y2=3.445
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%Y 1 3 4 15 17 18 21 25 28 37 38 43
c52 37 0 1.93333e-19 $X=1.54 $Y=2.48
r53 43 45 0.0917586 $w=2.9e-07 $l=1.2e-07 $layer=MET1_cond $X=1.55 $Y=1 $X2=1.55
+ $Y2=1.12
r54 38 45 1.40203 $w=1.5e-07 $l=1.245e-06 $layer=MET1_cond $X=1.56 $Y=2.365
+ $X2=1.56 $Y2=1.12
r55 37 38 0.0896135 $w=2.95e-07 $l=1.15e-07 $layer=MET1_cond $X=1.542 $Y=2.48
+ $X2=1.542 $Y2=2.365
r56 31 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r57 28 31 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.55 $Y=0.795
+ $X2=1.55 $Y2=1
r58 25 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.275
+ $X2=1.54 $Y2=3.19
r59 21 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.54 $Y=2.48
+ $X2=1.54 $Y2=2.48
r60 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.105
+ $X2=1.54 $Y2=3.19
r61 19 21 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.54 $Y=3.105
+ $X2=1.54 $Y2=2.48
r62 17 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=3.19
+ $X2=1.54 $Y2=3.19
r63 17 18 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.455 $Y=3.19
+ $X2=0.345 $Y2=3.19
r64 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.275
+ $X2=0.345 $Y2=3.19
r65 13 15 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.26 $Y=3.275
+ $X2=0.26 $Y2=3.63
r66 4 25 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=3.025 $X2=1.54 $Y2=3.275
r67 3 15 600 $w=1.7e-07 $l=1.0857e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.63
r68 1 28 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.57 $X2=1.55 $Y2=0.795
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OAI21_L%A_27_114# 1 2 11 13 14 17
r20 15 17 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.12 $Y=1.07 $X2=1.12
+ $Y2=0.75
r21 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.155
+ $X2=1.12 $Y2=1.07
r22 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.155
+ $X2=0.345 $Y2=1.155
r23 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.07
+ $X2=0.345 $Y2=1.155
r24 9 11 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.26 $Y=1.07 $X2=0.26
+ $Y2=0.75
r25 2 17 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.57
+ $X2=1.12 $Y2=0.75
r26 1 11 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.57 $X2=0.26 $Y2=0.75
.ends

