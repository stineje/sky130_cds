* File: sky130_osu_sc_15T_ls__xor2_l.pex.spice
* Created: Fri Nov 12 15:00:53 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%GND 1 2 33 35 43 45 55 67 69
r66 67 69 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r67 53 55 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.865
r68 46 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r69 41 59 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r70 41 43 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.865
r71 35 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r72 33 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r73 33 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r74 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r75 33 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r76 33 45 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r77 33 46 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r78 33 35 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r79 2 55 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.575 $X2=2.44 $Y2=0.865
r80 1 43 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%VDD 1 2 25 27 34 38 46 54 57 61
r45 57 61 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=2.38 $Y2=5.397
r46 54 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=5.36
+ $X2=2.38 $Y2=5.36
r47 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.44 $Y=3.885
+ $X2=2.44 $Y2=4.565
r48 44 54 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=5.245
+ $X2=2.44 $Y2=5.397
r49 44 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.44 $Y=5.245
+ $X2=2.44 $Y2=4.565
r50 41 43 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=5.397
+ $X2=1.7 $Y2=5.397
r51 39 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r52 39 41 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r53 38 54 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=5.397
+ $X2=2.44 $Y2=5.397
r54 38 43 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=5.397
+ $X2=1.7 $Y2=5.397
r55 34 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=3.885
+ $X2=0.69 $Y2=4.565
r56 32 52 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r57 32 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r58 29 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r59 27 52 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r60 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r61 25 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r62 25 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r63 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r64 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r65 2 49 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.825 $X2=2.44 $Y2=4.565
r66 2 46 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.825 $X2=2.44 $Y2=3.885
r67 1 37 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r68 1 34 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%A_27_115# 1 3 11 15 18 22 27 31 35 41 43
c76 41 0 6.74854e-20 $X=1.805 $Y=2.505
c77 35 0 1.52002e-20 $X=1.72 $Y=1.965
r78 39 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.805 $Y=2.05
+ $X2=1.805 $Y2=2.505
r79 36 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.965
+ $X2=0.26 $Y2=1.965
r80 36 38 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=1.965
+ $X2=0.845 $Y2=1.965
r81 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=1.965
+ $X2=1.805 $Y2=2.05
r82 35 38 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.72 $Y=1.965
+ $X2=0.845 $Y2=1.965
r83 31 33 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r84 29 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.05 $X2=0.26
+ $Y2=1.965
r85 29 31 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=0.26 $Y=2.05
+ $X2=0.26 $Y2=3.205
r86 25 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.88 $X2=0.26
+ $Y2=1.965
r87 25 27 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=0.26 $Y=1.88
+ $X2=0.26 $Y2=0.865
r88 22 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=2.505 $X2=1.805 $Y2=2.505
r89 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=2.505
+ $X2=1.805 $Y2=2.67
r90 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.965 $X2=0.845 $Y2=1.965
r91 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=1.965
+ $X2=0.845 $Y2=1.8
r92 15 24 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=1.865 $Y=3.825
+ $X2=1.865 $Y2=2.67
r93 11 19 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=1.8
r94 3 33 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r95 3 31 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r96 1 27 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%A 2 5 6 8 9 13 16 18 19 20 21 22 24 27
+ 28 34 37 40 45 50 52 53 58 61
c122 50 0 3.28297e-19 $X=2.235 $Y=1.96
r123 55 58 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=1.085 $Y=3.07
+ $X2=1.09 $Y2=3.07
r124 53 58 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=1.23 $Y=3.07
+ $X2=1.09 $Y2=3.07
r125 52 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2 $Y=3.07
+ $X2=2.145 $Y2=3.07
r126 52 53 0.741419 $w=1.7e-07 $l=7.7e-07 $layer=MET1_cond $X=2 $Y=3.07 $X2=1.23
+ $Y2=3.07
r127 47 50 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.145 $Y=1.96
+ $X2=2.235 $Y2=1.96
r128 45 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=3.07
+ $X2=1.085 $Y2=3.07
r129 42 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.845 $Y=3.07
+ $X2=1.085 $Y2=3.07
r130 37 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=3.07
+ $X2=2.145 $Y2=3.07
r131 35 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.045
+ $X2=2.145 $Y2=1.96
r132 35 37 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.145 $Y=2.045
+ $X2=2.145 $Y2=3.07
r133 34 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=2.985
+ $X2=0.845 $Y2=3.07
r134 33 40 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=2.59
+ $X2=0.845 $Y2=2.505
r135 33 34 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.845 $Y=2.59
+ $X2=0.845 $Y2=2.985
r136 31 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.96 $X2=2.235 $Y2=1.96
r137 28 31 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=1.825
+ $X2=2.235 $Y2=1.96
r138 26 27 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=2.675
+ $X2=0.845 $Y2=2.75
r139 24 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.505 $X2=0.845 $Y2=2.505
r140 24 26 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=0.845 $Y=2.505
+ $X2=0.845 $Y2=2.675
r141 20 21 41.4471 $w=2e-07 $l=1.25e-07 $layer=POLY_cond $X=0.45 $Y=1.39
+ $X2=0.45 $Y2=1.515
r142 18 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.1 $Y=1.825
+ $X2=2.235 $Y2=1.825
r143 18 19 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.1 $Y=1.825
+ $X2=1.94 $Y2=1.825
r144 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.865 $Y=1.75
+ $X2=1.94 $Y2=1.825
r145 14 16 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.865 $Y=1.75
+ $X2=1.865 $Y2=0.945
r146 13 27 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.75
r147 10 22 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=2.675
+ $X2=0.45 $Y2=2.675
r148 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=2.675
+ $X2=0.845 $Y2=2.675
r149 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=2.675
+ $X2=0.55 $Y2=2.675
r150 6 22 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.45 $Y2=2.675
r151 6 8 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=3.825
r152 5 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=1.39
r153 2 22 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=2.6
+ $X2=0.45 $Y2=2.675
r154 2 21 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=0.425 $Y=2.6
+ $X2=0.425 $Y2=1.515
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%A_238_89# 1 3 11 14 17 18 20 26 30 34
r64 30 32 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.87 $Y=3.205
+ $X2=2.87 $Y2=4.565
r65 28 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.675
+ $X2=2.87 $Y2=1.59
r66 28 30 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=2.87 $Y=1.675
+ $X2=2.87 $Y2=3.205
r67 24 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.505
+ $X2=2.87 $Y2=1.59
r68 24 26 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.87 $Y=1.505
+ $X2=2.87 $Y2=0.865
r69 20 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.59
+ $X2=2.87 $Y2=1.59
r70 20 22 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=1.59
+ $X2=1.325 $Y2=1.59
r71 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.59 $X2=1.325 $Y2=1.59
r72 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.59
+ $X2=1.325 $Y2=1.755
r73 17 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.59
+ $X2=1.325 $Y2=1.425
r74 14 19 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=1.265 $Y=3.825
+ $X2=1.265 $Y2=1.755
r75 11 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.265 $Y=0.945
+ $X2=1.265 $Y2=1.425
r76 3 32 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=2.825 $X2=2.87 $Y2=4.565
r77 3 30 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=2.825 $X2=2.87 $Y2=3.205
r78 1 26 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.575 $X2=2.87 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 20 21 23 29
c56 20 0 6.74854e-20 $X=2.655 $Y=2.545
c57 13 0 1.52002e-20 $X=2.655 $Y=2.34
c58 8 0 1.7901e-19 $X=2.3 $Y=1.465
c59 7 0 1.49287e-19 $X=2.58 $Y=1.465
r60 26 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.7 $X2=2.53
+ $Y2=2.7
r61 23 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.53 $Y=2.505
+ $X2=2.53 $Y2=2.7
r62 19 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=2.505 $X2=2.53 $Y2=2.505
r63 19 20 20.0833 $w=3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=2.545
+ $X2=2.655 $Y2=2.545
r64 14 20 18.9685 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.655 $Y=2.75
+ $X2=2.655 $Y2=2.545
r65 14 16 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.655 $Y=2.75
+ $X2=2.655 $Y2=3.825
r66 13 20 18.9685 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.655 $Y=2.34
+ $X2=2.655 $Y2=2.545
r67 12 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.54
+ $X2=2.655 $Y2=1.465
r68 12 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.655 $Y=1.54
+ $X2=2.655 $Y2=2.34
r69 9 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.39
+ $X2=2.655 $Y2=1.465
r70 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.655 $Y=1.39
+ $X2=2.655 $Y2=0.945
r71 7 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.465
+ $X2=2.655 $Y2=1.465
r72 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=1.465 $X2=2.3
+ $Y2=1.465
r73 4 19 49.0033 $w=3e-07 $l=3.94398e-07 $layer=POLY_cond $X=2.225 $Y=2.75
+ $X2=2.53 $Y2=2.545
r74 4 6 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.225 $Y=2.75
+ $X2=2.225 $Y2=3.825
r75 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=1.39
+ $X2=2.3 $Y2=1.465
r76 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.225 $Y=1.39
+ $X2=2.225 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__XOR2_L%Y 1 3 11 13 15 19 24 30 33 35
r58 35 37 0.0784753 $w=2.23e-07 $l=1.4e-07 $layer=MET1_cond $X=1.425 $Y=1.22
+ $X2=1.565 $Y2=1.22
r59 28 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=2.215
+ $X2=1.425 $Y2=2.33
r60 28 30 0.0433297 $w=1.7e-07 $l=4.5e-08 $layer=MET1_cond $X=1.425 $Y=2.215
+ $X2=1.425 $Y2=2.17
r61 27 35 0.0238602 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.335
+ $X2=1.425 $Y2=1.22
r62 27 30 0.804007 $w=1.7e-07 $l=8.35e-07 $layer=MET1_cond $X=1.425 $Y=1.335
+ $X2=1.425 $Y2=2.17
r63 26 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.565 $Y=1.22
+ $X2=1.565 $Y2=1.22
r64 23 24 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.537 $Y=2.945
+ $X2=1.537 $Y2=3.115
r65 19 21 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=1.565 $Y=3.205
+ $X2=1.565 $Y2=4.565
r66 19 24 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=1.565 $Y=3.205
+ $X2=1.565 $Y2=3.115
r67 13 26 9.13816 $w=3.4e-07 $l=2.35e-07 $layer=LI1_cond $X=1.565 $Y=0.985
+ $X2=1.565 $Y2=1.22
r68 13 15 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.565 $Y=0.985
+ $X2=1.565 $Y2=0.865
r69 11 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=2.33
+ $X2=1.425 $Y2=2.33
r70 11 23 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.425 $Y=2.33
+ $X2=1.425 $Y2=2.945
r71 3 21 240 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.565 $Y2=4.565
r72 3 19 240 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.565 $Y2=3.205
r73 1 15 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.865
.ends

