* File: sky130_osu_sc_12T_ls__xnor2_l.spice
* Created: Fri Nov 12 15:41:06 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__xnor2_l.pex.spice"
.subckt sky130_osu_sc_12T_ls__xnor2_l  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75002.4 A=0.078 P=1.34 MULT=1
MM1000 A_196_115# N_A_M1000_g N_GND_M1004_d N_GND_M1004_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1009 N_Y_M1009_d N_A_238_89#_M1009_g A_196_115# N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1006 A_388_115# N_A_27_115#_M1006_g N_Y_M1009_d N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_B_M1007_g A_388_115# N_GND_M1004_b NSHORT L=0.15 W=0.52
+ AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75001.9
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1005 N_A_238_89#_M1005_d N_B_M1005_g N_GND_M1007_d N_GND_M1004_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75002.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g N_A_27_115#_M1003_s N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1010 A_196_521# N_A_27_115#_M1010_g N_VDD_M1003_d N_VDD_M1003_b PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_A_238_89#_M1011_g A_196_521# N_VDD_M1003_b PHIGHVT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1001 A_388_521# N_A_M1001_g N_Y_M1011_d N_VDD_M1003_b PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1002 N_VDD_M1002_d N_B_M1002_g A_388_521# N_VDD_M1003_b PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_238_89#_M1008_d N_B_M1008_g N_VDD_M1002_d N_VDD_M1003_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1004_b N_VDD_M1003_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_12 A A PROBETYPE=1
pX14_noxref noxref_13 Y Y PROBETYPE=1
pX15_noxref noxref_14 B B PROBETYPE=1
c_503 A_388_115# 0 1.09094e-19 $X=1.94 $Y=0.575
*
.include "sky130_osu_sc_12T_ls__xnor2_l.pxi.spice"
*
.ends
*
*
