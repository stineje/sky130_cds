magic
tech sky130A
magscale 1 2
timestamp 1612373432
<< nwell >>
rect -9 529 814 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 252 115 282 243
rect 338 115 368 243
rect 424 115 454 243
rect 510 115 540 243
rect 596 115 626 243
rect 682 115 712 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
rect 338 565 368 965
rect 424 565 454 965
rect 510 565 540 965
rect 596 565 626 965
rect 682 565 712 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 166 243
rect 110 131 121 215
rect 155 131 166 215
rect 110 115 166 131
rect 196 215 252 243
rect 196 131 207 215
rect 241 131 252 215
rect 196 115 252 131
rect 282 215 338 243
rect 282 131 293 215
rect 327 131 338 215
rect 282 115 338 131
rect 368 215 424 243
rect 368 131 379 215
rect 413 131 424 215
rect 368 115 424 131
rect 454 215 510 243
rect 454 131 465 215
rect 499 131 510 215
rect 454 115 510 131
rect 540 215 596 243
rect 540 131 551 215
rect 585 131 596 215
rect 540 115 596 131
rect 626 215 682 243
rect 626 131 637 215
rect 671 131 682 215
rect 626 115 682 131
rect 712 215 765 243
rect 712 131 723 215
rect 757 131 765 215
rect 712 115 765 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 949 166 965
rect 110 605 121 949
rect 155 605 166 949
rect 110 565 166 605
rect 196 949 252 965
rect 196 605 207 949
rect 241 605 252 949
rect 196 565 252 605
rect 282 949 338 965
rect 282 605 293 949
rect 327 605 338 949
rect 282 565 338 605
rect 368 949 424 965
rect 368 605 379 949
rect 413 605 424 949
rect 368 565 424 605
rect 454 949 510 965
rect 454 605 465 949
rect 499 605 510 949
rect 454 565 510 605
rect 540 949 596 965
rect 540 605 551 949
rect 585 605 596 949
rect 540 565 596 605
rect 626 949 682 965
rect 626 605 637 949
rect 671 605 682 949
rect 626 565 682 605
rect 712 949 765 965
rect 712 605 723 949
rect 757 605 765 949
rect 712 565 765 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 207 131 241 215
rect 293 131 327 215
rect 379 131 413 215
rect 465 131 499 215
rect 551 131 585 215
rect 637 131 671 215
rect 723 131 757 215
<< pdiffc >>
rect 35 741 69 949
rect 121 605 155 949
rect 207 605 241 949
rect 293 605 327 949
rect 379 605 413 949
rect 465 605 499 949
rect 551 605 585 949
rect 637 605 671 949
rect 723 605 757 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
rect 571 1049 595 1083
rect 629 1049 653 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
rect 595 1049 629 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 991
rect 338 965 368 991
rect 424 965 454 991
rect 510 965 540 991
rect 596 965 626 991
rect 682 965 712 991
rect 80 540 110 565
rect 166 540 196 565
rect 252 540 282 565
rect 338 540 368 565
rect 424 540 454 565
rect 510 540 540 565
rect 596 540 626 565
rect 682 540 712 565
rect 80 510 712 540
rect 80 442 110 510
rect 80 426 134 442
rect 80 392 90 426
rect 124 392 134 426
rect 80 376 134 392
rect 80 318 110 376
rect 424 318 454 510
rect 80 288 712 318
rect 80 243 110 288
rect 166 243 196 288
rect 252 243 282 288
rect 338 243 368 288
rect 424 243 454 288
rect 510 243 540 288
rect 596 243 626 288
rect 682 243 712 288
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
rect 338 89 368 115
rect 424 89 454 115
rect 510 89 540 115
rect 596 89 626 115
rect 682 89 712 115
<< polycont >>
rect 90 392 124 426
<< locali >>
rect 0 1089 814 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 595 1089
rect 629 1049 814 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 121 949 155 965
rect 47 426 81 597
rect 121 557 155 605
rect 207 949 241 1049
rect 207 589 241 605
rect 293 949 327 965
rect 293 557 327 605
rect 379 949 413 1049
rect 379 589 413 605
rect 465 949 499 965
rect 465 557 499 605
rect 551 949 585 1049
rect 551 589 585 605
rect 637 949 671 965
rect 637 557 671 605
rect 723 949 757 1049
rect 723 589 757 605
rect 47 392 90 426
rect 124 392 140 426
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 227
rect 121 115 155 131
rect 207 215 241 231
rect 207 61 241 131
rect 293 215 327 227
rect 293 115 327 131
rect 379 215 413 231
rect 379 61 413 131
rect 465 215 499 227
rect 465 115 499 131
rect 551 215 585 231
rect 551 61 585 131
rect 637 215 671 227
rect 637 115 671 131
rect 723 215 757 231
rect 723 61 757 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 814 61
rect 0 0 814 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 595 1083 629 1089
rect 595 1055 629 1083
rect 47 597 81 631
rect 121 523 155 557
rect 293 523 327 557
rect 465 523 499 557
rect 637 523 671 557
rect 121 227 155 261
rect 293 227 327 261
rect 465 227 499 261
rect 637 227 671 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
<< metal1 >>
rect 0 1089 814 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 595 1089
rect 629 1055 814 1089
rect 0 1049 814 1055
rect 35 631 93 637
rect 35 597 47 631
rect 81 597 127 631
rect 35 591 93 597
rect 109 557 167 563
rect 281 557 339 563
rect 453 557 511 563
rect 625 557 683 563
rect 109 523 121 557
rect 155 523 293 557
rect 327 523 465 557
rect 499 523 637 557
rect 671 523 683 557
rect 109 517 167 523
rect 281 517 339 523
rect 453 517 511 523
rect 625 517 683 523
rect 121 267 155 517
rect 293 267 327 517
rect 465 267 499 517
rect 637 267 671 517
rect 109 261 167 267
rect 281 261 339 267
rect 453 261 511 267
rect 625 261 683 267
rect 109 227 121 261
rect 155 227 293 261
rect 327 227 465 261
rect 499 227 637 261
rect 671 227 683 261
rect 109 221 167 227
rect 281 221 339 227
rect 453 221 511 227
rect 625 221 683 227
rect 0 55 814 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 814 55
rect 0 0 814 21
<< labels >>
rlabel metal1 152 388 152 388 1 Y
port 1 n
rlabel viali 64 613 64 613 1 A
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
