* File: sky130_osu_sc_12T_ms__tnbufi_l.pxi.spice
* Created: Fri Nov 12 15:27:27 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_6_p
+ N_GND_c_2_p GND N_GND_c_3_p PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%GND
x_PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_33_p
+ N_VDD_c_37_p N_VDD_c_38_p VDD N_VDD_c_34_p
+ PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_c_52_n N_A_27_115#_c_53_n
+ N_A_27_115#_c_56_n N_A_27_115#_c_57_n N_A_27_115#_c_58_n N_A_27_115#_c_59_n
+ PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%OE N_OE_M1002_g N_OE_c_94_n N_OE_M1001_g
+ N_OE_M1005_g N_OE_c_95_n N_OE_c_96_n OE PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%OE
x_PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%A N_A_M1004_g N_A_M1003_g N_A_c_135_n
+ N_A_c_136_n A PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%A
x_PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%Y N_Y_M1004_d N_Y_M1003_d N_Y_c_168_n
+ N_Y_c_170_n Y N_Y_c_172_n N_Y_c_173_n PM_SKY130_OSU_SC_12T_MS__TNBUFI_L%Y
cc_1 N_GND_M1002_b N_A_27_115#_M1000_g 0.0674434f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.755
cc_2 N_GND_c_2_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905
+ $Y2=0.755
cc_3 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=0.755
cc_4 N_GND_M1002_b N_A_27_115#_c_52_n 0.0424934f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=2.06
cc_5 N_GND_M1002_b N_A_27_115#_c_53_n 0.0453036f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_6 N_GND_c_6_p N_A_27_115#_c_53_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_7 N_GND_c_3_p N_A_27_115#_c_53_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_8 N_GND_M1002_b N_A_27_115#_c_56_n 0.0221237f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.275
cc_9 N_GND_M1002_b N_A_27_115#_c_57_n 0.00869964f $X=-0.045 $Y=0 $X2=0.605
+ $Y2=2.062
cc_10 N_GND_M1002_b N_A_27_115#_c_58_n 0.00666352f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.062
cc_11 N_GND_M1002_b N_A_27_115#_c_59_n 0.00712065f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=2.06
cc_12 N_GND_M1002_b N_OE_M1002_g 0.0482623f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.755
cc_13 N_GND_c_6_p N_OE_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.755
cc_14 N_GND_c_2_p N_OE_M1002_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.755
cc_15 N_GND_c_3_p N_OE_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.755
cc_16 N_GND_M1002_b N_OE_c_94_n 0.0986588f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.9
cc_17 N_GND_M1002_b N_OE_c_95_n 0.0253092f $X=-0.045 $Y=0 $X2=0.27 $Y2=1.61
cc_18 N_GND_M1002_b N_OE_c_96_n 0.00225456f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.48
cc_19 N_GND_M1002_b OE 0.0102226f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.485
cc_20 N_GND_M1002_b N_A_M1004_g 0.0740802f $X=-0.045 $Y=0 $X2=1.265 $Y2=0.755
cc_21 N_GND_c_3_p N_A_M1004_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.265 $Y2=0.755
cc_22 N_GND_M1002_b N_A_M1003_g 0.0492565f $X=-0.045 $Y=0 $X2=1.265 $Y2=3.445
cc_23 N_GND_M1002_b N_A_c_135_n 0.032012f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.98
cc_24 N_GND_M1002_b N_A_c_136_n 0.0112497f $X=-0.045 $Y=0 $X2=1.14 $Y2=2.11
cc_25 N_GND_M1002_b A 0.0110418f $X=-0.045 $Y=0 $X2=1.14 $Y2=2.115
cc_26 N_GND_M1002_b N_Y_c_168_n 0.0330266f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.74
cc_27 N_GND_c_3_p N_Y_c_168_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.48 $Y2=0.74
cc_28 N_GND_M1002_b N_Y_c_170_n 0.00301383f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.85
cc_29 N_GND_M1002_b Y 0.0596048f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.71
cc_30 N_GND_M1002_b N_Y_c_172_n 0.00481997f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.85
cc_31 N_GND_M1002_b N_Y_c_173_n 0.0151505f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.37
cc_32 N_VDD_M1001_b N_A_27_115#_c_56_n 0.010588f $X=-0.045 $Y=2.795 $X2=0.26
+ $Y2=3.275
cc_33 N_VDD_c_33_p N_A_27_115#_c_56_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=3.275
cc_34 N_VDD_c_34_p N_A_27_115#_c_56_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26
+ $Y2=3.275
cc_35 N_VDD_M1001_b N_OE_c_94_n 0.0608086f $X=-0.045 $Y=2.795 $X2=0.475 $Y2=2.9
cc_36 N_VDD_c_33_p N_OE_c_94_n 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=2.9
cc_37 N_VDD_c_37_p N_OE_c_94_n 0.00972025f $X=0.69 $Y=3.275 $X2=0.475 $Y2=2.9
cc_38 N_VDD_c_38_p N_OE_c_94_n 0.00606474f $X=1.02 $Y=4.22 $X2=0.475 $Y2=2.9
cc_39 N_VDD_c_34_p N_OE_c_94_n 0.00937653f $X=1.02 $Y=4.25 $X2=0.475 $Y2=2.9
cc_40 N_VDD_c_37_p N_OE_c_96_n 0.0113232f $X=0.69 $Y=3.275 $X2=0.69 $Y2=2.48
cc_41 N_VDD_c_37_p OE 8.88903e-19 $X=0.69 $Y=3.275 $X2=0.69 $Y2=2.485
cc_42 N_VDD_M1001_b N_A_M1003_g 0.0286218f $X=-0.045 $Y=2.795 $X2=1.265
+ $Y2=3.445
cc_43 N_VDD_c_38_p N_A_M1003_g 0.00606474f $X=1.02 $Y=4.22 $X2=1.265 $Y2=3.445
cc_44 N_VDD_c_34_p N_A_M1003_g 0.00468827f $X=1.02 $Y=4.25 $X2=1.265 $Y2=3.445
cc_45 N_VDD_M1001_b N_Y_c_170_n 0.00984349f $X=-0.045 $Y=2.795 $X2=1.48 $Y2=2.85
cc_46 N_VDD_c_38_p N_Y_c_170_n 0.00757793f $X=1.02 $Y=4.22 $X2=1.48 $Y2=2.85
cc_47 N_VDD_c_34_p N_Y_c_170_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.48 $Y2=2.85
cc_48 N_VDD_M1001_b N_Y_c_172_n 0.0109393f $X=-0.045 $Y=2.795 $X2=1.48 $Y2=2.85
cc_49 N_A_27_115#_M1000_g N_OE_M1002_g 0.0398172f $X=0.905 $Y=0.755 $X2=0.475
+ $Y2=0.755
cc_50 N_A_27_115#_c_53_n N_OE_M1002_g 0.0232482f $X=0.26 $Y=0.74 $X2=0.475
+ $Y2=0.755
cc_51 N_A_27_115#_M1000_g N_OE_c_94_n 0.00301188f $X=0.905 $Y=0.755 $X2=0.475
+ $Y2=2.9
cc_52 N_A_27_115#_c_52_n N_OE_c_94_n 0.0386296f $X=0.905 $Y=2.06 $X2=0.475
+ $Y2=2.9
cc_53 N_A_27_115#_c_53_n N_OE_c_94_n 0.0121188f $X=0.26 $Y=0.74 $X2=0.475
+ $Y2=2.9
cc_54 N_A_27_115#_c_56_n N_OE_c_94_n 0.0476448f $X=0.26 $Y=3.275 $X2=0.475
+ $Y2=2.9
cc_55 N_A_27_115#_c_57_n N_OE_c_94_n 0.00105571f $X=0.605 $Y=2.062 $X2=0.475
+ $Y2=2.9
cc_56 N_A_27_115#_c_58_n N_OE_c_94_n 0.0065159f $X=0.26 $Y=2.062 $X2=0.475
+ $Y2=2.9
cc_57 N_A_27_115#_c_59_n N_OE_c_94_n 5.30096e-19 $X=0.69 $Y=2.06 $X2=0.475
+ $Y2=2.9
cc_58 N_A_27_115#_c_53_n N_OE_c_95_n 0.0104412f $X=0.26 $Y=0.74 $X2=0.27
+ $Y2=1.61
cc_59 N_A_27_115#_c_57_n N_OE_c_95_n 0.007138f $X=0.605 $Y=2.062 $X2=0.27
+ $Y2=1.61
cc_60 N_A_27_115#_c_52_n N_OE_c_96_n 4.76915e-19 $X=0.905 $Y=2.06 $X2=0.69
+ $Y2=2.48
cc_61 N_A_27_115#_c_56_n N_OE_c_96_n 0.0184316f $X=0.26 $Y=3.275 $X2=0.69
+ $Y2=2.48
cc_62 N_A_27_115#_c_59_n N_OE_c_96_n 0.011291f $X=0.69 $Y=2.06 $X2=0.69 $Y2=2.48
cc_63 N_A_27_115#_c_52_n OE 0.00302464f $X=0.905 $Y=2.06 $X2=0.69 $Y2=2.485
cc_64 N_A_27_115#_c_56_n OE 0.00724876f $X=0.26 $Y=3.275 $X2=0.69 $Y2=2.485
cc_65 N_A_27_115#_c_57_n OE 0.00255622f $X=0.605 $Y=2.062 $X2=0.69 $Y2=2.485
cc_66 N_A_27_115#_c_59_n OE 0.00476179f $X=0.69 $Y=2.06 $X2=0.69 $Y2=2.485
cc_67 N_A_27_115#_M1000_g N_A_M1004_g 0.0560234f $X=0.905 $Y=0.755 $X2=1.265
+ $Y2=0.755
cc_68 N_A_27_115#_c_52_n N_A_c_135_n 0.0560234f $X=0.905 $Y=2.06 $X2=1.325
+ $Y2=1.98
cc_69 N_A_27_115#_c_59_n N_A_c_135_n 2.32787e-19 $X=0.69 $Y=2.06 $X2=1.325
+ $Y2=1.98
cc_70 N_A_27_115#_c_52_n N_A_c_136_n 0.00227635f $X=0.905 $Y=2.06 $X2=1.14
+ $Y2=2.11
cc_71 N_A_27_115#_c_59_n N_A_c_136_n 0.0125821f $X=0.69 $Y=2.06 $X2=1.14
+ $Y2=2.11
cc_72 N_A_27_115#_c_52_n A 0.00865145f $X=0.905 $Y=2.06 $X2=1.14 $Y2=2.115
cc_73 N_A_27_115#_c_59_n A 0.00712629f $X=0.69 $Y=2.06 $X2=1.14 $Y2=2.115
cc_74 N_A_27_115#_M1000_g Y 3.12481e-19 $X=0.905 $Y=0.755 $X2=1.525 $Y2=1.71
cc_75 N_A_27_115#_M1000_g N_Y_c_173_n 0.00101819f $X=0.905 $Y=0.755 $X2=1.48
+ $Y2=1.37
cc_76 N_OE_c_94_n N_A_M1003_g 0.0836451f $X=0.475 $Y=2.9 $X2=1.265 $Y2=3.445
cc_77 N_OE_c_96_n N_A_M1003_g 0.00401208f $X=0.69 $Y=2.48 $X2=1.265 $Y2=3.445
cc_78 OE N_A_M1003_g 0.00290931f $X=0.69 $Y=2.485 $X2=1.265 $Y2=3.445
cc_79 N_OE_c_94_n A 2.29672e-19 $X=0.475 $Y=2.9 $X2=1.14 $Y2=2.115
cc_80 OE A 0.00500902f $X=0.69 $Y=2.485 $X2=1.14 $Y2=2.115
cc_81 N_OE_c_96_n N_Y_c_170_n 7.96059e-19 $X=0.69 $Y=2.48 $X2=1.48 $Y2=2.85
cc_82 OE Y 0.00979631f $X=0.69 $Y=2.485 $X2=1.525 $Y2=1.71
cc_83 N_OE_c_94_n N_Y_c_172_n 0.00114645f $X=0.475 $Y=2.9 $X2=1.48 $Y2=2.85
cc_84 N_OE_c_96_n N_Y_c_172_n 0.00179938f $X=0.69 $Y=2.48 $X2=1.48 $Y2=2.85
cc_85 N_A_M1004_g N_Y_c_168_n 0.0190376f $X=1.265 $Y=0.755 $X2=1.48 $Y2=0.74
cc_86 N_A_c_135_n N_Y_c_168_n 0.00104136f $X=1.325 $Y=1.98 $X2=1.48 $Y2=0.74
cc_87 N_A_c_136_n N_Y_c_168_n 0.00231375f $X=1.14 $Y=2.11 $X2=1.48 $Y2=0.74
cc_88 N_A_M1003_g N_Y_c_170_n 0.010524f $X=1.265 $Y=3.445 $X2=1.48 $Y2=2.85
cc_89 N_A_c_135_n N_Y_c_170_n 0.00107704f $X=1.325 $Y=1.98 $X2=1.48 $Y2=2.85
cc_90 N_A_M1004_g Y 0.00755346f $X=1.265 $Y=0.755 $X2=1.525 $Y2=1.71
cc_91 N_A_M1003_g Y 0.0113754f $X=1.265 $Y=3.445 $X2=1.525 $Y2=1.71
cc_92 N_A_c_135_n Y 0.00454161f $X=1.325 $Y=1.98 $X2=1.525 $Y2=1.71
cc_93 N_A_c_136_n Y 0.0137711f $X=1.14 $Y=2.11 $X2=1.525 $Y2=1.71
cc_94 A Y 0.0229562f $X=1.14 $Y=2.115 $X2=1.525 $Y2=1.71
cc_95 N_A_M1003_g N_Y_c_172_n 0.00729937f $X=1.265 $Y=3.445 $X2=1.48 $Y2=2.85
cc_96 N_A_c_135_n N_Y_c_172_n 0.00172008f $X=1.325 $Y=1.98 $X2=1.48 $Y2=2.85
cc_97 N_A_M1004_g N_Y_c_173_n 0.00707701f $X=1.265 $Y=0.755 $X2=1.48 $Y2=1.37
cc_98 N_A_c_135_n N_Y_c_173_n 0.0020015f $X=1.325 $Y=1.98 $X2=1.48 $Y2=1.37
cc_99 N_A_c_136_n N_Y_c_173_n 0.00274303f $X=1.14 $Y=2.11 $X2=1.48 $Y2=1.37
