* File: sky130_osu_sc_12T_hs__or2_2.pxi.spice
* Created: Fri Nov 12 15:12:43 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__OR2_2%GND N_GND_M1004_s N_GND_M1001_d N_GND_M1007_s
+ N_GND_M1004_b N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p N_GND_c_24_p
+ GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_HS__OR2_2%GND
x_PM_SKY130_OSU_SC_12T_HS__OR2_2%VDD N_VDD_M1005_d N_VDD_M1006_d N_VDD_M1000_b
+ N_VDD_c_45_p N_VDD_c_51_p N_VDD_c_58_p N_VDD_c_64_p VDD N_VDD_c_46_p
+ PM_SKY130_OSU_SC_12T_HS__OR2_2%VDD
x_PM_SKY130_OSU_SC_12T_HS__OR2_2%B N_B_M1004_g N_B_M1000_g N_B_c_79_n N_B_c_80_n
+ B PM_SKY130_OSU_SC_12T_HS__OR2_2%B
x_PM_SKY130_OSU_SC_12T_HS__OR2_2%A N_A_M1001_g N_A_M1005_g N_A_c_107_n
+ N_A_c_108_n A PM_SKY130_OSU_SC_12T_HS__OR2_2%A
x_PM_SKY130_OSU_SC_12T_HS__OR2_2%A_27_521# N_A_27_521#_M1004_d
+ N_A_27_521#_M1000_s N_A_27_521#_M1002_g N_A_27_521#_c_165_n
+ N_A_27_521#_M1003_g N_A_27_521#_c_150_n N_A_27_521#_c_151_n
+ N_A_27_521#_M1007_g N_A_27_521#_c_170_n N_A_27_521#_M1006_g
+ N_A_27_521#_c_156_n N_A_27_521#_c_157_n N_A_27_521#_c_176_n
+ N_A_27_521#_c_180_n N_A_27_521#_c_182_n N_A_27_521#_c_158_n
+ N_A_27_521#_c_159_n N_A_27_521#_c_162_n N_A_27_521#_c_164_n
+ PM_SKY130_OSU_SC_12T_HS__OR2_2%A_27_521#
x_PM_SKY130_OSU_SC_12T_HS__OR2_2%Y N_Y_M1002_d N_Y_M1003_s N_Y_c_236_n
+ N_Y_c_239_n Y N_Y_c_241_n N_Y_c_244_n PM_SKY130_OSU_SC_12T_HS__OR2_2%Y
cc_1 N_GND_M1004_b N_B_M1004_g 0.0813622f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_B_M1004_g 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_B_M1004_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.85
cc_4 N_GND_c_4_p N_B_M1004_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=0.85
cc_5 N_GND_M1004_b N_B_M1000_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_6 N_GND_M1004_b N_B_c_79_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.195
cc_7 N_GND_M1004_b N_B_c_80_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.195
cc_8 N_GND_M1004_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.48
cc_9 N_GND_M1004_b N_A_M1001_g 0.0424425f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.85
cc_10 N_GND_c_3_p N_A_M1001_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.85
cc_11 N_GND_c_11_p N_A_M1001_g 0.00308284f $X=1.12 $Y=0.755 $X2=0.905 $Y2=0.85
cc_12 N_GND_c_4_p N_A_M1001_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.905 $Y2=0.85
cc_13 N_GND_M1004_b N_A_M1005_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_14 N_GND_M1004_b N_A_c_107_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.905
cc_15 N_GND_M1004_b N_A_c_108_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.905
cc_16 N_GND_M1004_b N_A_27_521#_M1002_g 0.0192558f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.85
cc_17 N_GND_c_11_p N_A_27_521#_M1002_g 0.00308284f $X=1.12 $Y=0.755 $X2=1.335
+ $Y2=0.85
cc_18 N_GND_c_18_p N_A_27_521#_M1002_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.85
cc_19 N_GND_c_4_p N_A_27_521#_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335
+ $Y2=0.85
cc_20 N_GND_M1004_b N_A_27_521#_c_150_n 0.0466273f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.33
cc_21 N_GND_M1004_b N_A_27_521#_c_151_n 0.0244031f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.405
cc_22 N_GND_M1004_b N_A_27_521#_M1007_g 0.0241608f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.85
cc_23 N_GND_c_18_p N_A_27_521#_M1007_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.85
cc_24 N_GND_c_24_p N_A_27_521#_M1007_g 0.00502587f $X=1.98 $Y=0.755 $X2=1.765
+ $Y2=0.85
cc_25 N_GND_c_4_p N_A_27_521#_M1007_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765
+ $Y2=0.85
cc_26 N_GND_M1004_b N_A_27_521#_c_156_n 0.00567173f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.405
cc_27 N_GND_M1004_b N_A_27_521#_c_157_n 0.0539419f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_28 N_GND_M1004_b N_A_27_521#_c_158_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.065
cc_29 N_GND_M1004_b N_A_27_521#_c_159_n 0.00637039f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.755
cc_30 N_GND_c_3_p N_A_27_521#_c_159_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.755
cc_31 N_GND_c_4_p N_A_27_521#_c_159_n 0.00475776f $X=1.7 $Y=0.19 $X2=0.69
+ $Y2=0.755
cc_32 N_GND_M1004_b N_A_27_521#_c_162_n 0.0190355f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_33 N_GND_c_11_p N_A_27_521#_c_162_n 0.00702738f $X=1.12 $Y=0.755 $X2=1.43
+ $Y2=1.455
cc_34 N_GND_M1004_b N_A_27_521#_c_164_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.455
cc_35 N_GND_M1004_b N_Y_c_236_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_36 N_GND_c_18_p N_Y_c_236_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_37 N_GND_c_4_p N_Y_c_236_n 0.0047139f $X=1.7 $Y=0.19 $X2=1.55 $Y2=0.755
cc_38 N_GND_M1004_b N_Y_c_239_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_39 N_GND_M1004_b Y 0.0304196f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.74
cc_40 N_GND_c_11_p N_Y_c_241_n 0.00125659f $X=1.12 $Y=0.755 $X2=1.55 $Y2=1
cc_41 N_GND_c_18_p N_Y_c_241_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.55 $Y2=1
cc_42 N_GND_c_24_p N_Y_c_241_n 0.00125659f $X=1.98 $Y=0.755 $X2=1.55 $Y2=1
cc_43 N_GND_M1004_b N_Y_c_244_n 0.0111067f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_44 N_VDD_M1000_b N_B_M1000_g 0.0260091f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_45 N_VDD_c_45_p N_B_M1000_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.235
cc_46 N_VDD_c_46_p N_B_M1000_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.475 $Y2=3.235
cc_47 N_VDD_M1000_b N_B_c_80_n 0.00375034f $X=-0.045 $Y=2.425 $X2=0.27 $Y2=2.195
cc_48 N_VDD_M1000_b B 0.0108395f $X=-0.045 $Y=2.425 $X2=0.27 $Y2=2.48
cc_49 N_VDD_M1000_b N_A_M1005_g 0.0195137f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_50 N_VDD_c_45_p N_A_M1005_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.235
cc_51 N_VDD_c_51_p N_A_M1005_g 0.00337744f $X=1.12 $Y=3.635 $X2=0.905 $Y2=3.235
cc_52 N_VDD_c_46_p N_A_M1005_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.905 $Y2=3.235
cc_53 N_VDD_M1000_b N_A_c_108_n 0.00153494f $X=-0.045 $Y=2.425 $X2=0.95
+ $Y2=1.905
cc_54 N_VDD_M1005_d A 0.0077995f $X=0.98 $Y=2.605 $X2=0.95 $Y2=2.85
cc_55 N_VDD_c_51_p A 0.00247404f $X=1.12 $Y=3.635 $X2=0.95 $Y2=2.85
cc_56 N_VDD_M1000_b N_A_27_521#_c_165_n 0.0170965f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.48
cc_57 N_VDD_c_51_p N_A_27_521#_c_165_n 0.00337744f $X=1.12 $Y=3.635 $X2=1.335
+ $Y2=2.48
cc_58 N_VDD_c_58_p N_A_27_521#_c_165_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335
+ $Y2=2.48
cc_59 N_VDD_c_46_p N_A_27_521#_c_165_n 0.00468827f $X=1.7 $Y=4.25 $X2=1.335
+ $Y2=2.48
cc_60 N_VDD_M1000_b N_A_27_521#_c_151_n 0.00813142f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_61 N_VDD_M1000_b N_A_27_521#_c_170_n 0.0212198f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.48
cc_62 N_VDD_c_51_p N_A_27_521#_c_170_n 3.67508e-19 $X=1.12 $Y=3.635 $X2=1.765
+ $Y2=2.48
cc_63 N_VDD_c_58_p N_A_27_521#_c_170_n 0.00610567f $X=1.895 $Y=4.287 $X2=1.765
+ $Y2=2.48
cc_64 N_VDD_c_64_p N_A_27_521#_c_170_n 0.00656078f $X=1.98 $Y=2.955 $X2=1.765
+ $Y2=2.48
cc_65 N_VDD_c_46_p N_A_27_521#_c_170_n 0.00470215f $X=1.7 $Y=4.25 $X2=1.765
+ $Y2=2.48
cc_66 N_VDD_M1000_b N_A_27_521#_c_156_n 0.00216365f $X=-0.045 $Y=2.425 $X2=1.352
+ $Y2=2.405
cc_67 N_VDD_M1000_b N_A_27_521#_c_176_n 0.00156053f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=3.295
cc_68 N_VDD_c_45_p N_A_27_521#_c_176_n 0.00736239f $X=1.035 $Y=4.287 $X2=0.26
+ $Y2=3.295
cc_69 N_VDD_c_46_p N_A_27_521#_c_176_n 0.00476261f $X=1.7 $Y=4.25 $X2=0.26
+ $Y2=3.295
cc_70 N_VDD_M1000_b N_A_27_521#_c_158_n 0.00106577f $X=-0.045 $Y=2.425 $X2=0.61
+ $Y2=3.065
cc_71 N_VDD_M1000_b N_Y_c_239_n 0.00367096f $X=-0.045 $Y=2.425 $X2=1.55 $Y2=2.11
cc_72 N_VDD_c_58_p N_Y_c_239_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.11
cc_73 N_VDD_c_46_p N_Y_c_239_n 0.00475776f $X=1.7 $Y=4.25 $X2=1.55 $Y2=2.11
cc_74 N_B_M1004_g N_A_M1001_g 0.0358421f $X=0.475 $Y=0.85 $X2=0.905 $Y2=0.85
cc_75 N_B_c_79_n N_A_M1005_g 0.0819064f $X=0.475 $Y=2.195 $X2=0.905 $Y2=3.235
cc_76 N_B_M1004_g N_A_c_107_n 0.0148656f $X=0.475 $Y=0.85 $X2=0.95 $Y2=1.905
cc_77 N_B_M1004_g N_A_c_108_n 0.00121111f $X=0.475 $Y=0.85 $X2=0.95 $Y2=1.905
cc_78 N_B_M1000_g N_A_27_521#_c_180_n 0.0136492f $X=0.475 $Y=3.235 $X2=0.525
+ $Y2=3.15
cc_79 B N_A_27_521#_c_180_n 0.00520961f $X=0.27 $Y=2.48 $X2=0.525 $Y2=3.15
cc_80 N_B_c_80_n N_A_27_521#_c_182_n 0.00369517f $X=0.27 $Y=2.195 $X2=0.345
+ $Y2=3.15
cc_81 B N_A_27_521#_c_182_n 0.00431991f $X=0.27 $Y=2.48 $X2=0.345 $Y2=3.15
cc_82 N_B_M1004_g N_A_27_521#_c_158_n 0.0231435f $X=0.475 $Y=0.85 $X2=0.61
+ $Y2=3.065
cc_83 N_B_M1000_g N_A_27_521#_c_158_n 0.026563f $X=0.475 $Y=3.235 $X2=0.61
+ $Y2=3.065
cc_84 N_B_c_79_n N_A_27_521#_c_158_n 0.00764878f $X=0.475 $Y=2.195 $X2=0.61
+ $Y2=3.065
cc_85 N_B_c_80_n N_A_27_521#_c_158_n 0.0350086f $X=0.27 $Y=2.195 $X2=0.61
+ $Y2=3.065
cc_86 B N_A_27_521#_c_158_n 0.00758489f $X=0.27 $Y=2.48 $X2=0.61 $Y2=3.065
cc_87 N_B_M1004_g N_A_27_521#_c_159_n 0.00654421f $X=0.475 $Y=0.85 $X2=0.69
+ $Y2=0.755
cc_88 N_B_M1004_g N_A_27_521#_c_164_n 0.0113001f $X=0.475 $Y=0.85 $X2=0.65
+ $Y2=1.455
cc_89 N_A_M1001_g N_A_27_521#_M1002_g 0.0264543f $X=0.905 $Y=0.85 $X2=1.335
+ $Y2=0.85
cc_90 A N_A_27_521#_c_165_n 0.00374181f $X=0.95 $Y=2.85 $X2=1.335 $Y2=2.48
cc_91 N_A_M1005_g N_A_27_521#_c_150_n 0.00914307f $X=0.905 $Y=3.235 $X2=1.37
+ $Y2=2.33
cc_92 N_A_c_107_n N_A_27_521#_c_150_n 0.0204279f $X=0.95 $Y=1.905 $X2=1.37
+ $Y2=2.33
cc_93 N_A_c_108_n N_A_27_521#_c_150_n 0.00375034f $X=0.95 $Y=1.905 $X2=1.37
+ $Y2=2.33
cc_94 N_A_M1005_g N_A_27_521#_c_156_n 0.0532043f $X=0.905 $Y=3.235 $X2=1.352
+ $Y2=2.405
cc_95 N_A_c_108_n N_A_27_521#_c_156_n 0.00355256f $X=0.95 $Y=1.905 $X2=1.352
+ $Y2=2.405
cc_96 N_A_M1001_g N_A_27_521#_c_157_n 0.0119161f $X=0.905 $Y=0.85 $X2=1.43
+ $Y2=1.455
cc_97 N_A_M1005_g N_A_27_521#_c_180_n 0.00457566f $X=0.905 $Y=3.235 $X2=0.525
+ $Y2=3.15
cc_98 N_A_M1001_g N_A_27_521#_c_158_n 0.00429604f $X=0.905 $Y=0.85 $X2=0.61
+ $Y2=3.065
cc_99 N_A_M1005_g N_A_27_521#_c_158_n 0.00776428f $X=0.905 $Y=3.235 $X2=0.61
+ $Y2=3.065
cc_100 N_A_c_107_n N_A_27_521#_c_158_n 0.0021255f $X=0.95 $Y=1.905 $X2=0.61
+ $Y2=3.065
cc_101 N_A_c_108_n N_A_27_521#_c_158_n 0.0822139f $X=0.95 $Y=1.905 $X2=0.61
+ $Y2=3.065
cc_102 A N_A_27_521#_c_158_n 0.00866797f $X=0.95 $Y=2.85 $X2=0.61 $Y2=3.065
cc_103 N_A_M1001_g N_A_27_521#_c_159_n 0.00654421f $X=0.905 $Y=0.85 $X2=0.69
+ $Y2=0.755
cc_104 N_A_M1001_g N_A_27_521#_c_162_n 0.0163305f $X=0.905 $Y=0.85 $X2=1.43
+ $Y2=1.455
cc_105 N_A_c_107_n N_A_27_521#_c_162_n 0.00276813f $X=0.95 $Y=1.905 $X2=1.43
+ $Y2=1.455
cc_106 N_A_c_108_n N_A_27_521#_c_162_n 0.0114342f $X=0.95 $Y=1.905 $X2=1.43
+ $Y2=1.455
cc_107 A A_110_521# 0.0123256f $X=0.95 $Y=2.85 $X2=0.55 $Y2=2.605
cc_108 N_A_c_108_n N_Y_c_239_n 0.0206732f $X=0.95 $Y=1.905 $X2=1.55 $Y2=2.11
cc_109 A N_Y_c_239_n 0.00659455f $X=0.95 $Y=2.85 $X2=1.55 $Y2=2.11
cc_110 N_A_M1001_g Y 6.73508e-19 $X=0.905 $Y=0.85 $X2=1.555 $Y2=1.74
cc_111 N_A_c_108_n Y 0.00825539f $X=0.95 $Y=1.905 $X2=1.555 $Y2=1.74
cc_112 N_A_M1001_g N_Y_c_241_n 7.77582e-19 $X=0.905 $Y=0.85 $X2=1.55 $Y2=1
cc_113 N_A_c_107_n N_Y_c_244_n 3.65268e-19 $X=0.95 $Y=1.905 $X2=1.55 $Y2=2.11
cc_114 N_A_c_108_n N_Y_c_244_n 0.00535705f $X=0.95 $Y=1.905 $X2=1.55 $Y2=2.11
cc_115 N_A_27_521#_c_180_n A_110_521# 0.00613297f $X=0.525 $Y=3.15 $X2=0.55
+ $Y2=2.605
cc_116 N_A_27_521#_c_158_n A_110_521# 0.00377193f $X=0.61 $Y=3.065 $X2=0.55
+ $Y2=2.605
cc_117 N_A_27_521#_M1002_g N_Y_c_236_n 0.00182852f $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=0.755
cc_118 N_A_27_521#_M1007_g N_Y_c_236_n 0.00182852f $X=1.765 $Y=0.85 $X2=1.55
+ $Y2=0.755
cc_119 N_A_27_521#_c_157_n N_Y_c_236_n 0.0016986f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_120 N_A_27_521#_c_162_n N_Y_c_236_n 0.00498892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_121 N_A_27_521#_c_165_n N_Y_c_239_n 0.0020967f $X=1.335 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_122 N_A_27_521#_c_150_n N_Y_c_239_n 0.00744772f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_123 N_A_27_521#_c_151_n N_Y_c_239_n 0.0160452f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_124 N_A_27_521#_c_170_n N_Y_c_239_n 0.00375894f $X=1.765 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_125 N_A_27_521#_c_157_n N_Y_c_239_n 0.0013767f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_126 N_A_27_521#_c_162_n N_Y_c_239_n 0.00273485f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_127 N_A_27_521#_M1002_g Y 0.00251111f $X=1.335 $Y=0.85 $X2=1.555 $Y2=1.74
cc_128 N_A_27_521#_c_150_n Y 0.00892438f $X=1.37 $Y=2.33 $X2=1.555 $Y2=1.74
cc_129 N_A_27_521#_M1007_g Y 0.00251111f $X=1.765 $Y=0.85 $X2=1.555 $Y2=1.74
cc_130 N_A_27_521#_c_157_n Y 0.0120226f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_131 N_A_27_521#_c_162_n Y 0.0147088f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_132 N_A_27_521#_M1002_g N_Y_c_241_n 0.00466569f $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=1
cc_133 N_A_27_521#_M1007_g N_Y_c_241_n 0.0084691f $X=1.765 $Y=0.85 $X2=1.55
+ $Y2=1
cc_134 N_A_27_521#_c_162_n N_Y_c_241_n 0.00238892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1
cc_135 N_A_27_521#_c_150_n N_Y_c_244_n 0.00740115f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_136 N_A_27_521#_c_151_n N_Y_c_244_n 0.00229755f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_137 N_A_27_521#_c_157_n N_Y_c_244_n 0.00174847f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_138 N_A_27_521#_c_162_n N_Y_c_244_n 0.00181779f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
