* File: sky130_osu_sc_15T_hs__dffr_l.pex.spice
* Created: Fri Nov 12 14:29:19 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%GND 1 2 3 4 5 6 7 8 9 121 125 127 134
+ 136 143 152 154 164 166 176 178 185 187 194 196 203 230 232
c223 176 0 1.67294e-19 $X=6.09 $Y=0.865
c224 152 0 3.07193e-19 $X=2.59 $Y=0.865
c225 121 0 1.27355e-19 $X=-0.05 $Y=0
r226 230 232 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.175 $Y2=0.152
r227 205 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.152
+ $X2=8.85 $Y2=0.152
r228 201 226 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.152
r229 201 203 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.74
r230 196 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.152
+ $X2=8.85 $Y2=0.152
r231 192 194 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.74
r232 188 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.152
+ $X2=7.04 $Y2=0.152
r233 183 222 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.152
r234 183 185 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.74
r235 179 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.152
+ $X2=6.09 $Y2=0.152
r236 178 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.152
+ $X2=7.04 $Y2=0.152
r237 174 221 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.152
r238 174 176 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.865
r239 166 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.152
+ $X2=6.09 $Y2=0.152
r240 162 164 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.34 $Y=0.305
+ $X2=4.34 $Y2=0.74
r241 155 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.152
+ $X2=2.59 $Y2=0.152
r242 150 217 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.152
r243 150 152 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.865
r244 146 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.152
+ $X2=2.07 $Y2=0.152
r245 145 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.152
+ $X2=2.59 $Y2=0.152
r246 141 216 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.152
r247 141 143 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.74
r248 137 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.152
+ $X2=1.21 $Y2=0.152
r249 136 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.152
+ $X2=2.07 $Y2=0.152
r250 132 215 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.152
r251 132 134 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.74
r252 127 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.152
+ $X2=1.21 $Y2=0.152
r253 123 125 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r254 121 232 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=0.19 $X2=9.175 $Y2=0.19
r255 121 230 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=0.19 $X2=0.335 $Y2=0.19
r256 121 192 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r257 121 187 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r258 121 197 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.985 $Y2=0.152
r259 121 162 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.34 $Y2=0.305
r260 121 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.255 $Y2=0.152
r261 121 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.425 $Y2=0.152
r262 121 123 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r263 121 128 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r264 121 205 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.935 $Y2=0.152
r265 121 196 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.765 $Y2=0.152
r266 121 197 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=7.985 $Y2=0.152
r267 121 187 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r268 121 188 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.125 $Y2=0.152
r269 121 178 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.955 $Y2=0.152
r270 121 179 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.175 $Y2=0.152
r271 121 166 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.005 $Y2=0.152
r272 121 167 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.425 $Y2=0.152
r273 121 154 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=4.255 $Y2=0.152
r274 121 155 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=2.675 $Y2=0.152
r275 121 145 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.505 $Y2=0.152
r276 121 146 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.155 $Y2=0.152
r277 121 136 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.985 $Y2=0.152
r278 121 137 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.295 $Y2=0.152
r279 121 127 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.125 $Y2=0.152
r280 121 128 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r281 9 203 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.575 $X2=8.85 $Y2=0.74
r282 8 194 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.74
r283 7 185 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.575 $X2=7.04 $Y2=0.74
r284 6 176 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.575 $X2=6.09 $Y2=0.865
r285 5 164 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.575 $X2=4.34 $Y2=0.74
r286 4 152 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.575 $X2=2.59 $Y2=0.865
r287 3 143 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.74
r288 2 134 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.74
r289 1 125 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%VDD 1 2 3 4 5 6 7 85 89 93 101 109 113
+ 121 125 133 137 145 147 153 157 172 176
r118 172 176 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=5.397
+ $X2=9.175 $Y2=5.397
r119 161 172 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=5.36 $X2=0.335 $Y2=5.36
r120 157 176 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=5.36 $X2=9.175 $Y2=5.36
r121 155 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=5.397
+ $X2=8.85 $Y2=5.397
r122 155 157 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=8.935 $Y=5.397
+ $X2=9.175 $Y2=5.397
r123 151 170 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.85 $Y=5.245
+ $X2=8.85 $Y2=5.397
r124 151 153 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.85 $Y=5.245
+ $X2=8.85 $Y2=4.225
r125 148 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=5.397
+ $X2=7.83 $Y2=5.397
r126 148 150 21.9153 $w=3.03e-07 $l=5.8e-07 $layer=LI1_cond $X=7.915 $Y=5.397
+ $X2=8.495 $Y2=5.397
r127 147 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=5.397
+ $X2=8.85 $Y2=5.397
r128 147 150 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.765 $Y=5.397
+ $X2=8.495 $Y2=5.397
r129 143 169 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.83 $Y=5.245
+ $X2=7.83 $Y2=5.397
r130 143 145 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.83 $Y=5.245
+ $X2=7.83 $Y2=4.225
r131 140 142 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.455 $Y=5.397
+ $X2=7.135 $Y2=5.397
r132 138 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=5.397
+ $X2=6.09 $Y2=5.397
r133 138 140 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=5.397
+ $X2=6.455 $Y2=5.397
r134 137 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=5.397
+ $X2=7.83 $Y2=5.397
r135 137 142 23.0489 $w=3.03e-07 $l=6.1e-07 $layer=LI1_cond $X=7.745 $Y=5.397
+ $X2=7.135 $Y2=5.397
r136 133 136 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.09 $Y=3.205
+ $X2=6.09 $Y2=4.565
r137 131 167 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=5.245
+ $X2=6.09 $Y2=5.397
r138 131 136 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.09 $Y=5.245
+ $X2=6.09 $Y2=4.565
r139 128 130 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=5.397
+ $X2=5.775 $Y2=5.397
r140 126 166 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=5.397
+ $X2=4.34 $Y2=5.397
r141 126 128 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.425 $Y=5.397
+ $X2=5.095 $Y2=5.397
r142 125 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=5.397
+ $X2=6.09 $Y2=5.397
r143 125 130 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=5.397
+ $X2=5.775 $Y2=5.397
r144 121 124 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.34 $Y=3.545
+ $X2=4.34 $Y2=4.565
r145 119 166 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.34 $Y=5.245
+ $X2=4.34 $Y2=5.397
r146 119 124 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.34 $Y=5.245
+ $X2=4.34 $Y2=4.565
r147 116 118 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=5.397
+ $X2=3.735 $Y2=5.397
r148 114 164 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=5.397
+ $X2=2.59 $Y2=5.397
r149 114 116 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.675 $Y=5.397
+ $X2=3.055 $Y2=5.397
r150 113 166 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=5.397
+ $X2=4.34 $Y2=5.397
r151 113 118 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=4.255 $Y=5.397
+ $X2=3.735 $Y2=5.397
r152 109 112 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.59 $Y=3.545
+ $X2=2.59 $Y2=4.565
r153 107 164 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.59 $Y=5.245
+ $X2=2.59 $Y2=5.397
r154 107 112 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.59 $Y=5.245
+ $X2=2.59 $Y2=4.565
r155 104 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=5.397
+ $X2=2 $Y2=5.397
r156 104 106 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=2.085 $Y=5.397
+ $X2=2.375 $Y2=5.397
r157 103 164 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=5.397
+ $X2=2.59 $Y2=5.397
r158 103 106 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=5.397
+ $X2=2.375 $Y2=5.397
r159 99 163 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2 $Y=5.245 $X2=2
+ $Y2=5.397
r160 99 101 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2 $Y=5.245 $X2=2
+ $Y2=4.225
r161 96 98 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=5.397
+ $X2=1.695 $Y2=5.397
r162 94 161 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r163 94 96 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.015 $Y2=5.397
r164 93 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=5.397
+ $X2=2 $Y2=5.397
r165 93 98 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.915 $Y=5.397
+ $X2=1.695 $Y2=5.397
r166 89 92 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r167 87 161 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r168 87 92 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r169 85 157 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=5.245 $X2=9.175 $Y2=5.33
r170 85 150 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=5.245 $X2=8.495 $Y2=5.33
r171 85 169 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=5.245 $X2=7.815 $Y2=5.33
r172 85 142 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=5.245 $X2=7.135 $Y2=5.33
r173 85 140 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=5.245 $X2=6.455 $Y2=5.33
r174 85 130 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=5.245 $X2=5.775 $Y2=5.33
r175 85 128 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=5.245 $X2=5.095 $Y2=5.33
r176 85 166 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=5.245 $X2=4.415 $Y2=5.33
r177 85 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=5.245 $X2=3.735 $Y2=5.33
r178 85 116 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=5.245 $X2=3.055 $Y2=5.33
r179 85 106 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=5.245 $X2=2.375 $Y2=5.33
r180 85 98 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=5.245 $X2=1.695 $Y2=5.33
r181 85 96 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=5.245 $X2=1.015 $Y2=5.33
r182 85 161 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=5.245 $X2=0.335 $Y2=5.33
r183 7 153 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=3.565 $X2=8.85 $Y2=4.225
r184 6 145 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=3.565 $X2=7.83 $Y2=4.225
r185 5 136 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=5.95
+ $Y=2.825 $X2=6.09 $Y2=4.565
r186 5 133 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=5.95
+ $Y=2.825 $X2=6.09 $Y2=3.205
r187 4 124 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=2.825 $X2=4.34 $Y2=4.565
r188 4 121 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=2.825 $X2=4.34 $Y2=3.545
r189 3 112 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.825 $X2=2.59 $Y2=4.565
r190 3 109 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.825 $X2=2.59 $Y2=3.545
r191 2 101 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=3.565 $X2=2 $Y2=4.225
r192 1 92 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r193 1 89 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%RN 3 5 7 13 15 21
c39 21 0 7.48684e-20 $X=0.325 $Y=3.07
c40 3 0 1.0746e-19 $X=0.475 $Y=0.895
r41 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=3.07
+ $X2=0.325 $Y2=3.07
r42 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=2.045
+ $X2=0.53 $Y2=2.045
r43 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r44 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.21
+ $X2=0.32 $Y2=2.045
r45 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=2.21 $X2=0.32
+ $Y2=3.07
r46 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=2.045 $X2=0.53 $Y2=2.045
r47 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=2.21
+ $X2=0.53 $Y2=2.045
r48 5 7 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=0.475 $Y=2.21
+ $X2=0.475 $Y2=3.825
r49 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.875
+ $X2=0.53 $Y2=2.045
r50 1 3 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.475 $Y=1.875
+ $X2=0.475 $Y2=0.895
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%A_110_115# 1 3 11 15 19 23 27 30 31 35
+ 39 44 45 46 48 58 61 66 67 72
c175 67 0 1.63751e-20 $X=1.375 $Y=1.22
c176 66 0 1.94136e-20 $X=7.665 $Y=1.22
c177 61 0 9.10849e-20 $X=1.23 $Y=1.22
c178 58 0 7.48684e-20 $X=0.87 $Y=2.48
c179 48 0 7.745e-20 $X=7.81 $Y=1.22
r180 67 69 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.375 $Y=1.22
+ $X2=1.23 $Y2=1.22
r181 66 72 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.665 $Y=1.22
+ $X2=7.81 $Y2=1.22
r182 66 67 6.05653 $w=1.7e-07 $l=6.29e-06 $layer=MET1_cond $X=7.665 $Y=1.22
+ $X2=1.375 $Y2=1.22
r183 61 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.22
+ $X2=1.23 $Y2=1.22
r184 61 64 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.23 $Y=1.22
+ $X2=1.23 $Y2=1.37
r185 56 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.87 $Y2=2.48
r186 53 55 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.87 $Y2=1.37
r187 48 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.81 $Y=1.22
+ $X2=7.81 $Y2=1.22
r188 48 51 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.81 $Y=1.22
+ $X2=7.81 $Y2=1.37
r189 46 55 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.37
+ $X2=0.87 $Y2=1.37
r190 45 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.37
+ $X2=1.23 $Y2=1.37
r191 45 46 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.145 $Y=1.37
+ $X2=0.955 $Y2=1.37
r192 44 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.395
+ $X2=0.87 $Y2=2.48
r193 43 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.455
+ $X2=0.87 $Y2=1.37
r194 43 44 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.87 $Y=1.455
+ $X2=0.87 $Y2=2.395
r195 39 41 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r196 37 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.565
+ $X2=0.69 $Y2=2.48
r197 37 39 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.69 $Y=2.565
+ $X2=0.69 $Y2=3.205
r198 33 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.285
+ $X2=0.69 $Y2=1.37
r199 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.69 $Y=1.285
+ $X2=0.69 $Y2=0.865
r200 30 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.81
+ $Y=1.37 $X2=7.81 $Y2=1.37
r201 30 32 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=7.742 $Y=1.37
+ $X2=7.742 $Y2=1.535
r202 30 31 59.5222 $w=4.05e-07 $l=2.65e-07 $layer=POLY_cond $X=7.742 $Y=1.37
+ $X2=7.742 $Y2=1.105
r203 25 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.37 $X2=1.23 $Y2=1.37
r204 25 27 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.23 $Y=1.37
+ $X2=1.425 $Y2=1.37
r205 23 31 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.685 $Y=0.785
+ $X2=7.685 $Y2=1.105
r206 19 32 1363.96 $w=1.5e-07 $l=2.66e-06 $layer=POLY_cond $X=7.615 $Y=4.195
+ $X2=7.615 $Y2=1.535
r207 13 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.535
+ $X2=1.425 $Y2=1.37
r208 13 15 1363.96 $w=1.5e-07 $l=2.66e-06 $layer=POLY_cond $X=1.425 $Y=1.535
+ $X2=1.425 $Y2=4.195
r209 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.205
+ $X2=1.425 $Y2=1.37
r210 9 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.425 $Y=1.205
+ $X2=1.425 $Y2=0.785
r211 3 41 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r212 3 39 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r213 1 35 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%A_342_466# 1 3 11 15 18 22 24 25 26 27
+ 28 30 33 37 44 47
c86 47 0 1.71621e-19 $X=3.457 $Y=1.155
c87 25 0 1.29912e-19 $X=3.28 $Y=1.505
r88 46 47 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.457 $Y=0.985
+ $X2=3.457 $Y2=1.155
r89 42 44 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.94 $Y=2.495
+ $X2=2.11 $Y2=2.495
r90 37 39 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=3.465 $Y=3.205
+ $X2=3.465 $Y2=4.565
r91 35 37 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=3.465 $Y=3.01
+ $X2=3.465 $Y2=3.205
r92 33 46 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.465 $Y=0.865
+ $X2=3.465 $Y2=0.985
r93 30 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=1.42
+ $X2=3.365 $Y2=1.155
r94 27 35 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.295 $Y=2.925
+ $X2=3.465 $Y2=3.01
r95 27 28 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.295 $Y=2.925
+ $X2=2.195 $Y2=2.925
r96 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=1.505
+ $X2=3.365 $Y2=1.42
r97 25 26 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.28 $Y=1.505
+ $X2=2.195 $Y2=1.505
r98 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=2.84
+ $X2=2.195 $Y2=2.925
r99 23 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=2.66
+ $X2=2.11 $Y2=2.495
r100 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.11 $Y=2.66
+ $X2=2.11 $Y2=2.84
r101 22 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=2.33
+ $X2=2.11 $Y2=2.495
r102 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=1.59
+ $X2=2.195 $Y2=1.505
r103 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.11 $Y=1.59
+ $X2=2.11 $Y2=2.33
r104 18 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.495 $X2=1.94 $Y2=2.495
r105 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.495
+ $X2=1.892 $Y2=2.66
r106 18 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.495
+ $X2=1.892 $Y2=2.33
r107 15 19 792.223 $w=1.5e-07 $l=1.545e-06 $layer=POLY_cond $X=1.855 $Y=0.785
+ $X2=1.855 $Y2=2.33
r108 11 20 787.096 $w=1.5e-07 $l=1.535e-06 $layer=POLY_cond $X=1.785 $Y=4.195
+ $X2=1.785 $Y2=2.66
r109 3 39 240 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=3.24
+ $Y=2.825 $X2=3.465 $Y2=4.565
r110 3 37 240 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=2 $X=3.24
+ $Y=2.825 $X2=3.465 $Y2=3.205
r111 1 33 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.575 $X2=3.465 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%D 3 7 10 14 19
c41 19 0 1.41836e-19 $X=2.865 $Y=1.96
c42 10 0 1.12321e-19 $X=2.865 $Y=1.96
r43 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.865 $Y=1.96
+ $X2=2.865 $Y2=1.96
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.96 $X2=2.865 $Y2=1.96
r45 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.96
+ $X2=2.865 $Y2=2.125
r46 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.96
+ $X2=2.865 $Y2=1.795
r47 7 12 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=2.805 $Y=3.825
+ $X2=2.805 $Y2=2.125
r48 3 11 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.805 $Y=0.895
+ $X2=2.805 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%CK 3 7 11 15 19 21 23 26 28 32 36 40 44
+ 47 51 55 57 58 60 66 73 77 78 79 80 87
c219 58 0 6.79641e-20 $X=5.06 $Y=2.33
c220 51 0 1.98654e-19 $X=3.705 $Y=1.59
c221 47 0 1.86602e-19 $X=3.62 $Y=2.33
c222 28 0 1.41836e-19 $X=3.225 $Y=2.505
c223 7 0 1.29912e-19 $X=3.765 $Y=0.895
r224 80 85 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=2.33
+ $X2=5.455 $Y2=2.33
r225 79 87 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.305 $Y=2.33
+ $X2=6.45 $Y2=2.33
r226 79 80 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.305 $Y=2.33
+ $X2=5.6 $Y2=2.33
r227 78 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.37 $Y=2.33
+ $X2=3.225 $Y2=2.33
r228 77 85 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.31 $Y=2.33
+ $X2=5.455 $Y2=2.33
r229 77 78 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.31 $Y=2.33
+ $X2=3.37 $Y2=2.33
r230 73 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=2.33
+ $X2=5.455 $Y2=2.33
r231 73 75 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.455 $Y=2.33
+ $X2=5.455 $Y2=2.505
r232 66 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.225 $Y=2.33
+ $X2=3.225 $Y2=2.33
r233 66 69 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.225 $Y=2.33
+ $X2=3.225 $Y2=2.505
r234 60 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.45 $Y=2.33
+ $X2=6.45 $Y2=2.33
r235 60 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.45 $Y=2.33
+ $X2=6.45 $Y2=2.505
r236 57 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.33
+ $X2=5.455 $Y2=2.33
r237 57 58 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.37 $Y=2.33
+ $X2=5.06 $Y2=2.33
r238 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=2.245
+ $X2=5.06 $Y2=2.33
r239 53 55 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.975 $Y=2.245
+ $X2=4.975 $Y2=1.59
r240 49 51 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.705 $Y=2.245
+ $X2=3.705 $Y2=1.59
r241 48 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.33
+ $X2=3.225 $Y2=2.33
r242 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.33
+ $X2=3.705 $Y2=2.245
r243 47 48 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.62 $Y=2.33
+ $X2=3.31 $Y2=2.33
r244 46 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=2.505 $X2=6.45 $Y2=2.505
r245 43 44 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.332 $Y=1.425
+ $X2=6.332 $Y2=1.575
r246 40 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=2.505 $X2=5.455 $Y2=2.505
r247 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=2.505
+ $X2=5.455 $Y2=2.67
r248 36 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.59 $X2=4.975 $Y2=1.59
r249 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.59
+ $X2=4.975 $Y2=1.425
r250 32 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.59 $X2=3.705 $Y2=1.59
r251 32 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.59
+ $X2=3.705 $Y2=1.425
r252 28 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=2.505 $X2=3.225 $Y2=2.505
r253 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.505
+ $X2=3.225 $Y2=2.67
r254 26 46 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.36 $Y=2.34
+ $X2=6.407 $Y2=2.505
r255 26 44 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.36 $Y=2.34
+ $X2=6.36 $Y2=1.575
r256 21 46 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.305 $Y=2.67
+ $X2=6.407 $Y2=2.505
r257 21 23 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=6.305 $Y=2.67
+ $X2=6.305 $Y2=3.825
r258 19 43 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.305 $Y=0.895
+ $X2=6.305 $Y2=1.425
r259 15 42 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=5.515 $Y=3.825
+ $X2=5.515 $Y2=2.67
r260 11 37 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.915 $Y=0.895
+ $X2=4.915 $Y2=1.425
r261 7 33 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.765 $Y=0.895
+ $X2=3.765 $Y2=1.425
r262 3 30 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=3.165 $Y=3.825
+ $X2=3.165 $Y2=2.67
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%A_217_713# 1 3 11 15 17 18 21 22 27 31
+ 35 37 38 41 47 52 53 54 59
c140 53 0 1.35571e-19 $X=4.06 $Y=1.59
c141 47 0 1.5821e-19 $X=4.295 $Y=2.505
c142 31 0 6.36774e-20 $X=4.555 $Y=3.825
c143 22 0 1.86602e-19 $X=4.2 $Y=2.505
c144 21 0 6.79641e-20 $X=4.48 $Y=2.505
c145 15 0 6.36774e-20 $X=4.125 $Y=3.825
r146 54 56 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.785 $Y=1.59
+ $X2=1.64 $Y2=1.59
r147 53 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.59
+ $X2=4.205 $Y2=1.59
r148 53 54 2.19056 $w=1.7e-07 $l=2.275e-06 $layer=MET1_cond $X=4.06 $Y=1.59
+ $X2=1.785 $Y2=1.59
r149 50 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=1.59
+ $X2=4.205 $Y2=1.59
r150 50 52 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=1.55
+ $X2=4.295 $Y2=1.55
r151 45 52 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.295 $Y=1.675
+ $X2=4.295 $Y2=1.55
r152 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.295 $Y=1.675
+ $X2=4.295 $Y2=2.505
r153 44 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.59
+ $X2=1.64 $Y2=1.59
r154 41 44 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.64 $Y=0.74
+ $X2=1.64 $Y2=1.59
r155 39 44 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.64 $Y=1.715
+ $X2=1.64 $Y2=1.59
r156 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=1.8
+ $X2=1.64 $Y2=1.715
r157 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.555 $Y=1.8
+ $X2=1.295 $Y2=1.8
r158 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.885
+ $X2=1.295 $Y2=1.8
r159 33 35 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=1.21 $Y=1.885
+ $X2=1.21 $Y2=4.225
r160 29 31 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=4.555 $Y=2.64
+ $X2=4.555 $Y2=3.825
r161 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.555 $Y=1.455
+ $X2=4.555 $Y2=0.895
r162 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=2.505 $X2=4.295 $Y2=2.505
r163 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=2.505
+ $X2=4.295 $Y2=2.505
r164 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=2.505
+ $X2=4.555 $Y2=2.64
r165 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=2.505
+ $X2=4.295 $Y2=2.505
r166 20 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.59 $X2=4.295 $Y2=1.59
r167 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=1.59
+ $X2=4.295 $Y2=1.59
r168 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=1.59
+ $X2=4.555 $Y2=1.455
r169 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=1.59
+ $X2=4.295 $Y2=1.59
r170 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=2.64
+ $X2=4.2 $Y2=2.505
r171 13 15 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=4.125 $Y=2.64
+ $X2=4.125 $Y2=3.825
r172 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=1.455
+ $X2=4.2 $Y2=1.59
r173 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.125 $Y=1.455
+ $X2=4.125 $Y2=0.895
r174 3 35 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=3.565 $X2=1.21 $Y2=4.225
r175 1 41 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%A_618_89# 1 3 11 14 15 16 19 21 25 27 30
+ 33 37 39 40 42 45 51 54 57 62 63 66 70
c187 37 0 2.18068e-19 $X=3.285 $Y=1.5
c188 19 0 1.12321e-19 $X=3.765 $Y=3.825
r189 68 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=2.925
+ $X2=6.795 $Y2=2.925
r190 64 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=1.93
+ $X2=6.795 $Y2=1.93
r191 62 70 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.84
+ $X2=6.795 $Y2=2.925
r192 61 66 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.015
+ $X2=6.795 $Y2=1.93
r193 61 62 50.8333 $w=1.78e-07 $l=8.25e-07 $layer=LI1_cond $X=6.795 $Y=2.015
+ $X2=6.795 $Y2=2.84
r194 57 59 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.52 $Y=3.205
+ $X2=6.52 $Y2=4.565
r195 55 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=3.01
+ $X2=6.52 $Y2=2.925
r196 55 57 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.52 $Y=3.01
+ $X2=6.52 $Y2=3.205
r197 54 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.845
+ $X2=6.52 $Y2=1.93
r198 53 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.675
+ $X2=6.52 $Y2=1.59
r199 53 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=1.675
+ $X2=6.52 $Y2=1.845
r200 49 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.505
+ $X2=6.52 $Y2=1.59
r201 49 51 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.52 $Y=1.505
+ $X2=6.52 $Y2=0.865
r202 45 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=1.59
+ $X2=6.52 $Y2=1.59
r203 45 47 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.435 $Y=1.59
+ $X2=5.455 $Y2=1.59
r204 42 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.59 $X2=5.455 $Y2=1.59
r205 42 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.59
+ $X2=5.455 $Y2=1.755
r206 42 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.59
+ $X2=5.455 $Y2=1.425
r207 35 37 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.165 $Y=1.5
+ $X2=3.285 $Y2=1.5
r208 33 43 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.515 $Y=0.895
+ $X2=5.515 $Y2=1.425
r209 30 44 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.395 $Y=1.965
+ $X2=5.395 $Y2=1.755
r210 28 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.99 $Y=2.04
+ $X2=4.915 $Y2=2.04
r211 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.32 $Y=2.04
+ $X2=5.395 $Y2=1.965
r212 27 28 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.32 $Y=2.04
+ $X2=4.99 $Y2=2.04
r213 23 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.915 $Y=2.115
+ $X2=4.915 $Y2=2.04
r214 23 25 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=4.915 $Y=2.115
+ $X2=4.915 $Y2=3.825
r215 22 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.04
+ $X2=3.765 $Y2=2.04
r216 21 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=2.04
+ $X2=4.915 $Y2=2.04
r217 21 22 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.84 $Y=2.04 $X2=3.84
+ $Y2=2.04
r218 17 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=2.115
+ $X2=3.765 $Y2=2.04
r219 17 19 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=3.765 $Y=2.115
+ $X2=3.765 $Y2=3.825
r220 15 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=2.04
+ $X2=3.765 $Y2=2.04
r221 15 16 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.69 $Y=2.04
+ $X2=3.36 $Y2=2.04
r222 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.285 $Y=1.965
+ $X2=3.36 $Y2=2.04
r223 13 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.575
+ $X2=3.285 $Y2=1.5
r224 13 14 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.285 $Y=1.575
+ $X2=3.285 $Y2=1.965
r225 9 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.425
+ $X2=3.165 $Y2=1.5
r226 9 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.165 $Y=1.425
+ $X2=3.165 $Y2=0.895
r227 3 59 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=2.825 $X2=6.52 $Y2=4.565
r228 3 57 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=2.825 $X2=6.52 $Y2=3.205
r229 1 51 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%A_1160_89# 1 3 11 15 23 27 30 34 35 38
+ 39 40 42 48 50 51 54 57 60 63 64 65 70
c162 39 0 8.77106e-20 $X=8.61 $Y=2.595
c163 38 0 7.745e-20 $X=8.61 $Y=1.54
c164 34 0 2.20654e-19 $X=8.52 $Y=1.93
r165 65 67 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=1.93
+ $X2=5.935 $Y2=1.93
r166 64 70 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.375 $Y=1.93
+ $X2=8.52 $Y2=1.93
r167 64 65 2.20982 $w=1.7e-07 $l=2.295e-06 $layer=MET1_cond $X=8.375 $Y=1.93
+ $X2=6.08 $Y2=1.93
r168 60 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.52 $Y=1.93
+ $X2=8.52 $Y2=1.93
r169 58 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=1.93
+ $X2=7.47 $Y2=1.93
r170 58 60 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.555 $Y=1.93
+ $X2=8.52 $Y2=1.93
r171 56 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=2.015
+ $X2=7.47 $Y2=1.93
r172 56 57 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.47 $Y=2.015
+ $X2=7.47 $Y2=3.435
r173 52 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.845
+ $X2=7.47 $Y2=1.93
r174 52 54 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=7.47 $Y=1.845
+ $X2=7.47 $Y2=0.74
r175 50 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=3.52
+ $X2=7.47 $Y2=3.435
r176 50 51 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.385 $Y=3.52
+ $X2=7.125 $Y2=3.52
r177 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=3.605
+ $X2=7.125 $Y2=3.52
r178 46 48 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.04 $Y=3.605
+ $X2=7.04 $Y2=4.225
r179 42 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.935 $Y=1.93
+ $X2=5.935 $Y2=1.93
r180 39 40 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=2.595
+ $X2=8.61 $Y2=2.745
r181 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=1.39 $X2=8.61
+ $Y2=1.54
r182 36 39 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=8.585 $Y=2.095
+ $X2=8.585 $Y2=2.595
r183 35 38 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.585 $Y=1.765
+ $X2=8.585 $Y2=1.54
r184 34 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.52
+ $Y=1.93 $X2=8.52 $Y2=1.93
r185 34 36 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.93
+ $X2=8.522 $Y2=2.095
r186 34 35 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.93
+ $X2=8.522 $Y2=1.765
r187 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.935
+ $Y=1.93 $X2=5.935 $Y2=1.93
r188 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=1.93
+ $X2=5.935 $Y2=2.095
r189 30 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=1.93
+ $X2=5.935 $Y2=1.765
r190 27 40 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=8.635 $Y=4.195
+ $X2=8.635 $Y2=2.745
r191 23 37 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=8.635 $Y=0.785
+ $X2=8.635 $Y2=1.39
r192 15 32 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=5.875 $Y=3.825
+ $X2=5.875 $Y2=2.095
r193 11 31 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.875 $Y=0.895
+ $X2=5.875 $Y2=1.765
r194 3 48 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=3.565 $X2=7.04 $Y2=4.225
r195 1 54 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.575 $X2=7.47 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%A_998_115# 1 3 11 13 15 22 23 24 25 26
+ 29 33 38 42 43 48
c130 43 0 1.5821e-19 $X=4.78 $Y=1.59
c131 23 0 1.67294e-19 $X=5.045 $Y=1.17
c132 22 0 1.57671e-19 $X=4.635 $Y=1.59
r133 43 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.78 $Y=1.59
+ $X2=4.635 $Y2=1.59
r134 42 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=1.59
+ $X2=7.13 $Y2=1.59
r135 42 43 2.12316 $w=1.7e-07 $l=2.205e-06 $layer=MET1_cond $X=6.985 $Y=1.59
+ $X2=4.78 $Y2=1.59
r136 38 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=1.59
+ $X2=7.13 $Y2=1.59
r137 33 35 34.5733 $w=3.38e-07 $l=1.02e-06 $layer=LI1_cond $X=5.215 $Y=3.545
+ $X2=5.215 $Y2=4.565
r138 31 33 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=5.215 $Y=3.01
+ $X2=5.215 $Y2=3.545
r139 27 29 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=5.215 $Y=1.085
+ $X2=5.215 $Y2=0.865
r140 25 31 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=2.925
+ $X2=5.215 $Y2=3.01
r141 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=2.925
+ $X2=4.72 $Y2=2.925
r142 23 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=1.17
+ $X2=5.215 $Y2=1.085
r143 23 24 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=1.17
+ $X2=4.72 $Y2=1.17
r144 22 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.59
+ $X2=4.635 $Y2=1.59
r145 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=2.84
+ $X2=4.72 $Y2=2.925
r146 20 22 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.635 $Y=2.84
+ $X2=4.635 $Y2=1.59
r147 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=1.255
+ $X2=4.72 $Y2=1.17
r148 19 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.635 $Y=1.255
+ $X2=4.635 $Y2=1.59
r149 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.59 $X2=7.13 $Y2=1.59
r150 13 18 38.6212 $w=3.33e-07 $l=2.06325e-07 $layer=POLY_cond $X=7.255 $Y=1.755
+ $X2=7.162 $Y2=1.59
r151 13 15 1251.15 $w=1.5e-07 $l=2.44e-06 $layer=POLY_cond $X=7.255 $Y=1.755
+ $X2=7.255 $Y2=4.195
r152 9 18 39.3449 $w=3.33e-07 $l=2.11447e-07 $layer=POLY_cond $X=7.255 $Y=1.42
+ $X2=7.162 $Y2=1.59
r153 9 11 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.255 $Y=1.42
+ $X2=7.255 $Y2=0.785
r154 3 35 300 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.825 $X2=5.215 $Y2=4.565
r155 3 33 300 $w=1.7e-07 $l=8.24864e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.825 $X2=5.215 $Y2=3.545
r156 1 29 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.575 $X2=5.215 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c85 42 0 8.77106e-20 $X=8.425 $Y=2.7
c86 33 0 9.99996e-20 $X=8.92 $Y=2.505
c87 31 0 1.20654e-19 $X=8.92 $Y=1.59
r88 40 42 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=8.42 $Y=2.7
+ $X2=8.425 $Y2=2.7
r89 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.005 $Y=2.42
+ $X2=9.005 $Y2=2.135
r90 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.005 $Y=1.675
+ $X2=9.005 $Y2=2.135
r91 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=2.505
+ $X2=9.005 $Y2=2.42
r92 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=2.505
+ $X2=8.505 $Y2=2.505
r93 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=1.59
+ $X2=9.005 $Y2=1.675
r94 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=1.59
+ $X2=8.505 $Y2=1.59
r95 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.42 $Y=2.7 $X2=8.42
+ $Y2=2.7
r96 27 29 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=8.42 $Y=2.7
+ $X2=8.42 $Y2=4.225
r97 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=2.59
+ $X2=8.505 $Y2=2.505
r98 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.42 $Y=2.59
+ $X2=8.42 $Y2=2.7
r99 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=1.505
+ $X2=8.505 $Y2=1.59
r100 21 23 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=8.42 $Y=1.505
+ $X2=8.42 $Y2=0.74
r101 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=2.135 $X2=9.005 $Y2=2.135
r102 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=2.135
+ $X2=9.005 $Y2=2.3
r103 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=2.135
+ $X2=9.005 $Y2=1.97
r104 15 20 971.691 $w=1.5e-07 $l=1.895e-06 $layer=POLY_cond $X=9.065 $Y=4.195
+ $X2=9.065 $Y2=2.3
r105 11 19 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=9.065 $Y=0.785
+ $X2=9.065 $Y2=1.97
r106 3 29 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=3.565 $X2=8.42 $Y2=4.225
r107 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.575 $X2=8.42 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__DFFR_L%Q 1 3 11 15 18 21 25 28
r22 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=3.027
+ $X2=9.395 $Y2=3.027
r23 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=3.07
+ $X2=9.275 $Y2=3.07
r24 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=9.275 $Y=3.027
+ $X2=9.28 $Y2=3.027
r25 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=1.255
+ $X2=9.395 $Y2=1.255
r26 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.395 $Y=2.9
+ $X2=9.395 $Y2=3.027
r27 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.34
+ $X2=9.395 $Y2=1.255
r28 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=9.395 $Y=1.34
+ $X2=9.395 $Y2=2.9
r29 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.28 $Y=3.155
+ $X2=9.28 $Y2=3.027
r30 13 15 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=9.28 $Y=3.155
+ $X2=9.28 $Y2=4.225
r31 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=1.17 $X2=9.28
+ $Y2=1.255
r32 9 11 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.28 $Y=1.17 $X2=9.28
+ $Y2=0.74
r33 3 15 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=3.565 $X2=9.28 $Y2=4.225
r34 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.575 $X2=9.28 $Y2=0.74
.ends

