* File: sky130_osu_sc_12T_hs__inv_8.pxi.spice
* Created: Fri Nov 12 15:11:19 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__INV_8%GND N_GND_M1001_d N_GND_M1002_d N_GND_M1011_d
+ N_GND_M1013_d N_GND_M1015_d N_GND_M1001_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p
+ N_GND_c_17_p N_GND_c_23_p N_GND_c_30_p N_GND_c_37_p N_GND_c_44_p N_GND_c_50_p
+ GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_HS__INV_8%GND
x_PM_SKY130_OSU_SC_12T_HS__INV_8%VDD N_VDD_M1000_s N_VDD_M1003_s N_VDD_M1005_s
+ N_VDD_M1008_s N_VDD_M1010_s N_VDD_M1000_b N_VDD_c_118_p N_VDD_c_119_p
+ N_VDD_c_124_p N_VDD_c_130_p N_VDD_c_135_p N_VDD_c_141_p N_VDD_c_146_p
+ N_VDD_c_152_p N_VDD_c_157_p VDD N_VDD_c_120_p
+ PM_SKY130_OSU_SC_12T_HS__INV_8%VDD
x_PM_SKY130_OSU_SC_12T_HS__INV_8%A N_A_c_194_n N_A_M1001_g N_A_c_198_n
+ N_A_c_264_n N_A_M1000_g N_A_c_199_n N_A_c_200_n N_A_c_201_n N_A_M1002_g
+ N_A_c_269_n N_A_M1003_g N_A_c_205_n N_A_c_207_n N_A_c_208_n N_A_M1006_g
+ N_A_c_275_n N_A_M1004_g N_A_c_212_n N_A_c_213_n N_A_c_214_n N_A_M1011_g
+ N_A_c_280_n N_A_M1005_g N_A_c_218_n N_A_c_220_n N_A_c_221_n N_A_M1012_g
+ N_A_c_225_n N_A_c_286_n N_A_M1007_g N_A_c_226_n N_A_c_227_n N_A_c_228_n
+ N_A_M1013_g N_A_c_291_n N_A_M1008_g N_A_c_232_n N_A_c_234_n N_A_c_235_n
+ N_A_M1014_g N_A_c_297_n N_A_M1009_g N_A_c_239_n N_A_c_240_n N_A_c_241_n
+ N_A_M1015_g N_A_c_302_n N_A_M1010_g N_A_c_245_n N_A_c_246_n N_A_c_247_n
+ N_A_c_248_n N_A_c_249_n N_A_c_250_n N_A_c_251_n N_A_c_252_n N_A_c_253_n
+ N_A_c_254_n N_A_c_255_n N_A_c_256_n N_A_c_257_n N_A_c_258_n N_A_c_259_n
+ N_A_c_260_n N_A_c_261_n N_A_c_262_n N_A_c_263_n A
+ PM_SKY130_OSU_SC_12T_HS__INV_8%A
x_PM_SKY130_OSU_SC_12T_HS__INV_8%Y N_Y_M1001_s N_Y_M1006_s N_Y_M1012_s
+ N_Y_M1014_s N_Y_M1000_d N_Y_M1004_d N_Y_M1007_d N_Y_M1009_d N_Y_c_428_n
+ N_Y_c_474_n N_Y_c_432_n N_Y_c_477_n N_Y_c_437_n N_Y_c_480_n N_Y_c_442_n
+ N_Y_c_483_n N_Y_c_446_n N_Y_c_486_n Y N_Y_c_450_n N_Y_c_487_n N_Y_c_454_n
+ N_Y_c_455_n N_Y_c_459_n N_Y_c_489_n N_Y_c_491_n N_Y_c_462_n N_Y_c_463_n
+ N_Y_c_467_n N_Y_c_492_n N_Y_c_494_n N_Y_c_470_n N_Y_c_473_n
+ PM_SKY130_OSU_SC_12T_HS__INV_8%Y
cc_1 N_GND_M1001_b N_A_c_194_n 0.018528f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.22
cc_2 N_GND_c_2_p N_A_c_194_n 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=1.22
cc_3 N_GND_c_3_p N_A_c_194_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.22
cc_4 N_GND_c_4_p N_A_c_194_n 0.00468827f $X=3.06 $Y=0.19 $X2=0.475 $Y2=1.22
cc_5 N_GND_M1001_b N_A_c_198_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.33
cc_6 N_GND_M1001_b N_A_c_199_n 0.01476f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.295
cc_7 N_GND_M1001_b N_A_c_200_n 0.00981662f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.405
cc_8 N_GND_M1001_b N_A_c_201_n 0.0152079f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.22
cc_9 N_GND_c_3_p N_A_c_201_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.22
cc_10 N_GND_c_10_p N_A_c_201_n 0.00311745f $X=1.12 $Y=0.755 $X2=0.905 $Y2=1.22
cc_11 N_GND_c_4_p N_A_c_201_n 0.00468827f $X=3.06 $Y=0.19 $X2=0.905 $Y2=1.22
cc_12 N_GND_M1001_b N_A_c_205_n 0.0213783f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.295
cc_13 N_GND_c_10_p N_A_c_205_n 0.00283047f $X=1.12 $Y=0.755 $X2=1.26 $Y2=1.295
cc_14 N_GND_M1001_b N_A_c_207_n 0.0173499f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.405
cc_15 N_GND_M1001_b N_A_c_208_n 0.0152079f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.22
cc_16 N_GND_c_10_p N_A_c_208_n 0.00311745f $X=1.12 $Y=0.755 $X2=1.335 $Y2=1.22
cc_17 N_GND_c_17_p N_A_c_208_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.335 $Y2=1.22
cc_18 N_GND_c_4_p N_A_c_208_n 0.00468827f $X=3.06 $Y=0.19 $X2=1.335 $Y2=1.22
cc_19 N_GND_M1001_b N_A_c_212_n 0.0195339f $X=-0.045 $Y=0 $X2=1.69 $Y2=1.295
cc_20 N_GND_M1001_b N_A_c_213_n 0.0145324f $X=-0.045 $Y=0 $X2=1.69 $Y2=2.405
cc_21 N_GND_M1001_b N_A_c_214_n 0.0152079f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.22
cc_22 N_GND_c_17_p N_A_c_214_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.765 $Y2=1.22
cc_23 N_GND_c_23_p N_A_c_214_n 0.00311745f $X=1.98 $Y=0.755 $X2=1.765 $Y2=1.22
cc_24 N_GND_c_4_p N_A_c_214_n 0.00468827f $X=3.06 $Y=0.19 $X2=1.765 $Y2=1.22
cc_25 N_GND_M1001_b N_A_c_218_n 0.0164591f $X=-0.045 $Y=0 $X2=2.12 $Y2=1.295
cc_26 N_GND_c_23_p N_A_c_218_n 0.00283047f $X=1.98 $Y=0.755 $X2=2.12 $Y2=1.295
cc_27 N_GND_M1001_b N_A_c_220_n 0.0124307f $X=-0.045 $Y=0 $X2=2.12 $Y2=2.405
cc_28 N_GND_M1001_b N_A_c_221_n 0.0152079f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.22
cc_29 N_GND_c_23_p N_A_c_221_n 0.00311745f $X=1.98 $Y=0.755 $X2=2.195 $Y2=1.22
cc_30 N_GND_c_30_p N_A_c_221_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.195 $Y2=1.22
cc_31 N_GND_c_4_p N_A_c_221_n 0.00468827f $X=3.06 $Y=0.19 $X2=2.195 $Y2=1.22
cc_32 N_GND_M1001_b N_A_c_225_n 0.0685082f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.33
cc_33 N_GND_M1001_b N_A_c_226_n 0.0195339f $X=-0.045 $Y=0 $X2=2.55 $Y2=1.295
cc_34 N_GND_M1001_b N_A_c_227_n 0.0145324f $X=-0.045 $Y=0 $X2=2.55 $Y2=2.405
cc_35 N_GND_M1001_b N_A_c_228_n 0.0152079f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.22
cc_36 N_GND_c_30_p N_A_c_228_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.625 $Y2=1.22
cc_37 N_GND_c_37_p N_A_c_228_n 0.00311745f $X=2.84 $Y=0.755 $X2=2.625 $Y2=1.22
cc_38 N_GND_c_4_p N_A_c_228_n 0.00468827f $X=3.06 $Y=0.19 $X2=2.625 $Y2=1.22
cc_39 N_GND_M1001_b N_A_c_232_n 0.0213783f $X=-0.045 $Y=0 $X2=2.98 $Y2=1.295
cc_40 N_GND_c_37_p N_A_c_232_n 0.00283047f $X=2.84 $Y=0.755 $X2=2.98 $Y2=1.295
cc_41 N_GND_M1001_b N_A_c_234_n 0.0173499f $X=-0.045 $Y=0 $X2=2.98 $Y2=2.405
cc_42 N_GND_M1001_b N_A_c_235_n 0.0152079f $X=-0.045 $Y=0 $X2=3.055 $Y2=1.22
cc_43 N_GND_c_37_p N_A_c_235_n 0.00311745f $X=2.84 $Y=0.755 $X2=3.055 $Y2=1.22
cc_44 N_GND_c_44_p N_A_c_235_n 0.00606474f $X=3.615 $Y=0.152 $X2=3.055 $Y2=1.22
cc_45 N_GND_c_4_p N_A_c_235_n 0.00468827f $X=3.06 $Y=0.19 $X2=3.055 $Y2=1.22
cc_46 N_GND_M1001_b N_A_c_239_n 0.0385034f $X=-0.045 $Y=0 $X2=3.41 $Y2=1.295
cc_47 N_GND_M1001_b N_A_c_240_n 0.0295863f $X=-0.045 $Y=0 $X2=3.41 $Y2=2.405
cc_48 N_GND_M1001_b N_A_c_241_n 0.018528f $X=-0.045 $Y=0 $X2=3.485 $Y2=1.22
cc_49 N_GND_c_44_p N_A_c_241_n 0.00606474f $X=3.615 $Y=0.152 $X2=3.485 $Y2=1.22
cc_50 N_GND_c_50_p N_A_c_241_n 0.00502587f $X=3.7 $Y=0.755 $X2=3.485 $Y2=1.22
cc_51 N_GND_c_4_p N_A_c_241_n 0.00468827f $X=3.06 $Y=0.19 $X2=3.485 $Y2=1.22
cc_52 N_GND_M1001_b N_A_c_245_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.295
cc_53 N_GND_M1001_b N_A_c_246_n 0.0382476f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_54 N_GND_M1001_b N_A_c_247_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.66
cc_55 N_GND_M1001_b N_A_c_248_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.405
cc_56 N_GND_M1001_b N_A_c_249_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.295
cc_57 N_GND_M1001_b N_A_c_250_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.405
cc_58 N_GND_M1001_b N_A_c_251_n 0.0106787f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.295
cc_59 N_GND_M1001_b N_A_c_252_n 0.00980309f $X=-0.045 $Y=0 $X2=1.335 $Y2=2.405
cc_60 N_GND_M1001_b N_A_c_253_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.295
cc_61 N_GND_M1001_b N_A_c_254_n 0.00980309f $X=-0.045 $Y=0 $X2=1.765 $Y2=2.405
cc_62 N_GND_M1001_b N_A_c_255_n 0.0023879f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.295
cc_63 N_GND_M1001_b N_A_c_256_n 0.00151234f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.405
cc_64 N_GND_M1001_b N_A_c_257_n 0.0106787f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.295
cc_65 N_GND_M1001_b N_A_c_258_n 0.00980309f $X=-0.045 $Y=0 $X2=2.625 $Y2=2.405
cc_66 N_GND_M1001_b N_A_c_259_n 0.0106787f $X=-0.045 $Y=0 $X2=3.055 $Y2=1.295
cc_67 N_GND_M1001_b N_A_c_260_n 0.00980309f $X=-0.045 $Y=0 $X2=3.055 $Y2=2.405
cc_68 N_GND_M1001_b N_A_c_261_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.85
cc_69 N_GND_M1001_b N_A_c_262_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.825
cc_70 N_GND_M1001_b N_A_c_263_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_71 N_GND_M1001_b N_Y_c_428_n 0.00154299f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.755
cc_72 N_GND_c_3_p N_Y_c_428_n 0.00740081f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.755
cc_73 N_GND_c_10_p N_Y_c_428_n 8.14297e-19 $X=1.12 $Y=0.755 $X2=0.69 $Y2=0.755
cc_74 N_GND_c_4_p N_Y_c_428_n 0.0047139f $X=3.06 $Y=0.19 $X2=0.69 $Y2=0.755
cc_75 N_GND_M1001_b N_Y_c_432_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_76 N_GND_c_10_p N_Y_c_432_n 8.14297e-19 $X=1.12 $Y=0.755 $X2=1.55 $Y2=0.755
cc_77 N_GND_c_17_p N_Y_c_432_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_78 N_GND_c_23_p N_Y_c_432_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=0.755
cc_79 N_GND_c_4_p N_Y_c_432_n 0.0047139f $X=3.06 $Y=0.19 $X2=1.55 $Y2=0.755
cc_80 N_GND_M1001_b N_Y_c_437_n 0.00154299f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.755
cc_81 N_GND_c_23_p N_Y_c_437_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=2.41 $Y2=0.755
cc_82 N_GND_c_30_p N_Y_c_437_n 0.00718527f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.755
cc_83 N_GND_c_37_p N_Y_c_437_n 8.14297e-19 $X=2.84 $Y=0.755 $X2=2.41 $Y2=0.755
cc_84 N_GND_c_4_p N_Y_c_437_n 0.0047139f $X=3.06 $Y=0.19 $X2=2.41 $Y2=0.755
cc_85 N_GND_M1001_b N_Y_c_442_n 0.00154299f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.755
cc_86 N_GND_c_37_p N_Y_c_442_n 8.14297e-19 $X=2.84 $Y=0.755 $X2=3.27 $Y2=0.755
cc_87 N_GND_c_44_p N_Y_c_442_n 0.00729945f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.755
cc_88 N_GND_c_4_p N_Y_c_442_n 0.0047139f $X=3.06 $Y=0.19 $X2=3.27 $Y2=0.755
cc_89 N_GND_c_2_p N_Y_c_446_n 0.00134236f $X=0.26 $Y=0.755 $X2=0.69 $Y2=1.115
cc_90 N_GND_c_3_p N_Y_c_446_n 0.00245319f $X=1.035 $Y=0.152 $X2=0.69 $Y2=1.115
cc_91 N_GND_c_10_p N_Y_c_446_n 7.53951e-19 $X=1.12 $Y=0.755 $X2=0.69 $Y2=1.115
cc_92 N_GND_M1001_b Y 0.0453816f $X=-0.045 $Y=0 $X2=0.76 $Y2=1.72
cc_93 N_GND_M1002_d N_Y_c_450_n 0.0100144f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1
cc_94 N_GND_c_3_p N_Y_c_450_n 0.0028844f $X=1.035 $Y=0.152 $X2=1.405 $Y2=1
cc_95 N_GND_c_10_p N_Y_c_450_n 0.0142303f $X=1.12 $Y=0.755 $X2=1.405 $Y2=1
cc_96 N_GND_c_17_p N_Y_c_450_n 0.0028844f $X=1.895 $Y=0.152 $X2=1.405 $Y2=1
cc_97 N_GND_M1001_b N_Y_c_454_n 0.0589286f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.365
cc_98 N_GND_M1011_d N_Y_c_455_n 0.0100144f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1
cc_99 N_GND_c_17_p N_Y_c_455_n 0.0028844f $X=1.895 $Y=0.152 $X2=2.265 $Y2=1
cc_100 N_GND_c_23_p N_Y_c_455_n 0.0142303f $X=1.98 $Y=0.755 $X2=2.265 $Y2=1
cc_101 N_GND_c_30_p N_Y_c_455_n 0.0028844f $X=2.755 $Y=0.152 $X2=2.265 $Y2=1
cc_102 N_GND_c_10_p N_Y_c_459_n 7.53951e-19 $X=1.12 $Y=0.755 $X2=1.695 $Y2=1
cc_103 N_GND_c_17_p N_Y_c_459_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.695 $Y2=1
cc_104 N_GND_c_23_p N_Y_c_459_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=1.695 $Y2=1
cc_105 N_GND_M1001_b N_Y_c_462_n 0.0577603f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.365
cc_106 N_GND_M1013_d N_Y_c_463_n 0.0100144f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1
cc_107 N_GND_c_30_p N_Y_c_463_n 0.0028844f $X=2.755 $Y=0.152 $X2=3.125 $Y2=1
cc_108 N_GND_c_37_p N_Y_c_463_n 0.0142303f $X=2.84 $Y=0.755 $X2=3.125 $Y2=1
cc_109 N_GND_c_44_p N_Y_c_463_n 0.0028844f $X=3.615 $Y=0.152 $X2=3.125 $Y2=1
cc_110 N_GND_c_23_p N_Y_c_467_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=2.555 $Y2=1
cc_111 N_GND_c_30_p N_Y_c_467_n 0.00245319f $X=2.755 $Y=0.152 $X2=2.555 $Y2=1
cc_112 N_GND_c_37_p N_Y_c_467_n 7.53951e-19 $X=2.84 $Y=0.755 $X2=2.555 $Y2=1
cc_113 N_GND_c_37_p N_Y_c_470_n 7.53951e-19 $X=2.84 $Y=0.755 $X2=3.27 $Y2=1.115
cc_114 N_GND_c_44_p N_Y_c_470_n 0.00245319f $X=3.615 $Y=0.152 $X2=3.27 $Y2=1.115
cc_115 N_GND_c_50_p N_Y_c_470_n 0.00134236f $X=3.7 $Y=0.755 $X2=3.27 $Y2=1.115
cc_116 N_GND_M1001_b N_Y_c_473_n 0.07516f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.365
cc_117 N_VDD_M1000_b N_A_c_264_n 0.0181616f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.48
cc_118 N_VDD_c_118_p N_A_c_264_n 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=2.48
cc_119 N_VDD_c_119_p N_A_c_264_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.475
+ $Y2=2.48
cc_120 N_VDD_c_120_p N_A_c_264_n 0.00468827f $X=3.06 $Y=4.25 $X2=0.475 $Y2=2.48
cc_121 N_VDD_M1000_b N_A_c_200_n 0.00448664f $X=-0.045 $Y=2.425 $X2=0.83
+ $Y2=2.405
cc_122 N_VDD_M1000_b N_A_c_269_n 0.0159283f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.48
cc_123 N_VDD_c_119_p N_A_c_269_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.905
+ $Y2=2.48
cc_124 N_VDD_c_124_p N_A_c_269_n 0.00337744f $X=1.12 $Y=2.955 $X2=0.905 $Y2=2.48
cc_125 N_VDD_c_120_p N_A_c_269_n 0.00468827f $X=3.06 $Y=4.25 $X2=0.905 $Y2=2.48
cc_126 N_VDD_M1000_b N_A_c_207_n 0.00500158f $X=-0.045 $Y=2.425 $X2=1.26
+ $Y2=2.405
cc_127 N_VDD_c_124_p N_A_c_207_n 0.00341318f $X=1.12 $Y=2.955 $X2=1.26 $Y2=2.405
cc_128 N_VDD_M1000_b N_A_c_275_n 0.0159283f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.48
cc_129 N_VDD_c_124_p N_A_c_275_n 0.00337744f $X=1.12 $Y=2.955 $X2=1.335 $Y2=2.48
cc_130 N_VDD_c_130_p N_A_c_275_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335
+ $Y2=2.48
cc_131 N_VDD_c_120_p N_A_c_275_n 0.00468827f $X=3.06 $Y=4.25 $X2=1.335 $Y2=2.48
cc_132 N_VDD_M1000_b N_A_c_213_n 0.00448664f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_133 N_VDD_M1000_b N_A_c_280_n 0.0159283f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.48
cc_134 N_VDD_c_130_p N_A_c_280_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.765
+ $Y2=2.48
cc_135 N_VDD_c_135_p N_A_c_280_n 0.00337744f $X=1.98 $Y=2.955 $X2=1.765 $Y2=2.48
cc_136 N_VDD_c_120_p N_A_c_280_n 0.00468827f $X=3.06 $Y=4.25 $X2=1.765 $Y2=2.48
cc_137 N_VDD_M1000_b N_A_c_220_n 0.00500158f $X=-0.045 $Y=2.425 $X2=2.12
+ $Y2=2.405
cc_138 N_VDD_c_135_p N_A_c_220_n 0.00341318f $X=1.98 $Y=2.955 $X2=2.12 $Y2=2.405
cc_139 N_VDD_M1000_b N_A_c_286_n 0.0159283f $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.48
cc_140 N_VDD_c_135_p N_A_c_286_n 0.00337744f $X=1.98 $Y=2.955 $X2=2.195 $Y2=2.48
cc_141 N_VDD_c_141_p N_A_c_286_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.195
+ $Y2=2.48
cc_142 N_VDD_c_120_p N_A_c_286_n 0.00468827f $X=3.06 $Y=4.25 $X2=2.195 $Y2=2.48
cc_143 N_VDD_M1000_b N_A_c_227_n 0.00448664f $X=-0.045 $Y=2.425 $X2=2.55
+ $Y2=2.405
cc_144 N_VDD_M1000_b N_A_c_291_n 0.0159283f $X=-0.045 $Y=2.425 $X2=2.625
+ $Y2=2.48
cc_145 N_VDD_c_141_p N_A_c_291_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.625
+ $Y2=2.48
cc_146 N_VDD_c_146_p N_A_c_291_n 0.00337744f $X=2.84 $Y=2.955 $X2=2.625 $Y2=2.48
cc_147 N_VDD_c_120_p N_A_c_291_n 0.00468827f $X=3.06 $Y=4.25 $X2=2.625 $Y2=2.48
cc_148 N_VDD_M1000_b N_A_c_234_n 0.00500158f $X=-0.045 $Y=2.425 $X2=2.98
+ $Y2=2.405
cc_149 N_VDD_c_146_p N_A_c_234_n 0.00341318f $X=2.84 $Y=2.955 $X2=2.98 $Y2=2.405
cc_150 N_VDD_M1000_b N_A_c_297_n 0.0159283f $X=-0.045 $Y=2.425 $X2=3.055
+ $Y2=2.48
cc_151 N_VDD_c_146_p N_A_c_297_n 0.00337744f $X=2.84 $Y=2.955 $X2=3.055 $Y2=2.48
cc_152 N_VDD_c_152_p N_A_c_297_n 0.00606474f $X=3.615 $Y=4.287 $X2=3.055
+ $Y2=2.48
cc_153 N_VDD_c_120_p N_A_c_297_n 0.00468827f $X=3.06 $Y=4.25 $X2=3.055 $Y2=2.48
cc_154 N_VDD_M1000_b N_A_c_240_n 0.00840215f $X=-0.045 $Y=2.425 $X2=3.41
+ $Y2=2.405
cc_155 N_VDD_M1000_b N_A_c_302_n 0.0204783f $X=-0.045 $Y=2.425 $X2=3.485
+ $Y2=2.48
cc_156 N_VDD_c_152_p N_A_c_302_n 0.00606474f $X=3.615 $Y=4.287 $X2=3.485
+ $Y2=2.48
cc_157 N_VDD_c_157_p N_A_c_302_n 0.00636672f $X=3.7 $Y=2.955 $X2=3.485 $Y2=2.48
cc_158 N_VDD_c_120_p N_A_c_302_n 0.00468827f $X=3.06 $Y=4.25 $X2=3.485 $Y2=2.48
cc_159 N_VDD_M1000_b N_A_c_248_n 0.00244521f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.405
cc_160 N_VDD_M1000_b N_A_c_250_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.405
cc_161 N_VDD_M1000_b N_A_c_252_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.405
cc_162 N_VDD_M1000_b N_A_c_254_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.405
cc_163 N_VDD_M1000_b N_A_c_256_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.405
cc_164 N_VDD_M1000_b N_A_c_258_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=2.625
+ $Y2=2.405
cc_165 N_VDD_M1000_b N_A_c_260_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=3.055
+ $Y2=2.405
cc_166 N_VDD_M1000_s N_A_c_261_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.85
cc_167 N_VDD_M1000_b N_A_c_261_n 0.00618364f $X=-0.045 $Y=2.425 $X2=0.32
+ $Y2=2.85
cc_168 N_VDD_c_118_p N_A_c_261_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_169 N_VDD_M1000_s A 0.0162774f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.845
cc_170 N_VDD_c_118_p A 0.00522047f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.845
cc_171 N_VDD_c_124_p A 9.09141e-19 $X=1.12 $Y=2.955 $X2=0.32 $Y2=2.845
cc_172 N_VDD_M1000_b N_Y_c_474_n 0.00361433f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=2.48
cc_173 N_VDD_c_119_p N_Y_c_474_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69 $Y2=2.48
cc_174 N_VDD_c_120_p N_Y_c_474_n 0.00475776f $X=3.06 $Y=4.25 $X2=0.69 $Y2=2.48
cc_175 N_VDD_M1000_b N_Y_c_477_n 0.00465961f $X=-0.045 $Y=2.425 $X2=1.55
+ $Y2=2.48
cc_176 N_VDD_c_130_p N_Y_c_477_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.48
cc_177 N_VDD_c_120_p N_Y_c_477_n 0.00475776f $X=3.06 $Y=4.25 $X2=1.55 $Y2=2.48
cc_178 N_VDD_M1000_b N_Y_c_480_n 0.00465961f $X=-0.045 $Y=2.425 $X2=2.41
+ $Y2=2.48
cc_179 N_VDD_c_141_p N_Y_c_480_n 0.00734006f $X=2.755 $Y=4.287 $X2=2.41 $Y2=2.48
cc_180 N_VDD_c_120_p N_Y_c_480_n 0.00475776f $X=3.06 $Y=4.25 $X2=2.41 $Y2=2.48
cc_181 N_VDD_M1000_b N_Y_c_483_n 0.00465961f $X=-0.045 $Y=2.425 $X2=3.27
+ $Y2=2.48
cc_182 N_VDD_c_152_p N_Y_c_483_n 0.00745425f $X=3.615 $Y=4.287 $X2=3.27 $Y2=2.48
cc_183 N_VDD_c_120_p N_Y_c_483_n 0.00475776f $X=3.06 $Y=4.25 $X2=3.27 $Y2=2.48
cc_184 N_VDD_M1000_b N_Y_c_486_n 0.00248543f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=2.365
cc_185 N_VDD_M1000_b N_Y_c_487_n 0.00520877f $X=-0.045 $Y=2.425 $X2=1.405
+ $Y2=2.48
cc_186 N_VDD_c_124_p N_Y_c_487_n 0.0090257f $X=1.12 $Y=2.955 $X2=1.405 $Y2=2.48
cc_187 N_VDD_M1000_b N_Y_c_489_n 0.00520877f $X=-0.045 $Y=2.425 $X2=2.265
+ $Y2=2.48
cc_188 N_VDD_c_135_p N_Y_c_489_n 0.0090257f $X=1.98 $Y=2.955 $X2=2.265 $Y2=2.48
cc_189 N_VDD_M1000_b N_Y_c_491_n 0.00409378f $X=-0.045 $Y=2.425 $X2=1.695
+ $Y2=2.48
cc_190 N_VDD_M1000_b N_Y_c_492_n 0.00520877f $X=-0.045 $Y=2.425 $X2=3.125
+ $Y2=2.48
cc_191 N_VDD_c_146_p N_Y_c_492_n 0.0090257f $X=2.84 $Y=2.955 $X2=3.125 $Y2=2.48
cc_192 N_VDD_M1000_b N_Y_c_494_n 0.00409378f $X=-0.045 $Y=2.425 $X2=2.555
+ $Y2=2.48
cc_193 N_VDD_M1000_b N_Y_c_473_n 0.00409378f $X=-0.045 $Y=2.425 $X2=3.27
+ $Y2=2.365
cc_194 A N_Y_M1000_d 0.00250716f $X=0.32 $Y=2.845 $X2=0.55 $Y2=2.605
cc_195 N_A_c_194_n N_Y_c_428_n 0.00182852f $X=0.475 $Y=1.22 $X2=0.69 $Y2=0.755
cc_196 N_A_c_199_n N_Y_c_428_n 0.00251439f $X=0.83 $Y=1.295 $X2=0.69 $Y2=0.755
cc_197 N_A_c_201_n N_Y_c_428_n 0.00182852f $X=0.905 $Y=1.22 $X2=0.69 $Y2=0.755
cc_198 N_A_c_246_n N_Y_c_428_n 3.60975e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.755
cc_199 N_A_c_263_n N_Y_c_428_n 0.00109947f $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.755
cc_200 N_A_c_264_n N_Y_c_474_n 0.00183112f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.48
cc_201 N_A_c_200_n N_Y_c_474_n 0.00899372f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.48
cc_202 N_A_c_269_n N_Y_c_474_n 0.00335296f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.48
cc_203 N_A_c_246_n N_Y_c_474_n 5.06602e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_204 N_A_c_261_n N_Y_c_474_n 0.0226156f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_205 N_A_c_263_n N_Y_c_474_n 0.00165526f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_206 A N_Y_c_474_n 0.00938699f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.48
cc_207 N_A_c_208_n N_Y_c_432_n 0.00182852f $X=1.335 $Y=1.22 $X2=1.55 $Y2=0.755
cc_208 N_A_c_212_n N_Y_c_432_n 0.00310013f $X=1.69 $Y=1.295 $X2=1.55 $Y2=0.755
cc_209 N_A_c_214_n N_Y_c_432_n 0.00182852f $X=1.765 $Y=1.22 $X2=1.55 $Y2=0.755
cc_210 N_A_c_275_n N_Y_c_477_n 0.00335296f $X=1.335 $Y=2.48 $X2=1.55 $Y2=2.48
cc_211 N_A_c_213_n N_Y_c_477_n 0.0108863f $X=1.69 $Y=2.405 $X2=1.55 $Y2=2.48
cc_212 N_A_c_280_n N_Y_c_477_n 0.00335296f $X=1.765 $Y=2.48 $X2=1.55 $Y2=2.48
cc_213 N_A_c_221_n N_Y_c_437_n 0.00182852f $X=2.195 $Y=1.22 $X2=2.41 $Y2=0.755
cc_214 N_A_c_226_n N_Y_c_437_n 0.00310013f $X=2.55 $Y=1.295 $X2=2.41 $Y2=0.755
cc_215 N_A_c_228_n N_Y_c_437_n 0.00182852f $X=2.625 $Y=1.22 $X2=2.41 $Y2=0.755
cc_216 N_A_c_286_n N_Y_c_480_n 0.00335296f $X=2.195 $Y=2.48 $X2=2.41 $Y2=2.48
cc_217 N_A_c_227_n N_Y_c_480_n 0.0108863f $X=2.55 $Y=2.405 $X2=2.41 $Y2=2.48
cc_218 N_A_c_291_n N_Y_c_480_n 0.00335296f $X=2.625 $Y=2.48 $X2=2.41 $Y2=2.48
cc_219 N_A_c_235_n N_Y_c_442_n 0.00182852f $X=3.055 $Y=1.22 $X2=3.27 $Y2=0.755
cc_220 N_A_c_239_n N_Y_c_442_n 0.00310013f $X=3.41 $Y=1.295 $X2=3.27 $Y2=0.755
cc_221 N_A_c_241_n N_Y_c_442_n 0.00182852f $X=3.485 $Y=1.22 $X2=3.27 $Y2=0.755
cc_222 N_A_c_297_n N_Y_c_483_n 0.00335296f $X=3.055 $Y=2.48 $X2=3.27 $Y2=2.48
cc_223 N_A_c_240_n N_Y_c_483_n 0.0105836f $X=3.41 $Y=2.405 $X2=3.27 $Y2=2.48
cc_224 N_A_c_302_n N_Y_c_483_n 0.00335296f $X=3.485 $Y=2.48 $X2=3.27 $Y2=2.48
cc_225 N_A_c_194_n N_Y_c_446_n 0.00880716f $X=0.475 $Y=1.22 $X2=0.69 $Y2=1.115
cc_226 N_A_c_201_n N_Y_c_446_n 0.00198464f $X=0.905 $Y=1.22 $X2=0.69 $Y2=1.115
cc_227 N_A_c_246_n N_Y_c_446_n 0.0011424f $X=0.535 $Y=1.825 $X2=0.69 $Y2=1.115
cc_228 N_A_c_264_n N_Y_c_486_n 0.00169643f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.365
cc_229 N_A_c_200_n N_Y_c_486_n 0.00270155f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.365
cc_230 N_A_c_269_n N_Y_c_486_n 0.00144225f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.365
cc_231 N_A_c_246_n N_Y_c_486_n 8.31386e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.365
cc_232 N_A_c_248_n N_Y_c_486_n 0.00102602f $X=0.475 $Y=2.405 $X2=0.69 $Y2=2.365
cc_233 N_A_c_250_n N_Y_c_486_n 0.00150284f $X=0.905 $Y=2.405 $X2=0.69 $Y2=2.365
cc_234 N_A_c_261_n N_Y_c_486_n 0.0071561f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.365
cc_235 N_A_c_263_n N_Y_c_486_n 0.00173027f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.365
cc_236 A N_Y_c_486_n 0.00805971f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.365
cc_237 N_A_c_194_n Y 0.00150089f $X=0.475 $Y=1.22 $X2=0.76 $Y2=1.72
cc_238 N_A_c_198_n Y 0.00792324f $X=0.475 $Y=2.33 $X2=0.76 $Y2=1.72
cc_239 N_A_c_199_n Y 0.0161013f $X=0.83 $Y=1.295 $X2=0.76 $Y2=1.72
cc_240 N_A_c_200_n Y 0.00363305f $X=0.83 $Y=2.405 $X2=0.76 $Y2=1.72
cc_241 N_A_c_201_n Y 0.00150089f $X=0.905 $Y=1.22 $X2=0.76 $Y2=1.72
cc_242 N_A_c_246_n Y 0.00668675f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_243 N_A_c_247_n Y 0.00675469f $X=0.535 $Y=1.66 $X2=0.76 $Y2=1.72
cc_244 N_A_c_261_n Y 0.0182346f $X=0.32 $Y=2.85 $X2=0.76 $Y2=1.72
cc_245 N_A_c_263_n Y 0.0178517f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_246 N_A_c_201_n N_Y_c_450_n 0.00869047f $X=0.905 $Y=1.22 $X2=1.405 $Y2=1
cc_247 N_A_c_205_n N_Y_c_450_n 0.0022289f $X=1.26 $Y=1.295 $X2=1.405 $Y2=1
cc_248 N_A_c_208_n N_Y_c_450_n 0.00869047f $X=1.335 $Y=1.22 $X2=1.405 $Y2=1
cc_249 N_A_c_269_n N_Y_c_487_n 0.00693713f $X=0.905 $Y=2.48 $X2=1.405 $Y2=2.48
cc_250 N_A_c_207_n N_Y_c_487_n 0.0120397f $X=1.26 $Y=2.405 $X2=1.405 $Y2=2.48
cc_251 N_A_c_275_n N_Y_c_487_n 0.00693713f $X=1.335 $Y=2.48 $X2=1.405 $Y2=2.48
cc_252 N_A_c_250_n N_Y_c_487_n 0.00560085f $X=0.905 $Y=2.405 $X2=1.405 $Y2=2.48
cc_253 N_A_c_252_n N_Y_c_487_n 0.00560085f $X=1.335 $Y=2.405 $X2=1.405 $Y2=2.48
cc_254 N_A_c_208_n N_Y_c_454_n 0.00150089f $X=1.335 $Y=1.22 $X2=1.55 $Y2=2.365
cc_255 N_A_c_212_n N_Y_c_454_n 0.0177499f $X=1.69 $Y=1.295 $X2=1.55 $Y2=2.365
cc_256 N_A_c_213_n N_Y_c_454_n 0.00562481f $X=1.69 $Y=2.405 $X2=1.55 $Y2=2.365
cc_257 N_A_c_214_n N_Y_c_454_n 0.00150089f $X=1.765 $Y=1.22 $X2=1.55 $Y2=2.365
cc_258 N_A_c_225_n N_Y_c_454_n 0.0141566f $X=2.195 $Y=2.33 $X2=1.55 $Y2=2.365
cc_259 N_A_c_214_n N_Y_c_455_n 0.00869047f $X=1.765 $Y=1.22 $X2=2.265 $Y2=1
cc_260 N_A_c_218_n N_Y_c_455_n 0.0022289f $X=2.12 $Y=1.295 $X2=2.265 $Y2=1
cc_261 N_A_c_221_n N_Y_c_455_n 0.00938169f $X=2.195 $Y=1.22 $X2=2.265 $Y2=1
cc_262 N_A_c_208_n N_Y_c_459_n 0.00198464f $X=1.335 $Y=1.22 $X2=1.695 $Y2=1
cc_263 N_A_c_214_n N_Y_c_459_n 0.00198464f $X=1.765 $Y=1.22 $X2=1.695 $Y2=1
cc_264 N_A_c_280_n N_Y_c_489_n 0.00693713f $X=1.765 $Y=2.48 $X2=2.265 $Y2=2.48
cc_265 N_A_c_220_n N_Y_c_489_n 0.0125508f $X=2.12 $Y=2.405 $X2=2.265 $Y2=2.48
cc_266 N_A_c_286_n N_Y_c_489_n 0.00693713f $X=2.195 $Y=2.48 $X2=2.265 $Y2=2.48
cc_267 N_A_c_254_n N_Y_c_489_n 0.00560085f $X=1.765 $Y=2.405 $X2=2.265 $Y2=2.48
cc_268 N_A_c_256_n N_Y_c_489_n 0.00642784f $X=2.195 $Y=2.405 $X2=2.265 $Y2=2.48
cc_269 N_A_c_275_n N_Y_c_491_n 0.00144225f $X=1.335 $Y=2.48 $X2=1.695 $Y2=2.48
cc_270 N_A_c_213_n N_Y_c_491_n 0.00397642f $X=1.69 $Y=2.405 $X2=1.695 $Y2=2.48
cc_271 N_A_c_280_n N_Y_c_491_n 0.00144225f $X=1.765 $Y=2.48 $X2=1.695 $Y2=2.48
cc_272 N_A_c_252_n N_Y_c_491_n 0.00150284f $X=1.335 $Y=2.405 $X2=1.695 $Y2=2.48
cc_273 N_A_c_254_n N_Y_c_491_n 0.00150284f $X=1.765 $Y=2.405 $X2=1.695 $Y2=2.48
cc_274 N_A_c_221_n N_Y_c_462_n 0.00150089f $X=2.195 $Y=1.22 $X2=2.41 $Y2=2.365
cc_275 N_A_c_225_n N_Y_c_462_n 0.0182294f $X=2.195 $Y=2.33 $X2=2.41 $Y2=2.365
cc_276 N_A_c_226_n N_Y_c_462_n 0.0177499f $X=2.55 $Y=1.295 $X2=2.41 $Y2=2.365
cc_277 N_A_c_227_n N_Y_c_462_n 0.00562481f $X=2.55 $Y=2.405 $X2=2.41 $Y2=2.365
cc_278 N_A_c_228_n N_Y_c_462_n 0.00150089f $X=2.625 $Y=1.22 $X2=2.41 $Y2=2.365
cc_279 N_A_c_228_n N_Y_c_463_n 0.00869047f $X=2.625 $Y=1.22 $X2=3.125 $Y2=1
cc_280 N_A_c_232_n N_Y_c_463_n 0.0022289f $X=2.98 $Y=1.295 $X2=3.125 $Y2=1
cc_281 N_A_c_235_n N_Y_c_463_n 0.00869047f $X=3.055 $Y=1.22 $X2=3.125 $Y2=1
cc_282 N_A_c_221_n N_Y_c_467_n 0.00201073f $X=2.195 $Y=1.22 $X2=2.555 $Y2=1
cc_283 N_A_c_228_n N_Y_c_467_n 0.00198464f $X=2.625 $Y=1.22 $X2=2.555 $Y2=1
cc_284 N_A_c_291_n N_Y_c_492_n 0.00693713f $X=2.625 $Y=2.48 $X2=3.125 $Y2=2.48
cc_285 N_A_c_234_n N_Y_c_492_n 0.0120397f $X=2.98 $Y=2.405 $X2=3.125 $Y2=2.48
cc_286 N_A_c_297_n N_Y_c_492_n 0.00693713f $X=3.055 $Y=2.48 $X2=3.125 $Y2=2.48
cc_287 N_A_c_258_n N_Y_c_492_n 0.00560085f $X=2.625 $Y=2.405 $X2=3.125 $Y2=2.48
cc_288 N_A_c_260_n N_Y_c_492_n 0.00560085f $X=3.055 $Y=2.405 $X2=3.125 $Y2=2.48
cc_289 N_A_c_286_n N_Y_c_494_n 0.00144225f $X=2.195 $Y=2.48 $X2=2.555 $Y2=2.48
cc_290 N_A_c_227_n N_Y_c_494_n 0.00397642f $X=2.55 $Y=2.405 $X2=2.555 $Y2=2.48
cc_291 N_A_c_291_n N_Y_c_494_n 0.00144225f $X=2.625 $Y=2.48 $X2=2.555 $Y2=2.48
cc_292 N_A_c_256_n N_Y_c_494_n 0.00153387f $X=2.195 $Y=2.405 $X2=2.555 $Y2=2.48
cc_293 N_A_c_258_n N_Y_c_494_n 0.00150284f $X=2.625 $Y=2.405 $X2=2.555 $Y2=2.48
cc_294 N_A_c_235_n N_Y_c_470_n 0.00198464f $X=3.055 $Y=1.22 $X2=3.27 $Y2=1.115
cc_295 N_A_c_241_n N_Y_c_470_n 0.00878106f $X=3.485 $Y=1.22 $X2=3.27 $Y2=1.115
cc_296 N_A_c_235_n N_Y_c_473_n 0.00150089f $X=3.055 $Y=1.22 $X2=3.27 $Y2=2.365
cc_297 N_A_c_297_n N_Y_c_473_n 0.00144225f $X=3.055 $Y=2.48 $X2=3.27 $Y2=2.365
cc_298 N_A_c_239_n N_Y_c_473_n 0.0169795f $X=3.41 $Y=1.295 $X2=3.27 $Y2=2.365
cc_299 N_A_c_240_n N_Y_c_473_n 0.0141541f $X=3.41 $Y=2.405 $X2=3.27 $Y2=2.365
cc_300 N_A_c_241_n N_Y_c_473_n 0.00150089f $X=3.485 $Y=1.22 $X2=3.27 $Y2=2.365
cc_301 N_A_c_302_n N_Y_c_473_n 0.00541616f $X=3.485 $Y=2.48 $X2=3.27 $Y2=2.365
cc_302 N_A_c_260_n N_Y_c_473_n 0.00150284f $X=3.055 $Y=2.405 $X2=3.27 $Y2=2.365
