* File: sky130_osu_sc_12T_hs__dffsr_1.pxi.spice
* Created: Fri Nov 12 15:09:47 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%GND N_GND_M1016_s N_GND_M1034_s N_GND_M1003_d
+ N_GND_M1005_s N_GND_M1020_d N_GND_M1006_d N_GND_M1013_s N_GND_M1022_d
+ N_GND_M1007_d N_GND_M1016_b N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_13_p
+ N_GND_c_50_p N_GND_c_51_p N_GND_c_52_p N_GND_c_53_p N_GND_c_54_p N_GND_c_55_p
+ N_GND_c_56_p N_GND_c_57_p N_GND_c_58_p N_GND_c_16_p N_GND_c_17_p N_GND_c_61_p
+ N_GND_c_204_p GND N_GND_c_5_p PM_SKY130_OSU_SC_12T_HS__DFFSR_1%GND
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%VDD N_VDD_M1001_s N_VDD_M1024_d N_VDD_M1028_s
+ N_VDD_M1009_d N_VDD_M1029_d N_VDD_M1033_d N_VDD_M1030_d N_VDD_M1001_b
+ N_VDD_c_267_p N_VDD_c_268_p N_VDD_c_287_p N_VDD_c_311_p N_VDD_c_304_p
+ N_VDD_c_322_p N_VDD_c_305_p N_VDD_c_332_p N_VDD_c_306_p N_VDD_c_337_p
+ N_VDD_c_290_p N_VDD_c_279_p N_VDD_c_376_p N_VDD_c_399_p VDD N_VDD_c_269_p
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%VDD
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%RN N_RN_M1016_g N_RN_c_436_n N_RN_M1001_g
+ N_RN_c_438_n N_RN_c_439_n RN PM_SKY130_OSU_SC_12T_HS__DFFSR_1%RN
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_110_115# N_A_110_115#_M1016_d
+ N_A_110_115#_M1001_d N_A_110_115#_c_473_n N_A_110_115#_M1000_g
+ N_A_110_115#_c_474_n N_A_110_115#_M1034_g N_A_110_115#_c_478_n
+ N_A_110_115#_M1022_g N_A_110_115#_M1025_g N_A_110_115#_c_483_n
+ N_A_110_115#_c_484_n N_A_110_115#_c_485_n N_A_110_115#_c_487_n
+ N_A_110_115#_c_489_n N_A_110_115#_c_490_n N_A_110_115#_c_494_n
+ N_A_110_115#_c_495_n N_A_110_115#_c_496_n N_A_110_115#_c_497_n
+ N_A_110_115#_c_499_n N_A_110_115#_c_500_n N_A_110_115#_c_502_n
+ N_A_110_115#_c_503_n N_A_110_115#_c_525_n N_A_110_115#_c_527_n
+ N_A_110_115#_c_528_n N_A_110_115#_c_529_n
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_110_115#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%SN N_SN_c_703_n N_SN_c_704_n N_SN_M1024_g
+ N_SN_M1015_g N_SN_M1004_g N_SN_M1019_g N_SN_c_713_n N_SN_c_714_n N_SN_c_715_n
+ N_SN_c_716_n N_SN_c_730_n N_SN_c_717_n N_SN_c_732_n N_SN_c_718_n N_SN_c_719_n
+ N_SN_c_733_n N_SN_c_742_n SN PM_SKY130_OSU_SC_12T_HS__DFFSR_1%SN
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_432_424# N_A_432_424#_M1035_d
+ N_A_432_424#_M1018_d N_A_432_424#_M1003_g N_A_432_424#_M1027_g
+ N_A_432_424#_c_900_n N_A_432_424#_c_901_n N_A_432_424#_c_902_n
+ N_A_432_424#_c_905_n N_A_432_424#_c_906_n N_A_432_424#_c_907_n
+ N_A_432_424#_c_920_n N_A_432_424#_c_923_n N_A_432_424#_c_908_n
+ N_A_432_424#_c_924_n N_A_432_424#_c_909_n
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_432_424#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%D N_D_M1005_g N_D_M1028_g N_D_c_1010_n
+ N_D_c_1011_n D PM_SKY130_OSU_SC_12T_HS__DFFSR_1%D
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%CK N_CK_M1018_g N_CK_M1026_g N_CK_M1021_g
+ N_CK_M1002_g N_CK_M1011_g N_CK_c_1043_n N_CK_M1031_g N_CK_c_1044_n
+ N_CK_c_1045_n N_CK_c_1046_n N_CK_c_1047_n N_CK_c_1050_n N_CK_c_1051_n
+ N_CK_c_1054_n N_CK_c_1055_n N_CK_c_1060_n N_CK_c_1061_n N_CK_c_1062_n
+ N_CK_c_1063_n N_CK_c_1064_n N_CK_c_1065_n N_CK_c_1066_n N_CK_c_1067_n
+ N_CK_c_1068_n N_CK_c_1069_n N_CK_c_1070_n N_CK_c_1071_n N_CK_c_1072_n CK
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%CK
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_217_521# N_A_217_521#_M1034_d
+ N_A_217_521#_M1000_s N_A_217_521#_M1020_g N_A_217_521#_M1009_g
+ N_A_217_521#_c_1300_n N_A_217_521#_c_1302_n N_A_217_521#_c_1303_n
+ N_A_217_521#_c_1304_n N_A_217_521#_M1023_g N_A_217_521#_M1012_g
+ N_A_217_521#_c_1309_n N_A_217_521#_c_1310_n N_A_217_521#_c_1311_n
+ N_A_217_521#_c_1312_n N_A_217_521#_c_1315_n N_A_217_521#_c_1316_n
+ N_A_217_521#_c_1317_n N_A_217_521#_c_1319_n N_A_217_521#_c_1320_n
+ N_A_217_521#_c_1372_n PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_217_521#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_704_89# N_A_704_89#_M1011_d
+ N_A_704_89#_M1031_d N_A_704_89#_c_1460_n N_A_704_89#_M1035_g
+ N_A_704_89#_c_1463_n N_A_704_89#_c_1464_n N_A_704_89#_c_1465_n
+ N_A_704_89#_M1014_g N_A_704_89#_c_1467_n N_A_704_89#_M1010_g
+ N_A_704_89#_c_1469_n N_A_704_89#_M1017_g N_A_704_89#_c_1473_n
+ N_A_704_89#_c_1474_n N_A_704_89#_c_1475_n N_A_704_89#_c_1476_n
+ N_A_704_89#_c_1477_n N_A_704_89#_c_1478_n N_A_704_89#_c_1494_n
+ N_A_704_89#_c_1483_n N_A_704_89#_c_1484_n N_A_704_89#_c_1499_n
+ N_A_704_89#_c_1485_n N_A_704_89#_c_1486_n N_A_704_89#_c_1487_n
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_704_89#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1246_89# N_A_1246_89#_M1004_d
+ N_A_1246_89#_M1025_d N_A_1246_89#_M1006_g N_A_1246_89#_M1029_g
+ N_A_1246_89#_M1007_g N_A_1246_89#_M1030_g N_A_1246_89#_c_1677_n
+ N_A_1246_89#_c_1679_n N_A_1246_89#_c_1680_n N_A_1246_89#_c_1681_n
+ N_A_1246_89#_c_1686_n N_A_1246_89#_c_1687_n N_A_1246_89#_c_1688_n
+ N_A_1246_89#_c_1689_n N_A_1246_89#_c_1690_n N_A_1246_89#_c_1693_n
+ N_A_1246_89#_c_1694_n N_A_1246_89#_c_1695_n N_A_1246_89#_c_1696_n
+ N_A_1246_89#_c_1697_n N_A_1246_89#_c_1698_n N_A_1246_89#_c_1699_n
+ N_A_1246_89#_c_1700_n N_A_1246_89#_c_1701_n
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1246_89#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1084_115# N_A_1084_115#_M1021_d
+ N_A_1084_115#_M1010_d N_A_1084_115#_c_1883_n N_A_1084_115#_c_1884_n
+ N_A_1084_115#_M1013_g N_A_1084_115#_M1033_g N_A_1084_115#_c_1888_n
+ N_A_1084_115#_c_1890_n N_A_1084_115#_c_1891_n N_A_1084_115#_c_1941_n
+ N_A_1084_115#_c_1942_n N_A_1084_115#_c_1911_n N_A_1084_115#_c_1892_n
+ N_A_1084_115#_c_1893_n N_A_1084_115#_c_1895_n N_A_1084_115#_c_1898_n
+ N_A_1084_115#_c_1899_n N_A_1084_115#_c_1900_n N_A_1084_115#_c_1903_n
+ N_A_1084_115#_c_1904_n PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1084_115#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%QN N_QN_M1007_s N_QN_M1030_s N_QN_M1008_g
+ N_QN_M1032_g N_QN_c_2064_n N_QN_c_2065_n N_QN_c_2069_n N_QN_c_2070_n
+ N_QN_c_2072_n N_QN_c_2073_n N_QN_c_2074_n N_QN_c_2075_n QN
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%QN
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_300_521# N_A_300_521#_M1000_d
+ N_A_300_521#_M1027_d N_A_300_521#_c_2143_n N_A_300_521#_c_2146_n
+ N_A_300_521#_c_2159_n N_A_300_521#_c_2149_n
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_300_521#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1469_521# N_A_1469_521#_M1033_s
+ N_A_1469_521#_M1019_d N_A_1469_521#_c_2171_n N_A_1469_521#_c_2174_n
+ N_A_1469_521#_c_2184_n N_A_1469_521#_c_2176_n
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1469_521#
x_PM_SKY130_OSU_SC_12T_HS__DFFSR_1%Q N_Q_M1008_d N_Q_M1032_d N_Q_c_2191_n
+ N_Q_c_2195_n N_Q_c_2193_n N_Q_c_2194_n N_Q_c_2199_n Q
+ PM_SKY130_OSU_SC_12T_HS__DFFSR_1%Q
cc_1 N_GND_M1016_b N_RN_M1016_g 0.0605175f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_RN_M1016_g 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_RN_M1016_g 0.00606474f $X=1.135 $Y=0.152 $X2=0.475 $Y2=0.85
cc_4 N_GND_c_4_p N_RN_M1016_g 0.0035726f $X=1.22 $Y=0.74 $X2=0.475 $Y2=0.85
cc_5 N_GND_c_5_p N_RN_M1016_g 0.00468827f $X=9.855 $Y=0.19 $X2=0.475 $Y2=0.85
cc_6 N_GND_M1016_b N_RN_c_436_n 0.0366269f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.99
cc_7 N_GND_M1016_b N_RN_M1001_g 0.0318753f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.235
cc_8 N_GND_M1016_b N_RN_c_438_n 0.0149094f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_9 N_GND_M1016_b N_RN_c_439_n 0.0202952f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.825
cc_10 N_GND_M1016_b N_A_110_115#_c_473_n 0.05194f $X=-0.05 $Y=0 $X2=1.29
+ $Y2=2.32
cc_11 N_GND_M1016_b N_A_110_115#_c_474_n 0.0186674f $X=-0.05 $Y=0 $X2=1.435
+ $Y2=1.105
cc_12 N_GND_c_4_p N_A_110_115#_c_474_n 0.00502587f $X=1.22 $Y=0.74 $X2=1.435
+ $Y2=1.105
cc_13 N_GND_c_13_p N_A_110_115#_c_474_n 0.00606474f $X=2.415 $Y=0.152 $X2=1.435
+ $Y2=1.105
cc_14 N_GND_c_5_p N_A_110_115#_c_474_n 0.00468827f $X=9.855 $Y=0.19 $X2=1.435
+ $Y2=1.105
cc_15 N_GND_M1016_b N_A_110_115#_c_478_n 0.0186674f $X=-0.05 $Y=0 $X2=8.535
+ $Y2=1.105
cc_16 N_GND_c_16_p N_A_110_115#_c_478_n 0.00606474f $X=8.665 $Y=0.152 $X2=8.535
+ $Y2=1.105
cc_17 N_GND_c_17_p N_A_110_115#_c_478_n 0.00502587f $X=8.75 $Y=0.74 $X2=8.535
+ $Y2=1.105
cc_18 N_GND_c_5_p N_A_110_115#_c_478_n 0.00468827f $X=9.855 $Y=0.19 $X2=8.535
+ $Y2=1.105
cc_19 N_GND_M1016_b N_A_110_115#_M1025_g 5.06705e-19 $X=-0.05 $Y=0 $X2=8.545
+ $Y2=3.235
cc_20 N_GND_M1016_b N_A_110_115#_c_483_n 0.0419907f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=2.125
cc_21 N_GND_M1016_b N_A_110_115#_c_484_n 0.0124725f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=2.395
cc_22 N_GND_M1016_b N_A_110_115#_c_485_n 0.0425388f $X=-0.05 $Y=0 $X2=1.29
+ $Y2=1.27
cc_23 N_GND_c_4_p N_A_110_115#_c_485_n 0.00438982f $X=1.22 $Y=0.74 $X2=1.29
+ $Y2=1.27
cc_24 N_GND_M1016_b N_A_110_115#_c_487_n 0.0510808f $X=-0.05 $Y=0 $X2=8.8
+ $Y2=1.27
cc_25 N_GND_c_17_p N_A_110_115#_c_487_n 0.0043356f $X=8.75 $Y=0.74 $X2=8.8
+ $Y2=1.27
cc_26 N_GND_M1016_b N_A_110_115#_c_489_n 0.0393083f $X=-0.05 $Y=0 $X2=8.545
+ $Y2=2.27
cc_27 N_GND_M1016_b N_A_110_115#_c_490_n 0.00307511f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=0.755
cc_28 N_GND_c_3_p N_A_110_115#_c_490_n 0.00751834f $X=1.135 $Y=0.152 $X2=0.69
+ $Y2=0.755
cc_29 N_GND_c_4_p N_A_110_115#_c_490_n 0.013807f $X=1.22 $Y=0.74 $X2=0.69
+ $Y2=0.755
cc_30 N_GND_c_5_p N_A_110_115#_c_490_n 0.00474566f $X=9.855 $Y=0.19 $X2=0.69
+ $Y2=0.755
cc_31 N_GND_M1016_b N_A_110_115#_c_494_n 0.00213782f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=2.955
cc_32 N_GND_M1016_b N_A_110_115#_c_495_n 0.0176591f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=1.37
cc_33 N_GND_M1016_b N_A_110_115#_c_496_n 0.0102253f $X=-0.05 $Y=0 $X2=0.955
+ $Y2=1.27
cc_34 N_GND_M1016_b N_A_110_115#_c_497_n 0.00577265f $X=-0.05 $Y=0 $X2=1.23
+ $Y2=1.27
cc_35 N_GND_c_4_p N_A_110_115#_c_497_n 0.00544663f $X=1.22 $Y=0.74 $X2=1.23
+ $Y2=1.27
cc_36 N_GND_M1016_b N_A_110_115#_c_499_n 0.0161505f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.26
cc_37 N_GND_M1016_b N_A_110_115#_c_500_n 0.00388815f $X=-0.05 $Y=0 $X2=8.86
+ $Y2=1.27
cc_38 N_GND_c_17_p N_A_110_115#_c_500_n 0.00481479f $X=8.75 $Y=0.74 $X2=8.86
+ $Y2=1.27
cc_39 N_GND_M1016_b N_A_110_115#_c_502_n 0.00181375f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=1.255
cc_40 N_GND_M1034_s N_A_110_115#_c_503_n 0.00271747f $X=1.095 $Y=0.575 $X2=8.775
+ $Y2=1
cc_41 N_GND_M1003_d N_A_110_115#_c_503_n 0.00263306f $X=2.36 $Y=0.575 $X2=8.775
+ $Y2=1
cc_42 N_GND_M1005_s N_A_110_115#_c_503_n 0.00263312f $X=2.895 $Y=0.575 $X2=8.775
+ $Y2=1
cc_43 N_GND_M1020_d N_A_110_115#_c_503_n 0.00724592f $X=4.63 $Y=0.575 $X2=8.775
+ $Y2=1
cc_44 N_GND_M1006_d N_A_110_115#_c_503_n 0.00370555f $X=6.38 $Y=0.575 $X2=8.775
+ $Y2=1
cc_45 N_GND_M1013_s N_A_110_115#_c_503_n 0.00321993f $X=7.345 $Y=0.575 $X2=8.775
+ $Y2=1
cc_46 N_GND_M1022_d N_A_110_115#_c_503_n 0.00282782f $X=8.61 $Y=0.575 $X2=8.775
+ $Y2=1
cc_47 N_GND_M1016_b N_A_110_115#_c_503_n 0.0201213f $X=-0.05 $Y=0 $X2=8.775
+ $Y2=1
cc_48 N_GND_c_4_p N_A_110_115#_c_503_n 0.00597331f $X=1.22 $Y=0.74 $X2=8.775
+ $Y2=1
cc_49 N_GND_c_13_p N_A_110_115#_c_503_n 0.0148659f $X=2.415 $Y=0.152 $X2=8.775
+ $Y2=1
cc_50 N_GND_c_50_p N_A_110_115#_c_503_n 0.0118179f $X=2.5 $Y=0.755 $X2=8.775
+ $Y2=1
cc_51 N_GND_c_51_p N_A_110_115#_c_503_n 0.00599718f $X=2.935 $Y=0.152 $X2=8.775
+ $Y2=1
cc_52 N_GND_c_52_p N_A_110_115#_c_503_n 0.0118113f $X=3.02 $Y=0.755 $X2=8.775
+ $Y2=1
cc_53 N_GND_c_53_p N_A_110_115#_c_503_n 0.0196453f $X=4.685 $Y=0.152 $X2=8.775
+ $Y2=1
cc_54 N_GND_c_54_p N_A_110_115#_c_503_n 0.007301f $X=4.77 $Y=0.74 $X2=8.775
+ $Y2=1
cc_55 N_GND_c_55_p N_A_110_115#_c_503_n 0.0196423f $X=6.435 $Y=0.152 $X2=8.775
+ $Y2=1
cc_56 N_GND_c_56_p N_A_110_115#_c_503_n 0.0143043f $X=6.52 $Y=0.755 $X2=8.775
+ $Y2=1
cc_57 N_GND_c_57_p N_A_110_115#_c_503_n 0.0102455f $X=7.385 $Y=0.152 $X2=8.775
+ $Y2=1
cc_58 N_GND_c_58_p N_A_110_115#_c_503_n 0.0139059f $X=7.47 $Y=0.755 $X2=8.775
+ $Y2=1
cc_59 N_GND_c_16_p N_A_110_115#_c_503_n 0.0148659f $X=8.665 $Y=0.152 $X2=8.775
+ $Y2=1
cc_60 N_GND_c_17_p N_A_110_115#_c_503_n 0.00714169f $X=8.75 $Y=0.74 $X2=8.775
+ $Y2=1
cc_61 N_GND_c_61_p N_A_110_115#_c_503_n 0.00233122f $X=9.625 $Y=0.152 $X2=8.775
+ $Y2=1
cc_62 N_GND_M1016_b N_A_110_115#_c_525_n 0.00246937f $X=-0.05 $Y=0 $X2=0.955
+ $Y2=1
cc_63 N_GND_c_3_p N_A_110_115#_c_525_n 0.00667461f $X=1.135 $Y=0.152 $X2=0.955
+ $Y2=1
cc_64 N_GND_M1016_b N_A_110_115#_c_527_n 0.00747477f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=1.37
cc_65 N_GND_M1016_b N_A_110_115#_c_528_n 0.00268886f $X=-0.05 $Y=0 $X2=8.86
+ $Y2=1.37
cc_66 N_GND_M1016_b N_A_110_115#_c_529_n 3.28821e-19 $X=-0.05 $Y=0 $X2=8.862
+ $Y2=1.255
cc_67 N_GND_M1016_b N_SN_c_703_n 0.00804573f $X=-0.05 $Y=0 $X2=1.89 $Y2=1.405
cc_68 N_GND_M1016_b N_SN_c_704_n 0.0220657f $X=-0.05 $Y=0 $X2=1.89 $Y2=1.785
cc_69 N_GND_M1016_b N_SN_M1024_g 0.0152105f $X=-0.05 $Y=0 $X2=1.855 $Y2=3.235
cc_70 N_GND_M1016_b N_SN_M1015_g 0.0196935f $X=-0.05 $Y=0 $X2=1.925 $Y2=0.85
cc_71 N_GND_c_13_p N_SN_M1015_g 0.00606474f $X=2.415 $Y=0.152 $X2=1.925 $Y2=0.85
cc_72 N_GND_c_5_p N_SN_M1015_g 0.00468827f $X=9.855 $Y=0.19 $X2=1.925 $Y2=0.85
cc_73 N_GND_M1016_b N_SN_M1004_g 0.0405285f $X=-0.05 $Y=0 $X2=8.045 $Y2=0.85
cc_74 N_GND_c_16_p N_SN_M1004_g 0.00606474f $X=8.665 $Y=0.152 $X2=8.045 $Y2=0.85
cc_75 N_GND_c_5_p N_SN_M1004_g 0.00468827f $X=9.855 $Y=0.19 $X2=8.045 $Y2=0.85
cc_76 N_GND_M1016_b N_SN_M1019_g 0.0293574f $X=-0.05 $Y=0 $X2=8.115 $Y2=3.235
cc_77 N_GND_M1016_b N_SN_c_713_n 0.0384463f $X=-0.05 $Y=0 $X2=1.855 $Y2=1.95
cc_78 N_GND_M1016_b N_SN_c_714_n 0.0354748f $X=-0.05 $Y=0 $X2=8.02 $Y2=1.775
cc_79 N_GND_M1016_b N_SN_c_715_n 0.00238535f $X=-0.05 $Y=0 $X2=1.71 $Y2=2.62
cc_80 N_GND_M1016_b N_SN_c_716_n 6.25411e-19 $X=-0.05 $Y=0 $X2=7.937 $Y2=2.482
cc_81 N_GND_M1016_b N_SN_c_717_n 0.00242182f $X=-0.05 $Y=0 $X2=1.71 $Y2=1.95
cc_82 N_GND_M1016_b N_SN_c_718_n 0.00158638f $X=-0.05 $Y=0 $X2=8.02 $Y2=1.775
cc_83 N_GND_M1016_b N_SN_c_719_n 0.00848267f $X=-0.05 $Y=0 $X2=7.937 $Y2=2.395
cc_84 N_GND_M1016_b N_A_432_424#_M1003_g 0.0716031f $X=-0.05 $Y=0 $X2=2.285
+ $Y2=0.85
cc_85 N_GND_c_13_p N_A_432_424#_M1003_g 0.00606474f $X=2.415 $Y=0.152 $X2=2.285
+ $Y2=0.85
cc_86 N_GND_c_50_p N_A_432_424#_M1003_g 0.00509667f $X=2.5 $Y=0.755 $X2=2.285
+ $Y2=0.85
cc_87 N_GND_c_5_p N_A_432_424#_M1003_g 0.00468827f $X=9.855 $Y=0.19 $X2=2.285
+ $Y2=0.85
cc_88 N_GND_M1016_b N_A_432_424#_c_900_n 0.0299799f $X=-0.05 $Y=0 $X2=2.295
+ $Y2=2.285
cc_89 N_GND_M1016_b N_A_432_424#_c_901_n 0.0239207f $X=-0.05 $Y=0 $X2=2.295
+ $Y2=2.2
cc_90 N_GND_M1016_b N_A_432_424#_c_902_n 0.027997f $X=-0.05 $Y=0 $X2=3.71
+ $Y2=1.285
cc_91 N_GND_c_50_p N_A_432_424#_c_902_n 0.00673409f $X=2.5 $Y=0.755 $X2=3.71
+ $Y2=1.285
cc_92 N_GND_c_52_p N_A_432_424#_c_902_n 0.00673409f $X=3.02 $Y=0.755 $X2=3.71
+ $Y2=1.285
cc_93 N_GND_M1016_b N_A_432_424#_c_905_n 0.00154034f $X=-0.05 $Y=0 $X2=2.38
+ $Y2=1.285
cc_94 N_GND_M1016_b N_A_432_424#_c_906_n 0.0227986f $X=-0.05 $Y=0 $X2=2.685
+ $Y2=2.285
cc_95 N_GND_M1016_b N_A_432_424#_c_907_n 0.00124354f $X=-0.05 $Y=0 $X2=2.77
+ $Y2=2.62
cc_96 N_GND_M1016_b N_A_432_424#_c_908_n 0.00140975f $X=-0.05 $Y=0 $X2=3.795
+ $Y2=1.2
cc_97 N_GND_M1016_b N_A_432_424#_c_909_n 0.00311983f $X=-0.05 $Y=0 $X2=3.795
+ $Y2=0.755
cc_98 N_GND_c_53_p N_A_432_424#_c_909_n 0.0146486f $X=4.685 $Y=0.152 $X2=3.795
+ $Y2=0.755
cc_99 N_GND_c_5_p N_A_432_424#_c_909_n 0.0098977f $X=9.855 $Y=0.19 $X2=3.795
+ $Y2=0.755
cc_100 N_GND_M1016_b N_D_M1005_g 0.0417362f $X=-0.05 $Y=0 $X2=3.235 $Y2=0.85
cc_101 N_GND_c_52_p N_D_M1005_g 0.00509529f $X=3.02 $Y=0.755 $X2=3.235 $Y2=0.85
cc_102 N_GND_c_53_p N_D_M1005_g 0.00606474f $X=4.685 $Y=0.152 $X2=3.235 $Y2=0.85
cc_103 N_GND_c_5_p N_D_M1005_g 0.00468827f $X=9.855 $Y=0.19 $X2=3.235 $Y2=0.85
cc_104 N_GND_M1016_b N_D_M1028_g 0.0397275f $X=-0.05 $Y=0 $X2=3.235 $Y2=3.235
cc_105 N_GND_M1016_b N_D_c_1010_n 0.0342074f $X=-0.05 $Y=0 $X2=3.295 $Y2=1.74
cc_106 N_GND_M1016_b N_D_c_1011_n 0.00311208f $X=-0.05 $Y=0 $X2=3.295 $Y2=1.74
cc_107 N_GND_M1016_b D 0.0160302f $X=-0.05 $Y=0 $X2=3.295 $Y2=1.74
cc_108 N_GND_M1016_b N_CK_c_1043_n 0.0293731f $X=-0.05 $Y=0 $X2=6.735 $Y2=2.45
cc_109 N_GND_M1016_b N_CK_c_1044_n 0.0430736f $X=-0.05 $Y=0 $X2=6.79 $Y2=2.12
cc_110 N_GND_M1016_b N_CK_c_1045_n 0.0247714f $X=-0.05 $Y=0 $X2=3.685 $Y2=2.285
cc_111 N_GND_M1016_b N_CK_c_1046_n 0.0254952f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.4
cc_112 N_GND_M1016_b N_CK_c_1047_n 0.017381f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.235
cc_113 N_GND_c_53_p N_CK_c_1047_n 0.00606474f $X=4.685 $Y=0.152 $X2=4.135
+ $Y2=1.235
cc_114 N_GND_c_5_p N_CK_c_1047_n 0.00468827f $X=9.855 $Y=0.19 $X2=4.135
+ $Y2=1.235
cc_115 N_GND_M1016_b N_CK_c_1050_n 0.026818f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.4
cc_116 N_GND_M1016_b N_CK_c_1051_n 0.0174883f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.235
cc_117 N_GND_c_55_p N_CK_c_1051_n 0.00606474f $X=6.435 $Y=0.152 $X2=5.405
+ $Y2=1.235
cc_118 N_GND_c_5_p N_CK_c_1051_n 0.00468827f $X=9.855 $Y=0.19 $X2=5.405
+ $Y2=1.235
cc_119 N_GND_M1016_b N_CK_c_1054_n 0.0223817f $X=-0.05 $Y=0 $X2=5.855 $Y2=2.285
cc_120 N_GND_M1016_b N_CK_c_1055_n 0.0166942f $X=-0.05 $Y=0 $X2=6.762 $Y2=1.205
cc_121 N_GND_c_56_p N_CK_c_1055_n 0.00311745f $X=6.52 $Y=0.755 $X2=6.762
+ $Y2=1.205
cc_122 N_GND_c_57_p N_CK_c_1055_n 0.00606474f $X=7.385 $Y=0.152 $X2=6.762
+ $Y2=1.205
cc_123 N_GND_c_58_p N_CK_c_1055_n 0.00363995f $X=7.47 $Y=0.755 $X2=6.762
+ $Y2=1.205
cc_124 N_GND_c_5_p N_CK_c_1055_n 0.00468827f $X=9.855 $Y=0.19 $X2=6.762
+ $Y2=1.205
cc_125 N_GND_M1016_b N_CK_c_1060_n 0.0135081f $X=-0.05 $Y=0 $X2=6.762 $Y2=1.355
cc_126 N_GND_M1016_b N_CK_c_1061_n 0.00530209f $X=-0.05 $Y=0 $X2=4.05 $Y2=2.11
cc_127 N_GND_M1016_b N_CK_c_1062_n 0.00837891f $X=-0.05 $Y=0 $X2=4.135 $Y2=1.4
cc_128 N_GND_M1016_b N_CK_c_1063_n 0.0068355f $X=-0.05 $Y=0 $X2=5.405 $Y2=1.4
cc_129 N_GND_M1016_b N_CK_c_1064_n 0.00430942f $X=-0.05 $Y=0 $X2=5.77 $Y2=2.11
cc_130 N_GND_M1016_b N_CK_c_1065_n 5.00459e-19 $X=-0.05 $Y=0 $X2=5.49 $Y2=2.11
cc_131 N_GND_M1016_b N_CK_c_1066_n 7.36568e-19 $X=-0.05 $Y=0 $X2=6.88 $Y2=2.11
cc_132 N_GND_M1016_b N_CK_c_1067_n 0.00346455f $X=-0.05 $Y=0 $X2=3.655 $Y2=2.11
cc_133 N_GND_M1016_b N_CK_c_1068_n 0.00155168f $X=-0.05 $Y=0 $X2=5.885 $Y2=2.11
cc_134 N_GND_M1016_b N_CK_c_1069_n 0.0328755f $X=-0.05 $Y=0 $X2=5.74 $Y2=2.11
cc_135 N_GND_M1016_b N_CK_c_1070_n 0.00654989f $X=-0.05 $Y=0 $X2=3.8 $Y2=2.11
cc_136 N_GND_M1016_b N_CK_c_1071_n 0.0139116f $X=-0.05 $Y=0 $X2=6.735 $Y2=2.11
cc_137 N_GND_M1016_b N_CK_c_1072_n 0.00189466f $X=-0.05 $Y=0 $X2=6.03 $Y2=2.11
cc_138 N_GND_M1016_b CK 0.0014603f $X=-0.05 $Y=0 $X2=6.88 $Y2=2.11
cc_139 N_GND_M1016_b N_A_217_521#_M1020_g 0.0171592f $X=-0.05 $Y=0 $X2=4.555
+ $Y2=0.85
cc_140 N_GND_c_53_p N_A_217_521#_M1020_g 0.00606474f $X=4.685 $Y=0.152 $X2=4.555
+ $Y2=0.85
cc_141 N_GND_c_54_p N_A_217_521#_M1020_g 0.00308284f $X=4.77 $Y=0.74 $X2=4.555
+ $Y2=0.85
cc_142 N_GND_c_5_p N_A_217_521#_M1020_g 0.00468827f $X=9.855 $Y=0.19 $X2=4.555
+ $Y2=0.85
cc_143 N_GND_M1016_b N_A_217_521#_c_1300_n 0.0240372f $X=-0.05 $Y=0 $X2=4.91
+ $Y2=1.4
cc_144 N_GND_c_54_p N_A_217_521#_c_1300_n 9.75298e-19 $X=4.77 $Y=0.74 $X2=4.91
+ $Y2=1.4
cc_145 N_GND_M1016_b N_A_217_521#_c_1302_n 0.0105855f $X=-0.05 $Y=0 $X2=4.63
+ $Y2=1.4
cc_146 N_GND_M1016_b N_A_217_521#_c_1303_n 0.022671f $X=-0.05 $Y=0 $X2=4.91
+ $Y2=2.285
cc_147 N_GND_M1016_b N_A_217_521#_c_1304_n 0.0103324f $X=-0.05 $Y=0 $X2=4.63
+ $Y2=2.285
cc_148 N_GND_M1016_b N_A_217_521#_M1023_g 0.0170177f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=0.85
cc_149 N_GND_c_54_p N_A_217_521#_M1023_g 0.00308284f $X=4.77 $Y=0.74 $X2=4.985
+ $Y2=0.85
cc_150 N_GND_c_55_p N_A_217_521#_M1023_g 0.00606474f $X=6.435 $Y=0.152 $X2=4.985
+ $Y2=0.85
cc_151 N_GND_c_5_p N_A_217_521#_M1023_g 0.00468827f $X=9.855 $Y=0.19 $X2=4.985
+ $Y2=0.85
cc_152 N_GND_M1016_b N_A_217_521#_c_1309_n 0.00545065f $X=-0.05 $Y=0 $X2=1.21
+ $Y2=3.295
cc_153 N_GND_M1016_b N_A_217_521#_c_1310_n 0.00563276f $X=-0.05 $Y=0 $X2=1.565
+ $Y2=1.61
cc_154 N_GND_M1016_b N_A_217_521#_c_1311_n 0.0017406f $X=-0.05 $Y=0 $X2=1.295
+ $Y2=1.61
cc_155 N_GND_M1016_b N_A_217_521#_c_1312_n 0.00531957f $X=-0.05 $Y=0 $X2=1.71
+ $Y2=0.755
cc_156 N_GND_c_13_p N_A_217_521#_c_1312_n 0.00736239f $X=2.415 $Y=0.152 $X2=1.71
+ $Y2=0.755
cc_157 N_GND_c_5_p N_A_217_521#_c_1312_n 0.00476261f $X=9.855 $Y=0.19 $X2=1.71
+ $Y2=0.755
cc_158 N_GND_M1016_b N_A_217_521#_c_1315_n 0.00822335f $X=-0.05 $Y=0 $X2=4.725
+ $Y2=2.285
cc_159 N_GND_M1016_b N_A_217_521#_c_1316_n 0.0033417f $X=-0.05 $Y=0 $X2=1.68
+ $Y2=1.61
cc_160 N_GND_M1016_b N_A_217_521#_c_1317_n 0.00215364f $X=-0.05 $Y=0 $X2=4.725
+ $Y2=1.4
cc_161 N_GND_c_54_p N_A_217_521#_c_1317_n 0.00391768f $X=4.77 $Y=0.74 $X2=4.725
+ $Y2=1.4
cc_162 N_GND_M1016_b N_A_217_521#_c_1319_n 0.0479355f $X=-0.05 $Y=0 $X2=4.49
+ $Y2=1.37
cc_163 N_GND_M1016_b N_A_217_521#_c_1320_n 0.00251249f $X=-0.05 $Y=0 $X2=1.855
+ $Y2=1.37
cc_164 N_GND_M1016_b N_A_704_89#_c_1460_n 0.0156145f $X=-0.05 $Y=0 $X2=3.595
+ $Y2=1.205
cc_165 N_GND_c_53_p N_A_704_89#_c_1460_n 0.00606474f $X=4.685 $Y=0.152 $X2=3.595
+ $Y2=1.205
cc_166 N_GND_c_5_p N_A_704_89#_c_1460_n 0.00468827f $X=9.855 $Y=0.19 $X2=3.595
+ $Y2=1.205
cc_167 N_GND_M1016_b N_A_704_89#_c_1463_n 0.0217592f $X=-0.05 $Y=0 $X2=3.715
+ $Y2=1.775
cc_168 N_GND_M1016_b N_A_704_89#_c_1464_n 0.0182441f $X=-0.05 $Y=0 $X2=4.12
+ $Y2=1.85
cc_169 N_GND_M1016_b N_A_704_89#_c_1465_n 0.00766794f $X=-0.05 $Y=0 $X2=3.79
+ $Y2=1.85
cc_170 N_GND_M1016_b N_A_704_89#_M1014_g 0.0302127f $X=-0.05 $Y=0 $X2=4.195
+ $Y2=3.235
cc_171 N_GND_M1016_b N_A_704_89#_c_1467_n 0.0552247f $X=-0.05 $Y=0 $X2=5.27
+ $Y2=1.85
cc_172 N_GND_M1016_b N_A_704_89#_M1010_g 0.0297952f $X=-0.05 $Y=0 $X2=5.345
+ $Y2=3.235
cc_173 N_GND_M1016_b N_A_704_89#_c_1469_n 0.0182441f $X=-0.05 $Y=0 $X2=5.75
+ $Y2=1.85
cc_174 N_GND_M1016_b N_A_704_89#_M1017_g 0.0327555f $X=-0.05 $Y=0 $X2=5.945
+ $Y2=0.85
cc_175 N_GND_c_55_p N_A_704_89#_M1017_g 0.00606474f $X=6.435 $Y=0.152 $X2=5.945
+ $Y2=0.85
cc_176 N_GND_c_5_p N_A_704_89#_M1017_g 0.00468827f $X=9.855 $Y=0.19 $X2=5.945
+ $Y2=0.85
cc_177 N_GND_M1016_b N_A_704_89#_c_1473_n 0.0143258f $X=-0.05 $Y=0 $X2=3.715
+ $Y2=1.28
cc_178 N_GND_M1016_b N_A_704_89#_c_1474_n 0.00426513f $X=-0.05 $Y=0 $X2=4.195
+ $Y2=1.85
cc_179 N_GND_M1016_b N_A_704_89#_c_1475_n 0.00426513f $X=-0.05 $Y=0 $X2=5.345
+ $Y2=1.85
cc_180 N_GND_M1016_b N_A_704_89#_c_1476_n 0.0292692f $X=-0.05 $Y=0 $X2=5.885
+ $Y2=1.725
cc_181 N_GND_M1016_b N_A_704_89#_c_1477_n 0.00223816f $X=-0.05 $Y=0 $X2=5.885
+ $Y2=1.725
cc_182 N_GND_M1016_b N_A_704_89#_c_1478_n 0.014452f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=0.755
cc_183 N_GND_c_56_p N_A_704_89#_c_1478_n 4.65312e-19 $X=6.52 $Y=0.755 $X2=6.95
+ $Y2=0.755
cc_184 N_GND_c_57_p N_A_704_89#_c_1478_n 0.0074445f $X=7.385 $Y=0.152 $X2=6.95
+ $Y2=0.755
cc_185 N_GND_c_58_p N_A_704_89#_c_1478_n 0.0151608f $X=7.47 $Y=0.755 $X2=6.95
+ $Y2=0.755
cc_186 N_GND_c_5_p N_A_704_89#_c_1478_n 0.00476261f $X=9.855 $Y=0.19 $X2=6.95
+ $Y2=0.755
cc_187 N_GND_M1016_b N_A_704_89#_c_1483_n 0.0102727f $X=-0.05 $Y=0 $X2=7.22
+ $Y2=2.62
cc_188 N_GND_M1016_b N_A_704_89#_c_1484_n 0.0100174f $X=-0.05 $Y=0 $X2=7.22
+ $Y2=1.717
cc_189 N_GND_M1016_b N_A_704_89#_c_1485_n 0.00652814f $X=-0.05 $Y=0 $X2=6.835
+ $Y2=1.725
cc_190 N_GND_M1016_b N_A_704_89#_c_1486_n 0.00244571f $X=-0.05 $Y=0 $X2=6.05
+ $Y2=1.725
cc_191 N_GND_M1016_b N_A_704_89#_c_1487_n 0.00234408f $X=-0.05 $Y=0 $X2=6.95
+ $Y2=1.725
cc_192 N_GND_M1016_b N_A_1246_89#_M1006_g 0.0305867f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=0.85
cc_193 N_GND_c_55_p N_A_1246_89#_M1006_g 0.00606474f $X=6.435 $Y=0.152 $X2=6.305
+ $Y2=0.85
cc_194 N_GND_c_56_p N_A_1246_89#_M1006_g 0.00315235f $X=6.52 $Y=0.755 $X2=6.305
+ $Y2=0.85
cc_195 N_GND_c_5_p N_A_1246_89#_M1006_g 0.00468827f $X=9.855 $Y=0.19 $X2=6.305
+ $Y2=0.85
cc_196 N_GND_M1016_b N_A_1246_89#_M1029_g 0.0301968f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=3.235
cc_197 N_GND_M1016_b N_A_1246_89#_c_1677_n 0.0259391f $X=-0.05 $Y=0 $X2=6.365
+ $Y2=1.71
cc_198 N_GND_c_56_p N_A_1246_89#_c_1677_n 0.00109087f $X=6.52 $Y=0.755 $X2=6.365
+ $Y2=1.71
cc_199 N_GND_M1016_b N_A_1246_89#_c_1679_n 0.0270403f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=1.71
cc_200 N_GND_M1016_b N_A_1246_89#_c_1680_n 0.00921847f $X=-0.05 $Y=0 $X2=9.382
+ $Y2=1.545
cc_201 N_GND_M1016_b N_A_1246_89#_c_1681_n 0.0183502f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=1.23
cc_202 N_GND_c_17_p N_A_1246_89#_c_1681_n 0.0035726f $X=8.75 $Y=0.74 $X2=9.47
+ $Y2=1.23
cc_203 N_GND_c_61_p N_A_1246_89#_c_1681_n 0.00606474f $X=9.625 $Y=0.152 $X2=9.47
+ $Y2=1.23
cc_204 N_GND_c_204_p N_A_1246_89#_c_1681_n 0.00308284f $X=9.71 $Y=0.755 $X2=9.47
+ $Y2=1.23
cc_205 N_GND_c_5_p N_A_1246_89#_c_1681_n 0.00468827f $X=9.855 $Y=0.19 $X2=9.47
+ $Y2=1.23
cc_206 N_GND_M1016_b N_A_1246_89#_c_1686_n 0.0125076f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=1.38
cc_207 N_GND_M1016_b N_A_1246_89#_c_1687_n 0.0284927f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=2.375
cc_208 N_GND_M1016_b N_A_1246_89#_c_1688_n 0.00455162f $X=-0.05 $Y=0 $X2=9.47
+ $Y2=2.525
cc_209 N_GND_M1016_b N_A_1246_89#_c_1689_n 0.00491423f $X=-0.05 $Y=0 $X2=6.365
+ $Y2=1.71
cc_210 N_GND_M1016_b N_A_1246_89#_c_1690_n 0.00601598f $X=-0.05 $Y=0 $X2=8.26
+ $Y2=0.755
cc_211 N_GND_c_16_p N_A_1246_89#_c_1690_n 0.00750865f $X=8.665 $Y=0.152 $X2=8.26
+ $Y2=0.755
cc_212 N_GND_c_5_p N_A_1246_89#_c_1690_n 0.00476261f $X=9.855 $Y=0.19 $X2=8.26
+ $Y2=0.755
cc_213 N_GND_M1016_b N_A_1246_89#_c_1693_n 0.00495979f $X=-0.05 $Y=0 $X2=8.76
+ $Y2=3.295
cc_214 N_GND_M1016_b N_A_1246_89#_c_1694_n 0.0197717f $X=-0.05 $Y=0 $X2=8.845
+ $Y2=1.71
cc_215 N_GND_M1016_b N_A_1246_89#_c_1695_n 0.00907353f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=1.71
cc_216 N_GND_M1016_b N_A_1246_89#_c_1696_n 0.00254619f $X=-0.05 $Y=0 $X2=7.165
+ $Y2=2.482
cc_217 N_GND_M1016_b N_A_1246_89#_c_1697_n 0.00392233f $X=-0.05 $Y=0 $X2=7.305
+ $Y2=2.39
cc_218 N_GND_M1016_b N_A_1246_89#_c_1698_n 0.0436125f $X=-0.05 $Y=0 $X2=9.235
+ $Y2=1.71
cc_219 N_GND_M1016_b N_A_1246_89#_c_1699_n 0.00111647f $X=-0.05 $Y=0 $X2=7.375
+ $Y2=1.71
cc_220 N_GND_M1016_b N_A_1246_89#_c_1700_n 0.00129525f $X=-0.05 $Y=0 $X2=6.515
+ $Y2=2.48
cc_221 N_GND_M1016_b N_A_1246_89#_c_1701_n 0.0014645f $X=-0.05 $Y=0 $X2=9.38
+ $Y2=1.71
cc_222 N_GND_M1016_b N_A_1084_115#_c_1883_n 0.0449791f $X=-0.05 $Y=0 $X2=7.505
+ $Y2=2.15
cc_223 N_GND_M1016_b N_A_1084_115#_c_1884_n 0.0160302f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.21
cc_224 N_GND_c_58_p N_A_1084_115#_c_1884_n 0.00509667f $X=7.47 $Y=0.755
+ $X2=7.685 $Y2=1.21
cc_225 N_GND_c_16_p N_A_1084_115#_c_1884_n 0.00606474f $X=8.665 $Y=0.152
+ $X2=7.685 $Y2=1.21
cc_226 N_GND_c_5_p N_A_1084_115#_c_1884_n 0.00468827f $X=9.855 $Y=0.19 $X2=7.685
+ $Y2=1.21
cc_227 N_GND_M1016_b N_A_1084_115#_c_1888_n 0.0235095f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.29
cc_228 N_GND_c_58_p N_A_1084_115#_c_1888_n 0.00391038f $X=7.47 $Y=0.755
+ $X2=7.685 $Y2=1.29
cc_229 N_GND_M1016_b N_A_1084_115#_c_1890_n 0.0329441f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=2.285
cc_230 N_GND_M1016_b N_A_1084_115#_c_1891_n 0.0108511f $X=-0.05 $Y=0 $X2=5.065
+ $Y2=1.37
cc_231 N_GND_M1016_b N_A_1084_115#_c_1892_n 0.00800183f $X=-0.05 $Y=0 $X2=5.745
+ $Y2=1.34
cc_232 N_GND_M1016_b N_A_1084_115#_c_1893_n 0.00561499f $X=-0.05 $Y=0 $X2=7.595
+ $Y2=1.37
cc_233 N_GND_c_58_p N_A_1084_115#_c_1893_n 0.00131024f $X=7.47 $Y=0.755
+ $X2=7.595 $Y2=1.37
cc_234 N_GND_M1016_b N_A_1084_115#_c_1895_n 0.00312748f $X=-0.05 $Y=0 $X2=5.645
+ $Y2=0.755
cc_235 N_GND_c_55_p N_A_1084_115#_c_1895_n 0.0150277f $X=6.435 $Y=0.152
+ $X2=5.645 $Y2=0.755
cc_236 N_GND_c_5_p N_A_1084_115#_c_1895_n 0.00994746f $X=9.855 $Y=0.19 $X2=5.645
+ $Y2=0.755
cc_237 N_GND_M1016_b N_A_1084_115#_c_1898_n 0.00227051f $X=-0.05 $Y=0 $X2=5.6
+ $Y2=1.37
cc_238 N_GND_M1016_b N_A_1084_115#_c_1899_n 0.00135835f $X=-0.05 $Y=0 $X2=5.21
+ $Y2=1.37
cc_239 N_GND_M1016_b N_A_1084_115#_c_1900_n 0.0141417f $X=-0.05 $Y=0 $X2=7.45
+ $Y2=1.37
cc_240 N_GND_c_56_p N_A_1084_115#_c_1900_n 8.35925e-19 $X=6.52 $Y=0.755 $X2=7.45
+ $Y2=1.37
cc_241 N_GND_c_58_p N_A_1084_115#_c_1900_n 3.1624e-19 $X=7.47 $Y=0.755 $X2=7.45
+ $Y2=1.37
cc_242 N_GND_M1016_b N_A_1084_115#_c_1903_n 0.00325484f $X=-0.05 $Y=0 $X2=5.89
+ $Y2=1.37
cc_243 N_GND_M1016_b N_A_1084_115#_c_1904_n 0.00169121f $X=-0.05 $Y=0 $X2=7.595
+ $Y2=1.37
cc_244 N_GND_c_58_p N_A_1084_115#_c_1904_n 4.00959e-19 $X=7.47 $Y=0.755
+ $X2=7.595 $Y2=1.37
cc_245 N_GND_M1016_b N_QN_M1008_g 0.0543664f $X=-0.05 $Y=0 $X2=9.925 $Y2=0.85
cc_246 N_GND_c_204_p N_QN_M1008_g 0.00308284f $X=9.71 $Y=0.755 $X2=9.925
+ $Y2=0.85
cc_247 N_GND_c_5_p N_QN_M1008_g 0.00468827f $X=9.855 $Y=0.19 $X2=9.925 $Y2=0.85
cc_248 N_GND_M1016_b N_QN_M1032_g 0.0186095f $X=-0.05 $Y=0 $X2=9.925 $Y2=3.235
cc_249 N_GND_M1016_b N_QN_c_2064_n 0.0291912f $X=-0.05 $Y=0 $X2=9.865 $Y2=1.915
cc_250 N_GND_M1016_b N_QN_c_2065_n 0.00370057f $X=-0.05 $Y=0 $X2=9.28 $Y2=0.755
cc_251 N_GND_c_17_p N_QN_c_2065_n 0.013807f $X=8.75 $Y=0.74 $X2=9.28 $Y2=0.755
cc_252 N_GND_c_61_p N_QN_c_2065_n 0.00736239f $X=9.625 $Y=0.152 $X2=9.28
+ $Y2=0.755
cc_253 N_GND_c_5_p N_QN_c_2065_n 0.00476261f $X=9.855 $Y=0.19 $X2=9.28 $Y2=0.755
cc_254 N_GND_M1016_b N_QN_c_2069_n 0.00102655f $X=-0.05 $Y=0 $X2=9.28 $Y2=2.48
cc_255 N_GND_M1016_b N_QN_c_2070_n 0.0133445f $X=-0.05 $Y=0 $X2=9.78 $Y2=1.37
cc_256 N_GND_c_204_p N_QN_c_2070_n 0.00827206f $X=9.71 $Y=0.755 $X2=9.78
+ $Y2=1.37
cc_257 N_GND_M1016_b N_QN_c_2072_n 0.00188316f $X=-0.05 $Y=0 $X2=9.365 $Y2=1.37
cc_258 N_GND_M1016_b N_QN_c_2073_n 0.0138424f $X=-0.05 $Y=0 $X2=9.78 $Y2=2.285
cc_259 N_GND_M1016_b N_QN_c_2074_n 0.00301984f $X=-0.05 $Y=0 $X2=9.365 $Y2=2.285
cc_260 N_GND_M1016_b N_QN_c_2075_n 0.0034889f $X=-0.05 $Y=0 $X2=9.865 $Y2=1.915
cc_261 N_GND_M1016_b QN 0.00258296f $X=-0.05 $Y=0 $X2=9.285 $Y2=2.48
cc_262 N_GND_M1016_b N_Q_c_2191_n 0.00880132f $X=-0.05 $Y=0 $X2=10.14 $Y2=0.755
cc_263 N_GND_c_5_p N_Q_c_2191_n 0.00467398f $X=9.855 $Y=0.19 $X2=10.14 $Y2=0.755
cc_264 N_GND_M1016_b N_Q_c_2193_n 0.0622366f $X=-0.05 $Y=0 $X2=10.255 $Y2=2.525
cc_265 N_GND_M1016_b N_Q_c_2194_n 0.0106402f $X=-0.05 $Y=0 $X2=10.255 $Y2=1.035
cc_266 N_VDD_M1001_b N_RN_M1001_g 0.0269777f $X=-0.05 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_267 N_VDD_c_267_p N_RN_M1001_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_268 N_VDD_c_268_p N_RN_M1001_g 0.00606474f $X=1.985 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_269 N_VDD_c_269_p N_RN_M1001_g 0.00468827f $X=9.855 $Y=4.25 $X2=0.475
+ $Y2=3.235
cc_270 N_VDD_M1001_s N_RN_c_438_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32
+ $Y2=2.85
cc_271 N_VDD_M1001_b N_RN_c_438_n 0.00618364f $X=-0.05 $Y=2.425 $X2=0.32
+ $Y2=2.85
cc_272 N_VDD_c_267_p N_RN_c_438_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_273 N_VDD_M1001_s RN 0.0162774f $X=0.135 $Y=2.605 $X2=0.325 $Y2=2.85
cc_274 N_VDD_c_267_p RN 0.00522047f $X=0.26 $Y=3.635 $X2=0.325 $Y2=2.85
cc_275 N_VDD_M1001_b N_A_110_115#_M1000_g 0.022052f $X=-0.05 $Y=2.425 $X2=1.425
+ $Y2=3.235
cc_276 N_VDD_c_268_p N_A_110_115#_M1000_g 0.00606474f $X=1.985 $Y=4.287
+ $X2=1.425 $Y2=3.235
cc_277 N_VDD_c_269_p N_A_110_115#_M1000_g 0.00468827f $X=9.855 $Y=4.25 $X2=1.425
+ $Y2=3.235
cc_278 N_VDD_M1001_b N_A_110_115#_M1025_g 0.0246741f $X=-0.05 $Y=2.425 $X2=8.545
+ $Y2=3.235
cc_279 N_VDD_c_279_p N_A_110_115#_M1025_g 0.00606474f $X=9.625 $Y=4.287
+ $X2=8.545 $Y2=3.235
cc_280 N_VDD_c_269_p N_A_110_115#_M1025_g 0.00468827f $X=9.855 $Y=4.25 $X2=8.545
+ $Y2=3.235
cc_281 N_VDD_M1001_b N_A_110_115#_c_484_n 0.00862296f $X=-0.05 $Y=2.425
+ $X2=1.425 $Y2=2.395
cc_282 N_VDD_M1001_b N_A_110_115#_c_494_n 0.00546889f $X=-0.05 $Y=2.425 $X2=0.69
+ $Y2=2.955
cc_283 N_VDD_c_268_p N_A_110_115#_c_494_n 0.00757793f $X=1.985 $Y=4.287 $X2=0.69
+ $Y2=2.955
cc_284 N_VDD_c_269_p N_A_110_115#_c_494_n 0.00476261f $X=9.855 $Y=4.25 $X2=0.69
+ $Y2=2.955
cc_285 N_VDD_M1001_b N_SN_M1024_g 0.0195253f $X=-0.05 $Y=2.425 $X2=1.855
+ $Y2=3.235
cc_286 N_VDD_c_268_p N_SN_M1024_g 0.00606474f $X=1.985 $Y=4.287 $X2=1.855
+ $Y2=3.235
cc_287 N_VDD_c_287_p N_SN_M1024_g 0.00308284f $X=2.07 $Y=3.7 $X2=1.855 $Y2=3.235
cc_288 N_VDD_c_269_p N_SN_M1024_g 0.00468827f $X=9.855 $Y=4.25 $X2=1.855
+ $Y2=3.235
cc_289 N_VDD_M1001_b N_SN_M1019_g 0.0205652f $X=-0.05 $Y=2.425 $X2=8.115
+ $Y2=3.235
cc_290 N_VDD_c_290_p N_SN_M1019_g 0.00308284f $X=7.9 $Y=3.7 $X2=8.115 $Y2=3.235
cc_291 N_VDD_c_279_p N_SN_M1019_g 0.00606474f $X=9.625 $Y=4.287 $X2=8.115
+ $Y2=3.235
cc_292 N_VDD_c_269_p N_SN_M1019_g 0.00468827f $X=9.855 $Y=4.25 $X2=8.115
+ $Y2=3.235
cc_293 N_VDD_M1001_b N_SN_c_715_n 0.00132936f $X=-0.05 $Y=2.425 $X2=1.71
+ $Y2=2.62
cc_294 N_VDD_M1001_b N_SN_c_716_n 0.00126532f $X=-0.05 $Y=2.425 $X2=7.937
+ $Y2=2.482
cc_295 N_VDD_M1033_d N_SN_c_730_n 0.00754969f $X=7.76 $Y=2.605 $X2=7.935
+ $Y2=2.845
cc_296 N_VDD_M1001_b N_SN_c_730_n 0.00286365f $X=-0.05 $Y=2.425 $X2=7.935
+ $Y2=2.845
cc_297 N_VDD_M1024_d N_SN_c_732_n 0.0118947f $X=1.93 $Y=2.605 $X2=1.71 $Y2=2.777
cc_298 N_VDD_M1024_d N_SN_c_733_n 3.46903e-19 $X=1.93 $Y=2.605 $X2=7.79 $Y2=2.85
cc_299 N_VDD_M1028_s N_SN_c_733_n 0.00517585f $X=2.895 $Y=2.605 $X2=7.79
+ $Y2=2.85
cc_300 N_VDD_M1009_d N_SN_c_733_n 0.0113422f $X=4.63 $Y=2.605 $X2=7.79 $Y2=2.85
cc_301 N_VDD_M1029_d N_SN_c_733_n 0.0063778f $X=6.38 $Y=2.605 $X2=7.79 $Y2=2.85
cc_302 N_VDD_M1033_d N_SN_c_733_n 0.00135552f $X=7.76 $Y=2.605 $X2=7.79 $Y2=2.85
cc_303 N_VDD_M1001_b N_SN_c_733_n 0.0209311f $X=-0.05 $Y=2.425 $X2=7.79 $Y2=2.85
cc_304 N_VDD_c_304_p N_SN_c_733_n 0.00512495f $X=3.02 $Y=3.295 $X2=7.79 $Y2=2.85
cc_305 N_VDD_c_305_p N_SN_c_733_n 0.00697427f $X=4.77 $Y=3.295 $X2=7.79 $Y2=2.85
cc_306 N_VDD_c_306_p N_SN_c_733_n 0.0152728f $X=6.52 $Y=3.21 $X2=7.79 $Y2=2.85
cc_307 N_VDD_M1024_d N_SN_c_742_n 0.00440365f $X=1.93 $Y=2.605 $X2=2.195
+ $Y2=2.85
cc_308 N_VDD_M1033_d SN 0.00692874f $X=7.76 $Y=2.605 $X2=7.94 $Y2=2.845
cc_309 N_VDD_M1001_b N_A_432_424#_M1027_g 0.0214531f $X=-0.05 $Y=2.425 $X2=2.285
+ $Y2=3.235
cc_310 N_VDD_c_287_p N_A_432_424#_M1027_g 0.00308284f $X=2.07 $Y=3.7 $X2=2.285
+ $Y2=3.235
cc_311 N_VDD_c_311_p N_A_432_424#_M1027_g 0.00606474f $X=2.935 $Y=4.287
+ $X2=2.285 $Y2=3.235
cc_312 N_VDD_c_304_p N_A_432_424#_M1027_g 0.0041296f $X=3.02 $Y=3.295 $X2=2.285
+ $Y2=3.235
cc_313 N_VDD_c_269_p N_A_432_424#_M1027_g 0.00468827f $X=9.855 $Y=4.25 $X2=2.285
+ $Y2=3.235
cc_314 N_VDD_M1001_b N_A_432_424#_c_900_n 0.00572f $X=-0.05 $Y=2.425 $X2=2.295
+ $Y2=2.285
cc_315 N_VDD_M1001_b N_A_432_424#_c_901_n 2.73199e-19 $X=-0.05 $Y=2.425
+ $X2=2.295 $Y2=2.2
cc_316 N_VDD_M1001_b N_A_432_424#_c_907_n 0.00527983f $X=-0.05 $Y=2.425 $X2=2.77
+ $Y2=2.62
cc_317 N_VDD_M1028_s N_A_432_424#_c_920_n 0.0106534f $X=2.895 $Y=2.605 $X2=3.725
+ $Y2=2.705
cc_318 N_VDD_M1001_b N_A_432_424#_c_920_n 0.00208149f $X=-0.05 $Y=2.425
+ $X2=3.725 $Y2=2.705
cc_319 N_VDD_c_304_p N_A_432_424#_c_920_n 0.00682058f $X=3.02 $Y=3.295 $X2=3.725
+ $Y2=2.705
cc_320 N_VDD_M1001_b N_A_432_424#_c_923_n 0.00504431f $X=-0.05 $Y=2.425
+ $X2=2.855 $Y2=2.705
cc_321 N_VDD_M1001_b N_A_432_424#_c_924_n 0.00313975f $X=-0.05 $Y=2.425
+ $X2=3.895 $Y2=2.955
cc_322 N_VDD_c_322_p N_A_432_424#_c_924_n 0.0149718f $X=4.685 $Y=4.287 $X2=3.895
+ $Y2=2.955
cc_323 N_VDD_c_269_p N_A_432_424#_c_924_n 0.00958198f $X=9.855 $Y=4.25 $X2=3.895
+ $Y2=2.955
cc_324 N_VDD_M1001_b N_D_M1028_g 0.0210334f $X=-0.05 $Y=2.425 $X2=3.235
+ $Y2=3.235
cc_325 N_VDD_c_304_p N_D_M1028_g 0.00636672f $X=3.02 $Y=3.295 $X2=3.235
+ $Y2=3.235
cc_326 N_VDD_c_322_p N_D_M1028_g 0.00606474f $X=4.685 $Y=4.287 $X2=3.235
+ $Y2=3.235
cc_327 N_VDD_c_269_p N_D_M1028_g 0.00468827f $X=9.855 $Y=4.25 $X2=3.235
+ $Y2=3.235
cc_328 N_VDD_M1001_b N_CK_M1018_g 0.0201271f $X=-0.05 $Y=2.425 $X2=3.595
+ $Y2=3.235
cc_329 N_VDD_c_322_p N_CK_M1018_g 0.00606474f $X=4.685 $Y=4.287 $X2=3.595
+ $Y2=3.235
cc_330 N_VDD_c_269_p N_CK_M1018_g 0.00468827f $X=9.855 $Y=4.25 $X2=3.595
+ $Y2=3.235
cc_331 N_VDD_M1001_b N_CK_M1002_g 0.0201163f $X=-0.05 $Y=2.425 $X2=5.945
+ $Y2=3.235
cc_332 N_VDD_c_332_p N_CK_M1002_g 0.00606474f $X=6.435 $Y=4.287 $X2=5.945
+ $Y2=3.235
cc_333 N_VDD_c_269_p N_CK_M1002_g 0.00468827f $X=9.855 $Y=4.25 $X2=5.945
+ $Y2=3.235
cc_334 N_VDD_M1001_b N_CK_c_1043_n 0.007968f $X=-0.05 $Y=2.425 $X2=6.735
+ $Y2=2.45
cc_335 N_VDD_M1001_b N_CK_M1031_g 0.0241582f $X=-0.05 $Y=2.425 $X2=6.735
+ $Y2=3.235
cc_336 N_VDD_c_306_p N_CK_M1031_g 0.00413862f $X=6.52 $Y=3.21 $X2=6.735
+ $Y2=3.235
cc_337 N_VDD_c_337_p N_CK_M1031_g 0.00606474f $X=7.815 $Y=4.287 $X2=6.735
+ $Y2=3.235
cc_338 N_VDD_c_269_p N_CK_M1031_g 0.00468827f $X=9.855 $Y=4.25 $X2=6.735
+ $Y2=3.235
cc_339 N_VDD_M1001_b N_CK_c_1045_n 0.00654707f $X=-0.05 $Y=2.425 $X2=3.685
+ $Y2=2.285
cc_340 N_VDD_M1001_b N_CK_c_1054_n 0.00654388f $X=-0.05 $Y=2.425 $X2=5.855
+ $Y2=2.285
cc_341 N_VDD_M1001_b N_CK_c_1066_n 0.0010436f $X=-0.05 $Y=2.425 $X2=6.88
+ $Y2=2.11
cc_342 N_VDD_M1001_b N_CK_c_1067_n 8.09007e-19 $X=-0.05 $Y=2.425 $X2=3.655
+ $Y2=2.11
cc_343 N_VDD_M1001_b N_CK_c_1068_n 0.00115766f $X=-0.05 $Y=2.425 $X2=5.885
+ $Y2=2.11
cc_344 N_VDD_M1001_b N_A_217_521#_M1009_g 0.0192219f $X=-0.05 $Y=2.425 $X2=4.555
+ $Y2=3.235
cc_345 N_VDD_c_322_p N_A_217_521#_M1009_g 0.00606474f $X=4.685 $Y=4.287
+ $X2=4.555 $Y2=3.235
cc_346 N_VDD_c_305_p N_A_217_521#_M1009_g 0.00337744f $X=4.77 $Y=3.295 $X2=4.555
+ $Y2=3.235
cc_347 N_VDD_c_269_p N_A_217_521#_M1009_g 0.00468827f $X=9.855 $Y=4.25 $X2=4.555
+ $Y2=3.235
cc_348 N_VDD_c_305_p N_A_217_521#_c_1303_n 8.24975e-19 $X=4.77 $Y=3.295 $X2=4.91
+ $Y2=2.285
cc_349 N_VDD_M1001_b N_A_217_521#_M1012_g 0.0181098f $X=-0.05 $Y=2.425 $X2=4.985
+ $Y2=3.235
cc_350 N_VDD_c_305_p N_A_217_521#_M1012_g 0.00337744f $X=4.77 $Y=3.295 $X2=4.985
+ $Y2=3.235
cc_351 N_VDD_c_332_p N_A_217_521#_M1012_g 0.00606474f $X=6.435 $Y=4.287
+ $X2=4.985 $Y2=3.235
cc_352 N_VDD_c_269_p N_A_217_521#_M1012_g 0.00468827f $X=9.855 $Y=4.25 $X2=4.985
+ $Y2=3.235
cc_353 N_VDD_M1001_b N_A_217_521#_c_1309_n 0.00426107f $X=-0.05 $Y=2.425
+ $X2=1.21 $Y2=3.295
cc_354 N_VDD_c_268_p N_A_217_521#_c_1309_n 0.00745733f $X=1.985 $Y=4.287
+ $X2=1.21 $Y2=3.295
cc_355 N_VDD_c_269_p N_A_217_521#_c_1309_n 0.00476261f $X=9.855 $Y=4.25 $X2=1.21
+ $Y2=3.295
cc_356 N_VDD_M1001_b N_A_217_521#_c_1315_n 0.00269632f $X=-0.05 $Y=2.425
+ $X2=4.725 $Y2=2.285
cc_357 N_VDD_c_305_p N_A_217_521#_c_1315_n 0.00176301f $X=4.77 $Y=3.295
+ $X2=4.725 $Y2=2.285
cc_358 N_VDD_M1001_b N_A_704_89#_M1014_g 0.0214581f $X=-0.05 $Y=2.425 $X2=4.195
+ $Y2=3.235
cc_359 N_VDD_c_322_p N_A_704_89#_M1014_g 0.00606474f $X=4.685 $Y=4.287 $X2=4.195
+ $Y2=3.235
cc_360 N_VDD_c_269_p N_A_704_89#_M1014_g 0.00468827f $X=9.855 $Y=4.25 $X2=4.195
+ $Y2=3.235
cc_361 N_VDD_M1001_b N_A_704_89#_M1010_g 0.0214271f $X=-0.05 $Y=2.425 $X2=5.345
+ $Y2=3.235
cc_362 N_VDD_c_332_p N_A_704_89#_M1010_g 0.00606474f $X=6.435 $Y=4.287 $X2=5.345
+ $Y2=3.235
cc_363 N_VDD_c_269_p N_A_704_89#_M1010_g 0.00468827f $X=9.855 $Y=4.25 $X2=5.345
+ $Y2=3.235
cc_364 N_VDD_M1001_b N_A_704_89#_c_1494_n 0.00156053f $X=-0.05 $Y=2.425 $X2=6.95
+ $Y2=2.955
cc_365 N_VDD_c_306_p N_A_704_89#_c_1494_n 9.30625e-19 $X=6.52 $Y=3.21 $X2=6.95
+ $Y2=2.955
cc_366 N_VDD_c_337_p N_A_704_89#_c_1494_n 0.0074445f $X=7.815 $Y=4.287 $X2=6.95
+ $Y2=2.955
cc_367 N_VDD_c_269_p N_A_704_89#_c_1494_n 0.00476261f $X=9.855 $Y=4.25 $X2=6.95
+ $Y2=2.955
cc_368 N_VDD_M1001_b N_A_704_89#_c_1483_n 0.00531414f $X=-0.05 $Y=2.425 $X2=7.22
+ $Y2=2.62
cc_369 N_VDD_M1001_b N_A_704_89#_c_1499_n 0.00687104f $X=-0.05 $Y=2.425 $X2=7.22
+ $Y2=2.705
cc_370 N_VDD_M1001_b N_A_1246_89#_M1029_g 0.0178558f $X=-0.05 $Y=2.425 $X2=6.305
+ $Y2=3.235
cc_371 N_VDD_c_332_p N_A_1246_89#_M1029_g 0.00606474f $X=6.435 $Y=4.287
+ $X2=6.305 $Y2=3.235
cc_372 N_VDD_c_306_p N_A_1246_89#_M1029_g 0.00421098f $X=6.52 $Y=3.21 $X2=6.305
+ $Y2=3.235
cc_373 N_VDD_c_269_p N_A_1246_89#_M1029_g 0.00468827f $X=9.855 $Y=4.25 $X2=6.305
+ $Y2=3.235
cc_374 N_VDD_M1001_b N_A_1246_89#_c_1688_n 0.0289507f $X=-0.05 $Y=2.425 $X2=9.47
+ $Y2=2.525
cc_375 N_VDD_c_279_p N_A_1246_89#_c_1688_n 0.00606474f $X=9.625 $Y=4.287
+ $X2=9.47 $Y2=2.525
cc_376 N_VDD_c_376_p N_A_1246_89#_c_1688_n 0.00337744f $X=9.71 $Y=2.955 $X2=9.47
+ $Y2=2.525
cc_377 N_VDD_c_269_p N_A_1246_89#_c_1688_n 0.00468827f $X=9.855 $Y=4.25 $X2=9.47
+ $Y2=2.525
cc_378 N_VDD_M1001_b N_A_1246_89#_c_1689_n 0.00242843f $X=-0.05 $Y=2.425
+ $X2=6.365 $Y2=1.71
cc_379 N_VDD_c_306_p N_A_1246_89#_c_1689_n 4.80241e-19 $X=6.52 $Y=3.21 $X2=6.365
+ $Y2=1.71
cc_380 N_VDD_M1001_b N_A_1246_89#_c_1693_n 0.00467454f $X=-0.05 $Y=2.425
+ $X2=8.76 $Y2=3.295
cc_381 N_VDD_c_279_p N_A_1246_89#_c_1693_n 0.00754714f $X=9.625 $Y=4.287
+ $X2=8.76 $Y2=3.295
cc_382 N_VDD_c_269_p N_A_1246_89#_c_1693_n 0.00476261f $X=9.855 $Y=4.25 $X2=8.76
+ $Y2=3.295
cc_383 N_VDD_M1001_b N_A_1246_89#_c_1696_n 0.00441981f $X=-0.05 $Y=2.425
+ $X2=7.165 $Y2=2.482
cc_384 N_VDD_c_306_p N_A_1246_89#_c_1696_n 4.71502e-19 $X=6.52 $Y=3.21 $X2=7.165
+ $Y2=2.482
cc_385 N_VDD_M1001_b N_A_1246_89#_c_1700_n 0.00375232f $X=-0.05 $Y=2.425
+ $X2=6.515 $Y2=2.48
cc_386 N_VDD_c_306_p N_A_1246_89#_c_1700_n 3.96997e-19 $X=6.52 $Y=3.21 $X2=6.515
+ $Y2=2.48
cc_387 N_VDD_M1001_b N_A_1084_115#_M1033_g 0.025099f $X=-0.05 $Y=2.425 $X2=7.685
+ $Y2=3.235
cc_388 N_VDD_c_337_p N_A_1084_115#_M1033_g 0.00606474f $X=7.815 $Y=4.287
+ $X2=7.685 $Y2=3.235
cc_389 N_VDD_c_290_p N_A_1084_115#_M1033_g 0.00308284f $X=7.9 $Y=3.7 $X2=7.685
+ $Y2=3.235
cc_390 N_VDD_c_269_p N_A_1084_115#_M1033_g 0.00468827f $X=9.855 $Y=4.25
+ $X2=7.685 $Y2=3.235
cc_391 N_VDD_M1001_b N_A_1084_115#_c_1891_n 0.00167876f $X=-0.05 $Y=2.425
+ $X2=5.065 $Y2=1.37
cc_392 N_VDD_M1001_b N_A_1084_115#_c_1911_n 0.00313975f $X=-0.05 $Y=2.425
+ $X2=5.645 $Y2=3.295
cc_393 N_VDD_c_332_p N_A_1084_115#_c_1911_n 0.0149333f $X=6.435 $Y=4.287
+ $X2=5.645 $Y2=3.295
cc_394 N_VDD_c_306_p N_A_1084_115#_c_1911_n 3.30052e-19 $X=6.52 $Y=3.21
+ $X2=5.645 $Y2=3.295
cc_395 N_VDD_c_269_p N_A_1084_115#_c_1911_n 0.00958198f $X=9.855 $Y=4.25
+ $X2=5.645 $Y2=3.295
cc_396 N_VDD_M1001_b N_A_1084_115#_c_1893_n 0.00148487f $X=-0.05 $Y=2.425
+ $X2=7.595 $Y2=1.37
cc_397 N_VDD_M1001_b N_QN_M1032_g 0.0247184f $X=-0.05 $Y=2.425 $X2=9.925
+ $Y2=3.235
cc_398 N_VDD_c_376_p N_QN_M1032_g 0.00337744f $X=9.71 $Y=2.955 $X2=9.925
+ $Y2=3.235
cc_399 N_VDD_c_399_p N_QN_M1032_g 0.00606474f $X=9.855 $Y=4.22 $X2=9.925
+ $Y2=3.235
cc_400 N_VDD_c_269_p N_QN_M1032_g 0.00468827f $X=9.855 $Y=4.25 $X2=9.925
+ $Y2=3.235
cc_401 N_VDD_M1001_b N_QN_c_2069_n 0.00531805f $X=-0.05 $Y=2.425 $X2=9.28
+ $Y2=2.48
cc_402 N_VDD_c_279_p N_QN_c_2069_n 0.00736239f $X=9.625 $Y=4.287 $X2=9.28
+ $Y2=2.48
cc_403 N_VDD_c_269_p N_QN_c_2069_n 0.00476261f $X=9.855 $Y=4.25 $X2=9.28
+ $Y2=2.48
cc_404 N_VDD_c_376_p N_QN_c_2073_n 0.00818856f $X=9.71 $Y=2.955 $X2=9.78
+ $Y2=2.285
cc_405 N_VDD_M1001_b QN 0.0101088f $X=-0.05 $Y=2.425 $X2=9.285 $Y2=2.48
cc_406 N_VDD_M1001_b N_A_300_521#_c_2143_n 0.00155118f $X=-0.05 $Y=2.425
+ $X2=1.64 $Y2=3.295
cc_407 N_VDD_c_268_p N_A_300_521#_c_2143_n 0.00734006f $X=1.985 $Y=4.287
+ $X2=1.64 $Y2=3.295
cc_408 N_VDD_c_269_p N_A_300_521#_c_2143_n 0.00475776f $X=9.855 $Y=4.25 $X2=1.64
+ $Y2=3.295
cc_409 N_VDD_M1024_d N_A_300_521#_c_2146_n 0.00376542f $X=1.93 $Y=2.605
+ $X2=2.415 $Y2=3.19
cc_410 N_VDD_c_287_p N_A_300_521#_c_2146_n 0.0090579f $X=2.07 $Y=3.7 $X2=2.415
+ $Y2=3.19
cc_411 N_VDD_c_304_p N_A_300_521#_c_2146_n 0.00982979f $X=3.02 $Y=3.295
+ $X2=2.415 $Y2=3.19
cc_412 N_VDD_M1001_b N_A_300_521#_c_2149_n 0.00156053f $X=-0.05 $Y=2.425 $X2=2.5
+ $Y2=3.295
cc_413 N_VDD_c_311_p N_A_300_521#_c_2149_n 0.00736752f $X=2.935 $Y=4.287 $X2=2.5
+ $Y2=3.295
cc_414 N_VDD_c_304_p N_A_300_521#_c_2149_n 0.0251825f $X=3.02 $Y=3.295 $X2=2.5
+ $Y2=3.295
cc_415 N_VDD_c_269_p N_A_300_521#_c_2149_n 0.00476261f $X=9.855 $Y=4.25 $X2=2.5
+ $Y2=3.295
cc_416 N_VDD_M1001_b N_A_1469_521#_c_2171_n 0.00156053f $X=-0.05 $Y=2.425
+ $X2=7.47 $Y2=3.295
cc_417 N_VDD_c_337_p N_A_1469_521#_c_2171_n 0.00757793f $X=7.815 $Y=4.287
+ $X2=7.47 $Y2=3.295
cc_418 N_VDD_c_269_p N_A_1469_521#_c_2171_n 0.00476261f $X=9.855 $Y=4.25
+ $X2=7.47 $Y2=3.295
cc_419 N_VDD_M1033_d N_A_1469_521#_c_2174_n 0.0038492f $X=7.76 $Y=2.605
+ $X2=8.245 $Y2=3.185
cc_420 N_VDD_c_290_p N_A_1469_521#_c_2174_n 0.00891306f $X=7.9 $Y=3.7 $X2=8.245
+ $Y2=3.185
cc_421 N_VDD_M1001_b N_A_1469_521#_c_2176_n 0.00155118f $X=-0.05 $Y=2.425
+ $X2=8.33 $Y2=3.295
cc_422 N_VDD_c_279_p N_A_1469_521#_c_2176_n 0.00739652f $X=9.625 $Y=4.287
+ $X2=8.33 $Y2=3.295
cc_423 N_VDD_c_269_p N_A_1469_521#_c_2176_n 0.00475776f $X=9.855 $Y=4.25
+ $X2=8.33 $Y2=3.295
cc_424 N_VDD_M1001_b N_Q_c_2195_n 0.00156053f $X=-0.05 $Y=2.425 $X2=10.14
+ $Y2=2.85
cc_425 N_VDD_c_399_p N_Q_c_2195_n 0.0075728f $X=9.855 $Y=4.22 $X2=10.14 $Y2=2.85
cc_426 N_VDD_c_269_p N_Q_c_2195_n 0.00476261f $X=9.855 $Y=4.25 $X2=10.14
+ $Y2=2.85
cc_427 N_VDD_M1001_b N_Q_c_2193_n 0.00544948f $X=-0.05 $Y=2.425 $X2=10.255
+ $Y2=2.525
cc_428 N_VDD_M1001_b N_Q_c_2199_n 0.0144447f $X=-0.05 $Y=2.425 $X2=10.255
+ $Y2=2.61
cc_429 N_VDD_M1001_b Q 0.00983408f $X=-0.05 $Y=2.425 $X2=10.14 $Y2=2.85
cc_430 N_VDD_c_376_p Q 0.00673193f $X=9.71 $Y=2.955 $X2=10.14 $Y2=2.85
cc_431 RN N_A_110_115#_M1001_d 0.00410657f $X=0.325 $Y=2.85 $X2=0.55 $Y2=2.605
cc_432 N_RN_M1016_g N_A_110_115#_c_473_n 0.00226126f $X=0.475 $Y=0.85 $X2=1.29
+ $Y2=2.32
cc_433 N_RN_c_436_n N_A_110_115#_c_473_n 0.00491604f $X=0.475 $Y=1.99 $X2=1.29
+ $Y2=2.32
cc_434 N_RN_M1001_g N_A_110_115#_c_473_n 0.00480617f $X=0.475 $Y=3.235 $X2=1.29
+ $Y2=2.32
cc_435 N_RN_M1016_g N_A_110_115#_c_485_n 0.00475169f $X=0.475 $Y=0.85 $X2=1.29
+ $Y2=1.27
cc_436 N_RN_M1016_g N_A_110_115#_c_490_n 0.0047157f $X=0.475 $Y=0.85 $X2=0.69
+ $Y2=0.755
cc_437 N_RN_M1001_g N_A_110_115#_c_494_n 0.00835855f $X=0.475 $Y=3.235 $X2=0.69
+ $Y2=2.955
cc_438 N_RN_c_438_n N_A_110_115#_c_494_n 0.0282684f $X=0.32 $Y=2.85 $X2=0.69
+ $Y2=2.955
cc_439 RN N_A_110_115#_c_494_n 0.00974028f $X=0.325 $Y=2.85 $X2=0.69 $Y2=2.955
cc_440 N_RN_M1016_g N_A_110_115#_c_495_n 0.00620105f $X=0.475 $Y=0.85 $X2=0.87
+ $Y2=1.37
cc_441 N_RN_c_436_n N_A_110_115#_c_495_n 0.00325637f $X=0.475 $Y=1.99 $X2=0.87
+ $Y2=1.37
cc_442 N_RN_M1001_g N_A_110_115#_c_495_n 0.00186244f $X=0.475 $Y=3.235 $X2=0.87
+ $Y2=1.37
cc_443 N_RN_c_438_n N_A_110_115#_c_495_n 0.0072511f $X=0.32 $Y=2.85 $X2=0.87
+ $Y2=1.37
cc_444 N_RN_c_439_n N_A_110_115#_c_495_n 0.0248372f $X=0.32 $Y=1.825 $X2=0.87
+ $Y2=1.37
cc_445 N_RN_M1016_g N_A_110_115#_c_496_n 0.00584255f $X=0.475 $Y=0.85 $X2=0.955
+ $Y2=1.27
cc_446 N_RN_c_436_n N_A_110_115#_c_496_n 0.00168842f $X=0.475 $Y=1.99 $X2=0.955
+ $Y2=1.27
cc_447 N_RN_c_439_n N_A_110_115#_c_496_n 4.87394e-19 $X=0.32 $Y=1.825 $X2=0.955
+ $Y2=1.27
cc_448 N_RN_c_436_n N_A_110_115#_c_499_n 0.00191737f $X=0.475 $Y=1.99 $X2=0.87
+ $Y2=2.26
cc_449 N_RN_M1001_g N_A_110_115#_c_499_n 0.00207383f $X=0.475 $Y=3.235 $X2=0.87
+ $Y2=2.26
cc_450 N_RN_c_438_n N_A_110_115#_c_499_n 0.0113366f $X=0.32 $Y=2.85 $X2=0.87
+ $Y2=2.26
cc_451 N_RN_c_439_n N_A_110_115#_c_499_n 7.08415e-19 $X=0.32 $Y=1.825 $X2=0.87
+ $Y2=2.26
cc_452 N_RN_M1016_g N_A_110_115#_c_527_n 0.00223114f $X=0.475 $Y=0.85 $X2=0.87
+ $Y2=1.37
cc_453 N_RN_M1001_g N_A_217_521#_c_1309_n 0.00351056f $X=0.475 $Y=3.235 $X2=1.21
+ $Y2=3.295
cc_454 RN N_A_217_521#_c_1309_n 9.10636e-19 $X=0.325 $Y=2.85 $X2=1.21 $Y2=3.295
cc_455 N_A_110_115#_c_485_n N_SN_c_703_n 0.00643294f $X=1.29 $Y=1.27 $X2=1.89
+ $Y2=1.405
cc_456 N_A_110_115#_c_503_n N_SN_c_703_n 2.91248e-19 $X=8.775 $Y=1 $X2=1.89
+ $Y2=1.405
cc_457 N_A_110_115#_c_473_n N_SN_c_704_n 0.00643294f $X=1.29 $Y=2.32 $X2=1.89
+ $Y2=1.785
cc_458 N_A_110_115#_c_473_n N_SN_M1024_g 0.0048371f $X=1.29 $Y=2.32 $X2=1.855
+ $Y2=3.235
cc_459 N_A_110_115#_c_484_n N_SN_M1024_g 0.0396474f $X=1.425 $Y=2.395 $X2=1.855
+ $Y2=3.235
cc_460 N_A_110_115#_c_474_n N_SN_M1015_g 0.0208493f $X=1.435 $Y=1.105 $X2=1.925
+ $Y2=0.85
cc_461 N_A_110_115#_c_485_n N_SN_M1015_g 6.85742e-19 $X=1.29 $Y=1.27 $X2=1.925
+ $Y2=0.85
cc_462 N_A_110_115#_c_503_n N_SN_M1015_g 0.00618821f $X=8.775 $Y=1 $X2=1.925
+ $Y2=0.85
cc_463 N_A_110_115#_c_478_n N_SN_M1004_g 0.0205825f $X=8.535 $Y=1.105 $X2=8.045
+ $Y2=0.85
cc_464 N_A_110_115#_c_487_n N_SN_M1004_g 0.00449705f $X=8.8 $Y=1.27 $X2=8.045
+ $Y2=0.85
cc_465 N_A_110_115#_c_503_n N_SN_M1004_g 0.00660386f $X=8.775 $Y=1 $X2=8.045
+ $Y2=0.85
cc_466 N_A_110_115#_c_489_n N_SN_M1019_g 0.0463249f $X=8.545 $Y=2.27 $X2=8.115
+ $Y2=3.235
cc_467 N_A_110_115#_c_473_n N_SN_c_713_n 0.0200438f $X=1.29 $Y=2.32 $X2=1.855
+ $Y2=1.95
cc_468 N_A_110_115#_c_483_n N_SN_c_714_n 0.00935305f $X=8.8 $Y=2.125 $X2=8.02
+ $Y2=1.775
cc_469 N_A_110_115#_c_503_n N_SN_c_714_n 0.00219437f $X=8.775 $Y=1 $X2=8.02
+ $Y2=1.775
cc_470 N_A_110_115#_c_473_n N_SN_c_715_n 0.00173691f $X=1.29 $Y=2.32 $X2=1.71
+ $Y2=2.62
cc_471 N_A_110_115#_c_484_n N_SN_c_715_n 0.00247884f $X=1.425 $Y=2.395 $X2=1.71
+ $Y2=2.62
cc_472 N_A_110_115#_c_473_n N_SN_c_717_n 0.00103414f $X=1.29 $Y=2.32 $X2=1.71
+ $Y2=1.95
cc_473 N_A_110_115#_M1000_g N_SN_c_732_n 0.0018081f $X=1.425 $Y=3.235 $X2=1.71
+ $Y2=2.777
cc_474 N_A_110_115#_c_483_n N_SN_c_718_n 2.69784e-19 $X=8.8 $Y=2.125 $X2=8.02
+ $Y2=1.775
cc_475 N_A_110_115#_c_503_n N_SN_c_718_n 0.00344841f $X=8.775 $Y=1 $X2=8.02
+ $Y2=1.775
cc_476 N_A_110_115#_M1000_g N_SN_c_742_n 7.05054e-19 $X=1.425 $Y=3.235 $X2=2.195
+ $Y2=2.85
cc_477 N_A_110_115#_M1025_g SN 0.00109708f $X=8.545 $Y=3.235 $X2=7.94 $Y2=2.845
cc_478 N_A_110_115#_c_503_n N_A_432_424#_M1035_d 0.00324609f $X=8.775 $Y=1
+ $X2=3.67 $Y2=0.575
cc_479 N_A_110_115#_c_503_n N_A_432_424#_M1003_g 0.00683876f $X=8.775 $Y=1
+ $X2=2.285 $Y2=0.85
cc_480 N_A_110_115#_c_503_n N_A_432_424#_c_902_n 0.0295499f $X=8.775 $Y=1
+ $X2=3.71 $Y2=1.285
cc_481 N_A_110_115#_c_503_n N_A_432_424#_c_905_n 0.00540043f $X=8.775 $Y=1
+ $X2=2.38 $Y2=1.285
cc_482 N_A_110_115#_c_503_n N_A_432_424#_c_908_n 0.0151351f $X=8.775 $Y=1
+ $X2=3.795 $Y2=1.2
cc_483 N_A_110_115#_c_503_n N_A_432_424#_c_909_n 0.0133933f $X=8.775 $Y=1
+ $X2=3.795 $Y2=0.755
cc_484 N_A_110_115#_c_503_n N_D_M1005_g 0.00683925f $X=8.775 $Y=1 $X2=3.235
+ $Y2=0.85
cc_485 N_A_110_115#_c_503_n N_CK_c_1046_n 7.89968e-19 $X=8.775 $Y=1 $X2=4.135
+ $Y2=1.4
cc_486 N_A_110_115#_c_503_n N_CK_c_1047_n 0.0064365f $X=8.775 $Y=1 $X2=4.135
+ $Y2=1.235
cc_487 N_A_110_115#_c_503_n N_CK_c_1050_n 7.89968e-19 $X=8.775 $Y=1 $X2=5.405
+ $Y2=1.4
cc_488 N_A_110_115#_c_503_n N_CK_c_1051_n 0.00634331f $X=8.775 $Y=1 $X2=5.405
+ $Y2=1.235
cc_489 N_A_110_115#_c_503_n N_CK_c_1055_n 0.00713721f $X=8.775 $Y=1 $X2=6.762
+ $Y2=1.205
cc_490 N_A_110_115#_c_503_n N_CK_c_1060_n 0.00107886f $X=8.775 $Y=1 $X2=6.762
+ $Y2=1.355
cc_491 N_A_110_115#_c_503_n N_CK_c_1062_n 0.00475893f $X=8.775 $Y=1 $X2=4.135
+ $Y2=1.4
cc_492 N_A_110_115#_c_503_n N_CK_c_1063_n 0.00475709f $X=8.775 $Y=1 $X2=5.405
+ $Y2=1.4
cc_493 N_A_110_115#_c_503_n N_A_217_521#_M1034_d 0.00288434f $X=8.775 $Y=1
+ $X2=1.51 $Y2=0.575
cc_494 N_A_110_115#_c_503_n N_A_217_521#_M1020_g 0.00607163f $X=8.775 $Y=1
+ $X2=4.555 $Y2=0.85
cc_495 N_A_110_115#_c_503_n N_A_217_521#_c_1300_n 2.38222e-19 $X=8.775 $Y=1
+ $X2=4.91 $Y2=1.4
cc_496 N_A_110_115#_c_503_n N_A_217_521#_M1023_g 0.00633529f $X=8.775 $Y=1
+ $X2=4.985 $Y2=0.85
cc_497 N_A_110_115#_c_473_n N_A_217_521#_c_1309_n 0.0184538f $X=1.29 $Y=2.32
+ $X2=1.21 $Y2=3.295
cc_498 N_A_110_115#_M1000_g N_A_217_521#_c_1309_n 0.0133902f $X=1.425 $Y=3.235
+ $X2=1.21 $Y2=3.295
cc_499 N_A_110_115#_c_484_n N_A_217_521#_c_1309_n 0.00692138f $X=1.425 $Y=2.395
+ $X2=1.21 $Y2=3.295
cc_500 N_A_110_115#_c_494_n N_A_217_521#_c_1309_n 0.0646924f $X=0.69 $Y=2.955
+ $X2=1.21 $Y2=3.295
cc_501 N_A_110_115#_c_495_n N_A_217_521#_c_1309_n 0.0361025f $X=0.87 $Y=1.37
+ $X2=1.21 $Y2=3.295
cc_502 N_A_110_115#_c_499_n N_A_217_521#_c_1309_n 0.0134429f $X=0.87 $Y=2.26
+ $X2=1.21 $Y2=3.295
cc_503 N_A_110_115#_c_473_n N_A_217_521#_c_1310_n 0.00698097f $X=1.29 $Y=2.32
+ $X2=1.565 $Y2=1.61
cc_504 N_A_110_115#_c_484_n N_A_217_521#_c_1310_n 0.00349831f $X=1.425 $Y=2.395
+ $X2=1.565 $Y2=1.61
cc_505 N_A_110_115#_c_485_n N_A_217_521#_c_1310_n 0.00449938f $X=1.29 $Y=1.27
+ $X2=1.565 $Y2=1.61
cc_506 N_A_110_115#_c_497_n N_A_217_521#_c_1310_n 0.00666591f $X=1.23 $Y=1.27
+ $X2=1.565 $Y2=1.61
cc_507 N_A_110_115#_c_503_n N_A_217_521#_c_1310_n 0.00580834f $X=8.775 $Y=1
+ $X2=1.565 $Y2=1.61
cc_508 N_A_110_115#_c_473_n N_A_217_521#_c_1311_n 0.00443913f $X=1.29 $Y=2.32
+ $X2=1.295 $Y2=1.61
cc_509 N_A_110_115#_c_485_n N_A_217_521#_c_1311_n 0.00231083f $X=1.29 $Y=1.27
+ $X2=1.295 $Y2=1.61
cc_510 N_A_110_115#_c_495_n N_A_217_521#_c_1311_n 0.0138602f $X=0.87 $Y=1.37
+ $X2=1.295 $Y2=1.61
cc_511 N_A_110_115#_c_497_n N_A_217_521#_c_1311_n 0.0126994f $X=1.23 $Y=1.27
+ $X2=1.295 $Y2=1.61
cc_512 N_A_110_115#_c_474_n N_A_217_521#_c_1312_n 0.00936975f $X=1.435 $Y=1.105
+ $X2=1.71 $Y2=0.755
cc_513 N_A_110_115#_c_485_n N_A_217_521#_c_1312_n 0.00114928f $X=1.29 $Y=1.27
+ $X2=1.71 $Y2=0.755
cc_514 N_A_110_115#_c_495_n N_A_217_521#_c_1312_n 0.00143024f $X=0.87 $Y=1.37
+ $X2=1.71 $Y2=0.755
cc_515 N_A_110_115#_c_497_n N_A_217_521#_c_1312_n 0.00961285f $X=1.23 $Y=1.27
+ $X2=1.71 $Y2=0.755
cc_516 N_A_110_115#_c_503_n N_A_217_521#_c_1312_n 0.0198038f $X=8.775 $Y=1
+ $X2=1.71 $Y2=0.755
cc_517 N_A_110_115#_c_527_n N_A_217_521#_c_1312_n 5.78004e-19 $X=0.87 $Y=1.37
+ $X2=1.71 $Y2=0.755
cc_518 N_A_110_115#_c_473_n N_A_217_521#_c_1316_n 9.49852e-19 $X=1.29 $Y=2.32
+ $X2=1.68 $Y2=1.61
cc_519 N_A_110_115#_c_495_n N_A_217_521#_c_1316_n 0.00179145f $X=0.87 $Y=1.37
+ $X2=1.68 $Y2=1.61
cc_520 N_A_110_115#_c_503_n N_A_217_521#_c_1316_n 2.82351e-19 $X=8.775 $Y=1
+ $X2=1.68 $Y2=1.61
cc_521 N_A_110_115#_c_503_n N_A_217_521#_c_1317_n 0.00469682f $X=8.775 $Y=1
+ $X2=4.725 $Y2=1.4
cc_522 N_A_110_115#_c_503_n N_A_217_521#_c_1319_n 0.212989f $X=8.775 $Y=1
+ $X2=4.49 $Y2=1.37
cc_523 N_A_110_115#_c_485_n N_A_217_521#_c_1320_n 0.00123792f $X=1.29 $Y=1.27
+ $X2=1.855 $Y2=1.37
cc_524 N_A_110_115#_c_495_n N_A_217_521#_c_1320_n 7.31862e-19 $X=0.87 $Y=1.37
+ $X2=1.855 $Y2=1.37
cc_525 N_A_110_115#_c_497_n N_A_217_521#_c_1320_n 0.00150041f $X=1.23 $Y=1.27
+ $X2=1.855 $Y2=1.37
cc_526 N_A_110_115#_c_503_n N_A_217_521#_c_1320_n 0.0252928f $X=8.775 $Y=1
+ $X2=1.855 $Y2=1.37
cc_527 N_A_110_115#_c_527_n N_A_217_521#_c_1320_n 0.0119249f $X=0.87 $Y=1.37
+ $X2=1.855 $Y2=1.37
cc_528 N_A_110_115#_c_503_n N_A_217_521#_c_1372_n 0.0259855f $X=8.775 $Y=1
+ $X2=4.635 $Y2=1.37
cc_529 N_A_110_115#_c_503_n N_A_704_89#_M1011_d 0.00194184f $X=8.775 $Y=1
+ $X2=6.81 $Y2=0.575
cc_530 N_A_110_115#_c_503_n N_A_704_89#_c_1460_n 0.00599689f $X=8.775 $Y=1
+ $X2=3.595 $Y2=1.205
cc_531 N_A_110_115#_c_503_n N_A_704_89#_M1017_g 0.00631343f $X=8.775 $Y=1
+ $X2=5.945 $Y2=0.85
cc_532 N_A_110_115#_c_503_n N_A_704_89#_c_1478_n 0.0194702f $X=8.775 $Y=1
+ $X2=6.95 $Y2=0.755
cc_533 N_A_110_115#_c_503_n N_A_1246_89#_M1004_d 0.00313302f $X=8.775 $Y=1
+ $X2=8.12 $Y2=0.575
cc_534 N_A_110_115#_c_503_n N_A_1246_89#_M1006_g 0.0058983f $X=8.775 $Y=1
+ $X2=6.305 $Y2=0.85
cc_535 N_A_110_115#_c_483_n N_A_1246_89#_c_1679_n 0.0112463f $X=8.8 $Y=2.125
+ $X2=9.38 $Y2=1.71
cc_536 N_A_110_115#_c_483_n N_A_1246_89#_c_1680_n 0.00290928f $X=8.8 $Y=2.125
+ $X2=9.382 $Y2=1.545
cc_537 N_A_110_115#_c_528_n N_A_1246_89#_c_1680_n 4.37027e-19 $X=8.86 $Y=1.37
+ $X2=9.382 $Y2=1.545
cc_538 N_A_110_115#_c_487_n N_A_1246_89#_c_1681_n 0.00268913f $X=8.8 $Y=1.27
+ $X2=9.47 $Y2=1.23
cc_539 N_A_110_115#_c_487_n N_A_1246_89#_c_1686_n 0.00630476f $X=8.8 $Y=1.27
+ $X2=9.47 $Y2=1.38
cc_540 N_A_110_115#_c_500_n N_A_1246_89#_c_1686_n 3.89361e-19 $X=8.86 $Y=1.27
+ $X2=9.47 $Y2=1.38
cc_541 N_A_110_115#_c_483_n N_A_1246_89#_c_1687_n 0.00978182f $X=8.8 $Y=2.125
+ $X2=9.47 $Y2=2.375
cc_542 N_A_110_115#_c_489_n N_A_1246_89#_c_1687_n 0.00180274f $X=8.545 $Y=2.27
+ $X2=9.47 $Y2=2.375
cc_543 N_A_110_115#_c_478_n N_A_1246_89#_c_1690_n 0.00942337f $X=8.535 $Y=1.105
+ $X2=8.26 $Y2=0.755
cc_544 N_A_110_115#_c_487_n N_A_1246_89#_c_1690_n 3.37028e-19 $X=8.8 $Y=1.27
+ $X2=8.26 $Y2=0.755
cc_545 N_A_110_115#_c_500_n N_A_1246_89#_c_1690_n 0.0062056f $X=8.86 $Y=1.27
+ $X2=8.26 $Y2=0.755
cc_546 N_A_110_115#_c_503_n N_A_1246_89#_c_1690_n 0.0216418f $X=8.775 $Y=1
+ $X2=8.26 $Y2=0.755
cc_547 N_A_110_115#_c_528_n N_A_1246_89#_c_1690_n 5.9368e-19 $X=8.86 $Y=1.37
+ $X2=8.26 $Y2=0.755
cc_548 N_A_110_115#_c_529_n N_A_1246_89#_c_1690_n 0.00371946f $X=8.862 $Y=1.255
+ $X2=8.26 $Y2=0.755
cc_549 N_A_110_115#_M1025_g N_A_1246_89#_c_1693_n 0.0154027f $X=8.545 $Y=3.235
+ $X2=8.76 $Y2=3.295
cc_550 N_A_110_115#_c_483_n N_A_1246_89#_c_1693_n 0.0115916f $X=8.8 $Y=2.125
+ $X2=8.76 $Y2=3.295
cc_551 N_A_110_115#_c_489_n N_A_1246_89#_c_1693_n 0.0174845f $X=8.545 $Y=2.27
+ $X2=8.76 $Y2=3.295
cc_552 N_A_110_115#_c_483_n N_A_1246_89#_c_1694_n 0.00574194f $X=8.8 $Y=2.125
+ $X2=8.845 $Y2=1.71
cc_553 N_A_110_115#_c_487_n N_A_1246_89#_c_1694_n 0.0128134f $X=8.8 $Y=1.27
+ $X2=8.845 $Y2=1.71
cc_554 N_A_110_115#_c_489_n N_A_1246_89#_c_1694_n 0.00546847f $X=8.545 $Y=2.27
+ $X2=8.845 $Y2=1.71
cc_555 N_A_110_115#_c_500_n N_A_1246_89#_c_1694_n 0.0130331f $X=8.86 $Y=1.27
+ $X2=8.845 $Y2=1.71
cc_556 N_A_110_115#_c_503_n N_A_1246_89#_c_1694_n 0.0067495f $X=8.775 $Y=1
+ $X2=8.845 $Y2=1.71
cc_557 N_A_110_115#_c_528_n N_A_1246_89#_c_1694_n 0.00526093f $X=8.86 $Y=1.37
+ $X2=8.845 $Y2=1.71
cc_558 N_A_110_115#_c_483_n N_A_1246_89#_c_1695_n 0.00377526f $X=8.8 $Y=2.125
+ $X2=9.38 $Y2=1.71
cc_559 N_A_110_115#_c_487_n N_A_1246_89#_c_1695_n 0.00127281f $X=8.8 $Y=1.27
+ $X2=9.38 $Y2=1.71
cc_560 N_A_110_115#_c_500_n N_A_1246_89#_c_1695_n 0.0103258f $X=8.86 $Y=1.27
+ $X2=9.38 $Y2=1.71
cc_561 N_A_110_115#_c_528_n N_A_1246_89#_c_1695_n 6.55882e-19 $X=8.86 $Y=1.37
+ $X2=9.38 $Y2=1.71
cc_562 N_A_110_115#_c_483_n N_A_1246_89#_c_1698_n 0.00196012f $X=8.8 $Y=2.125
+ $X2=9.235 $Y2=1.71
cc_563 N_A_110_115#_c_487_n N_A_1246_89#_c_1698_n 2.4916e-19 $X=8.8 $Y=1.27
+ $X2=9.235 $Y2=1.71
cc_564 N_A_110_115#_c_500_n N_A_1246_89#_c_1698_n 0.00128974f $X=8.86 $Y=1.27
+ $X2=9.235 $Y2=1.71
cc_565 N_A_110_115#_c_503_n N_A_1246_89#_c_1698_n 0.0444699f $X=8.775 $Y=1
+ $X2=9.235 $Y2=1.71
cc_566 N_A_110_115#_c_528_n N_A_1246_89#_c_1698_n 0.0300972f $X=8.86 $Y=1.37
+ $X2=9.235 $Y2=1.71
cc_567 N_A_110_115#_c_483_n N_A_1246_89#_c_1701_n 8.29185e-19 $X=8.8 $Y=2.125
+ $X2=9.38 $Y2=1.71
cc_568 N_A_110_115#_c_503_n N_A_1084_115#_M1021_d 0.00325279f $X=8.775 $Y=1
+ $X2=5.42 $Y2=0.575
cc_569 N_A_110_115#_c_503_n N_A_1084_115#_c_1884_n 0.00717782f $X=8.775 $Y=1
+ $X2=7.685 $Y2=1.21
cc_570 N_A_110_115#_c_503_n N_A_1084_115#_c_1888_n 0.00328689f $X=8.775 $Y=1
+ $X2=7.685 $Y2=1.29
cc_571 N_A_110_115#_c_503_n N_A_1084_115#_c_1891_n 0.00535229f $X=8.775 $Y=1
+ $X2=5.065 $Y2=1.37
cc_572 N_A_110_115#_c_503_n N_A_1084_115#_c_1892_n 0.00625719f $X=8.775 $Y=1
+ $X2=5.745 $Y2=1.34
cc_573 N_A_110_115#_c_503_n N_A_1084_115#_c_1893_n 0.00241187f $X=8.775 $Y=1
+ $X2=7.595 $Y2=1.37
cc_574 N_A_110_115#_c_503_n N_A_1084_115#_c_1895_n 0.0230942f $X=8.775 $Y=1
+ $X2=5.645 $Y2=0.755
cc_575 N_A_110_115#_c_503_n N_A_1084_115#_c_1898_n 0.0320068f $X=8.775 $Y=1
+ $X2=5.6 $Y2=1.37
cc_576 N_A_110_115#_c_503_n N_A_1084_115#_c_1899_n 0.0259535f $X=8.775 $Y=1
+ $X2=5.21 $Y2=1.37
cc_577 N_A_110_115#_c_503_n N_A_1084_115#_c_1900_n 0.130211f $X=8.775 $Y=1
+ $X2=7.45 $Y2=1.37
cc_578 N_A_110_115#_c_503_n N_A_1084_115#_c_1903_n 0.0270067f $X=8.775 $Y=1
+ $X2=5.89 $Y2=1.37
cc_579 N_A_110_115#_c_503_n N_A_1084_115#_c_1904_n 0.0265552f $X=8.775 $Y=1
+ $X2=7.595 $Y2=1.37
cc_580 N_A_110_115#_c_478_n N_QN_c_2065_n 0.00411421f $X=8.535 $Y=1.105 $X2=9.28
+ $Y2=0.755
cc_581 N_A_110_115#_c_487_n N_QN_c_2065_n 0.00214646f $X=8.8 $Y=1.27 $X2=9.28
+ $Y2=0.755
cc_582 N_A_110_115#_c_500_n N_QN_c_2065_n 0.00731463f $X=8.86 $Y=1.27 $X2=9.28
+ $Y2=0.755
cc_583 N_A_110_115#_c_503_n N_QN_c_2065_n 0.0123459f $X=8.775 $Y=1 $X2=9.28
+ $Y2=0.755
cc_584 N_A_110_115#_c_528_n N_QN_c_2065_n 2.14408e-19 $X=8.86 $Y=1.37 $X2=9.28
+ $Y2=0.755
cc_585 N_A_110_115#_c_529_n N_QN_c_2065_n 4.33654e-19 $X=8.862 $Y=1.255 $X2=9.28
+ $Y2=0.755
cc_586 N_A_110_115#_c_487_n N_QN_c_2072_n 8.77889e-19 $X=8.8 $Y=1.27 $X2=9.365
+ $Y2=1.37
cc_587 N_A_110_115#_c_500_n N_QN_c_2072_n 0.0102707f $X=8.86 $Y=1.27 $X2=9.365
+ $Y2=1.37
cc_588 N_A_110_115#_c_528_n N_QN_c_2072_n 0.00363844f $X=8.86 $Y=1.37 $X2=9.365
+ $Y2=1.37
cc_589 N_A_110_115#_c_489_n N_QN_c_2074_n 0.00115295f $X=8.545 $Y=2.27 $X2=9.365
+ $Y2=2.285
cc_590 N_A_110_115#_c_503_n A_400_115# 0.00473401f $X=8.775 $Y=1 $X2=2 $Y2=0.575
cc_591 N_A_110_115#_c_503_n A_662_115# 0.00381028f $X=8.775 $Y=1 $X2=3.31
+ $Y2=0.575
cc_592 N_A_110_115#_c_503_n A_854_115# 0.00473401f $X=8.775 $Y=1 $X2=4.27
+ $Y2=0.575
cc_593 N_A_110_115#_c_503_n A_1012_115# 0.00430069f $X=8.775 $Y=1 $X2=5.06
+ $Y2=0.575
cc_594 N_A_110_115#_c_503_n A_1204_115# 0.00466077f $X=8.775 $Y=1 $X2=6.02
+ $Y2=0.575
cc_595 N_A_110_115#_c_503_n A_1552_115# 0.00533054f $X=8.775 $Y=1 $X2=7.76
+ $Y2=0.575
cc_596 N_SN_c_733_n N_A_432_424#_M1018_d 0.004688f $X=7.79 $Y=2.85 $X2=3.67
+ $Y2=2.605
cc_597 N_SN_M1015_g N_A_432_424#_M1003_g 0.0939126f $X=1.925 $Y=0.85 $X2=2.285
+ $Y2=0.85
cc_598 N_SN_c_713_n N_A_432_424#_M1003_g 0.00639789f $X=1.855 $Y=1.95 $X2=2.285
+ $Y2=0.85
cc_599 N_SN_c_715_n N_A_432_424#_M1003_g 2.30594e-19 $X=1.71 $Y=2.62 $X2=2.285
+ $Y2=0.85
cc_600 N_SN_c_717_n N_A_432_424#_M1003_g 4.68111e-19 $X=1.71 $Y=1.95 $X2=2.285
+ $Y2=0.85
cc_601 N_SN_M1024_g N_A_432_424#_M1027_g 0.0520248f $X=1.855 $Y=3.235 $X2=2.285
+ $Y2=3.235
cc_602 N_SN_c_715_n N_A_432_424#_M1027_g 8.16515e-19 $X=1.71 $Y=2.62 $X2=2.285
+ $Y2=3.235
cc_603 N_SN_c_732_n N_A_432_424#_M1027_g 0.00503122f $X=1.71 $Y=2.777 $X2=2.285
+ $Y2=3.235
cc_604 N_SN_c_733_n N_A_432_424#_M1027_g 0.0077142f $X=7.79 $Y=2.85 $X2=2.285
+ $Y2=3.235
cc_605 N_SN_c_742_n N_A_432_424#_M1027_g 0.00102878f $X=2.195 $Y=2.85 $X2=2.285
+ $Y2=3.235
cc_606 N_SN_M1024_g N_A_432_424#_c_900_n 0.0173689f $X=1.855 $Y=3.235 $X2=2.295
+ $Y2=2.285
cc_607 N_SN_c_715_n N_A_432_424#_c_900_n 9.68052e-19 $X=1.71 $Y=2.62 $X2=2.295
+ $Y2=2.285
cc_608 N_SN_c_733_n N_A_432_424#_c_900_n 0.0014689f $X=7.79 $Y=2.85 $X2=2.295
+ $Y2=2.285
cc_609 N_SN_c_742_n N_A_432_424#_c_900_n 8.46214e-19 $X=2.195 $Y=2.85 $X2=2.295
+ $Y2=2.285
cc_610 N_SN_c_703_n N_A_432_424#_c_901_n 0.00287608f $X=1.89 $Y=1.405 $X2=2.295
+ $Y2=2.2
cc_611 N_SN_M1024_g N_A_432_424#_c_901_n 7.93818e-19 $X=1.855 $Y=3.235 $X2=2.295
+ $Y2=2.2
cc_612 N_SN_c_713_n N_A_432_424#_c_901_n 8.91506e-19 $X=1.855 $Y=1.95 $X2=2.295
+ $Y2=2.2
cc_613 N_SN_c_715_n N_A_432_424#_c_901_n 0.0142773f $X=1.71 $Y=2.62 $X2=2.295
+ $Y2=2.2
cc_614 N_SN_c_717_n N_A_432_424#_c_901_n 0.00704932f $X=1.71 $Y=1.95 $X2=2.295
+ $Y2=2.2
cc_615 N_SN_c_733_n N_A_432_424#_c_901_n 0.00424733f $X=7.79 $Y=2.85 $X2=2.295
+ $Y2=2.2
cc_616 N_SN_M1015_g N_A_432_424#_c_905_n 6.84827e-19 $X=1.925 $Y=0.85 $X2=2.38
+ $Y2=1.285
cc_617 N_SN_c_733_n N_A_432_424#_c_906_n 0.0111257f $X=7.79 $Y=2.85 $X2=2.685
+ $Y2=2.285
cc_618 N_SN_c_733_n N_A_432_424#_c_920_n 0.0722563f $X=7.79 $Y=2.85 $X2=3.725
+ $Y2=2.705
cc_619 N_SN_c_732_n N_A_432_424#_c_923_n 0.0056303f $X=1.71 $Y=2.777 $X2=2.855
+ $Y2=2.705
cc_620 N_SN_c_733_n N_A_432_424#_c_923_n 0.0150027f $X=7.79 $Y=2.85 $X2=2.855
+ $Y2=2.705
cc_621 N_SN_c_742_n N_A_432_424#_c_923_n 7.56538e-19 $X=2.195 $Y=2.85 $X2=2.855
+ $Y2=2.705
cc_622 N_SN_c_733_n N_A_432_424#_c_924_n 0.0225196f $X=7.79 $Y=2.85 $X2=3.895
+ $Y2=2.955
cc_623 N_SN_c_733_n N_D_M1028_g 0.00954918f $X=7.79 $Y=2.85 $X2=3.235 $Y2=3.235
cc_624 N_SN_c_733_n N_CK_M1018_g 0.00848309f $X=7.79 $Y=2.85 $X2=3.595 $Y2=3.235
cc_625 N_SN_c_733_n N_CK_M1002_g 0.011385f $X=7.79 $Y=2.85 $X2=5.945 $Y2=3.235
cc_626 N_SN_c_733_n N_CK_M1031_g 0.0092737f $X=7.79 $Y=2.85 $X2=6.735 $Y2=3.235
cc_627 N_SN_c_733_n N_CK_c_1061_n 0.00366725f $X=7.79 $Y=2.85 $X2=4.05 $Y2=2.11
cc_628 N_SN_c_733_n N_CK_c_1064_n 7.28286e-19 $X=7.79 $Y=2.85 $X2=5.77 $Y2=2.11
cc_629 N_SN_c_733_n N_CK_c_1065_n 5.66698e-19 $X=7.79 $Y=2.85 $X2=5.49 $Y2=2.11
cc_630 N_SN_c_733_n N_CK_c_1066_n 0.00112396f $X=7.79 $Y=2.85 $X2=6.88 $Y2=2.11
cc_631 N_SN_c_733_n N_CK_c_1067_n 6.09336e-19 $X=7.79 $Y=2.85 $X2=3.655 $Y2=2.11
cc_632 N_SN_c_733_n N_CK_c_1068_n 0.00366727f $X=7.79 $Y=2.85 $X2=5.885 $Y2=2.11
cc_633 N_SN_c_733_n N_CK_c_1070_n 0.0119585f $X=7.79 $Y=2.85 $X2=3.8 $Y2=2.11
cc_634 N_SN_c_733_n N_CK_c_1072_n 0.0128795f $X=7.79 $Y=2.85 $X2=6.03 $Y2=2.11
cc_635 N_SN_c_733_n N_A_217_521#_M1009_g 0.0155696f $X=7.79 $Y=2.85 $X2=4.555
+ $Y2=3.235
cc_636 N_SN_c_733_n N_A_217_521#_c_1303_n 2.37802e-19 $X=7.79 $Y=2.85 $X2=4.91
+ $Y2=2.285
cc_637 N_SN_c_733_n N_A_217_521#_M1012_g 0.0112548f $X=7.79 $Y=2.85 $X2=4.985
+ $Y2=3.235
cc_638 N_SN_c_704_n N_A_217_521#_c_1309_n 4.72187e-19 $X=1.89 $Y=1.785 $X2=1.21
+ $Y2=3.295
cc_639 N_SN_M1024_g N_A_217_521#_c_1309_n 3.15481e-19 $X=1.855 $Y=3.235 $X2=1.21
+ $Y2=3.295
cc_640 N_SN_c_713_n N_A_217_521#_c_1309_n 9.48304e-19 $X=1.855 $Y=1.95 $X2=1.21
+ $Y2=3.295
cc_641 N_SN_c_715_n N_A_217_521#_c_1309_n 0.0253396f $X=1.71 $Y=2.62 $X2=1.21
+ $Y2=3.295
cc_642 N_SN_c_717_n N_A_217_521#_c_1309_n 0.00963813f $X=1.71 $Y=1.95 $X2=1.21
+ $Y2=3.295
cc_643 N_SN_c_742_n N_A_217_521#_c_1309_n 0.00373659f $X=2.195 $Y=2.85 $X2=1.21
+ $Y2=3.295
cc_644 N_SN_c_717_n N_A_217_521#_c_1310_n 0.00143797f $X=1.71 $Y=1.95 $X2=1.565
+ $Y2=1.61
cc_645 N_SN_c_703_n N_A_217_521#_c_1312_n 0.00283874f $X=1.89 $Y=1.405 $X2=1.71
+ $Y2=0.755
cc_646 N_SN_c_704_n N_A_217_521#_c_1312_n 0.00108565f $X=1.89 $Y=1.785 $X2=1.71
+ $Y2=0.755
cc_647 N_SN_M1015_g N_A_217_521#_c_1312_n 0.00495342f $X=1.925 $Y=0.85 $X2=1.71
+ $Y2=0.755
cc_648 N_SN_c_733_n N_A_217_521#_c_1315_n 0.00567928f $X=7.79 $Y=2.85 $X2=4.725
+ $Y2=2.285
cc_649 N_SN_c_704_n N_A_217_521#_c_1316_n 0.00675404f $X=1.89 $Y=1.785 $X2=1.68
+ $Y2=1.61
cc_650 N_SN_c_713_n N_A_217_521#_c_1316_n 0.00522003f $X=1.855 $Y=1.95 $X2=1.68
+ $Y2=1.61
cc_651 N_SN_c_717_n N_A_217_521#_c_1316_n 0.0184565f $X=1.71 $Y=1.95 $X2=1.68
+ $Y2=1.61
cc_652 N_SN_c_703_n N_A_217_521#_c_1319_n 0.00106582f $X=1.89 $Y=1.405 $X2=4.49
+ $Y2=1.37
cc_653 N_SN_c_704_n N_A_217_521#_c_1319_n 0.00569141f $X=1.89 $Y=1.785 $X2=4.49
+ $Y2=1.37
cc_654 N_SN_M1015_g N_A_217_521#_c_1319_n 0.00153565f $X=1.925 $Y=0.85 $X2=4.49
+ $Y2=1.37
cc_655 N_SN_c_717_n N_A_217_521#_c_1319_n 5.4793e-19 $X=1.71 $Y=1.95 $X2=4.49
+ $Y2=1.37
cc_656 N_SN_c_703_n N_A_217_521#_c_1320_n 4.80352e-19 $X=1.89 $Y=1.405 $X2=1.855
+ $Y2=1.37
cc_657 N_SN_c_704_n N_A_217_521#_c_1320_n 0.00104555f $X=1.89 $Y=1.785 $X2=1.855
+ $Y2=1.37
cc_658 N_SN_M1015_g N_A_217_521#_c_1320_n 5.56399e-19 $X=1.925 $Y=0.85 $X2=1.855
+ $Y2=1.37
cc_659 N_SN_c_717_n N_A_217_521#_c_1320_n 0.00302218f $X=1.71 $Y=1.95 $X2=1.855
+ $Y2=1.37
cc_660 N_SN_c_733_n N_A_704_89#_M1031_d 0.00393081f $X=7.79 $Y=2.85 $X2=6.81
+ $Y2=2.605
cc_661 N_SN_c_733_n N_A_704_89#_M1014_g 0.0128833f $X=7.79 $Y=2.85 $X2=4.195
+ $Y2=3.235
cc_662 N_SN_c_733_n N_A_704_89#_M1010_g 0.00850479f $X=7.79 $Y=2.85 $X2=5.345
+ $Y2=3.235
cc_663 N_SN_c_733_n N_A_704_89#_c_1494_n 0.0204742f $X=7.79 $Y=2.85 $X2=6.95
+ $Y2=2.955
cc_664 N_SN_c_716_n N_A_704_89#_c_1483_n 0.00393268f $X=7.937 $Y=2.482 $X2=7.22
+ $Y2=2.62
cc_665 N_SN_c_730_n N_A_704_89#_c_1499_n 0.00365476f $X=7.935 $Y=2.845 $X2=7.22
+ $Y2=2.705
cc_666 N_SN_c_733_n N_A_704_89#_c_1499_n 0.0140011f $X=7.79 $Y=2.85 $X2=7.22
+ $Y2=2.705
cc_667 SN N_A_704_89#_c_1499_n 0.00270579f $X=7.94 $Y=2.845 $X2=7.22 $Y2=2.705
cc_668 N_SN_c_733_n N_A_1246_89#_M1029_g 0.0101037f $X=7.79 $Y=2.85 $X2=6.305
+ $Y2=3.235
cc_669 N_SN_c_733_n N_A_1246_89#_c_1689_n 0.00210214f $X=7.79 $Y=2.85 $X2=6.365
+ $Y2=1.71
cc_670 N_SN_M1004_g N_A_1246_89#_c_1690_n 0.00700354f $X=8.045 $Y=0.85 $X2=8.26
+ $Y2=0.755
cc_671 N_SN_M1019_g N_A_1246_89#_c_1693_n 8.82637e-19 $X=8.115 $Y=3.235 $X2=8.76
+ $Y2=3.295
cc_672 N_SN_c_714_n N_A_1246_89#_c_1693_n 0.0024079f $X=8.02 $Y=1.775 $X2=8.76
+ $Y2=3.295
cc_673 N_SN_c_716_n N_A_1246_89#_c_1693_n 0.00705921f $X=7.937 $Y=2.482 $X2=8.76
+ $Y2=3.295
cc_674 N_SN_c_718_n N_A_1246_89#_c_1693_n 0.00488332f $X=8.02 $Y=1.775 $X2=8.76
+ $Y2=3.295
cc_675 N_SN_c_719_n N_A_1246_89#_c_1693_n 0.0122081f $X=7.937 $Y=2.395 $X2=8.76
+ $Y2=3.295
cc_676 SN N_A_1246_89#_c_1693_n 0.00504458f $X=7.94 $Y=2.845 $X2=8.76 $Y2=3.295
cc_677 N_SN_M1004_g N_A_1246_89#_c_1694_n 0.0039039f $X=8.045 $Y=0.85 $X2=8.845
+ $Y2=1.71
cc_678 N_SN_c_714_n N_A_1246_89#_c_1694_n 0.00231499f $X=8.02 $Y=1.775 $X2=8.845
+ $Y2=1.71
cc_679 N_SN_c_718_n N_A_1246_89#_c_1694_n 0.00799131f $X=8.02 $Y=1.775 $X2=8.845
+ $Y2=1.71
cc_680 N_SN_c_719_n N_A_1246_89#_c_1696_n 0.00416618f $X=7.937 $Y=2.395
+ $X2=7.165 $Y2=2.482
cc_681 N_SN_c_733_n N_A_1246_89#_c_1696_n 0.0715704f $X=7.79 $Y=2.85 $X2=7.165
+ $Y2=2.482
cc_682 N_SN_c_714_n N_A_1246_89#_c_1698_n 0.00639634f $X=8.02 $Y=1.775 $X2=9.235
+ $Y2=1.71
cc_683 N_SN_c_718_n N_A_1246_89#_c_1698_n 0.0201609f $X=8.02 $Y=1.775 $X2=9.235
+ $Y2=1.71
cc_684 N_SN_c_719_n N_A_1246_89#_c_1698_n 9.1164e-19 $X=7.937 $Y=2.395 $X2=9.235
+ $Y2=1.71
cc_685 N_SN_c_733_n N_A_1246_89#_c_1700_n 0.0272012f $X=7.79 $Y=2.85 $X2=6.515
+ $Y2=2.48
cc_686 N_SN_c_733_n N_A_1084_115#_M1010_d 0.0046196f $X=7.79 $Y=2.85 $X2=5.42
+ $Y2=2.605
cc_687 N_SN_M1004_g N_A_1084_115#_c_1883_n 0.00627778f $X=8.045 $Y=0.85
+ $X2=7.505 $Y2=2.15
cc_688 N_SN_M1019_g N_A_1084_115#_c_1883_n 0.00402616f $X=8.115 $Y=3.235
+ $X2=7.505 $Y2=2.15
cc_689 N_SN_c_714_n N_A_1084_115#_c_1883_n 0.0141258f $X=8.02 $Y=1.775 $X2=7.505
+ $Y2=2.15
cc_690 N_SN_c_718_n N_A_1084_115#_c_1883_n 6.29389e-19 $X=8.02 $Y=1.775
+ $X2=7.505 $Y2=2.15
cc_691 N_SN_c_719_n N_A_1084_115#_c_1883_n 5.97554e-19 $X=7.937 $Y=2.395
+ $X2=7.505 $Y2=2.15
cc_692 N_SN_M1004_g N_A_1084_115#_c_1884_n 0.0574115f $X=8.045 $Y=0.85 $X2=7.685
+ $Y2=1.21
cc_693 N_SN_c_716_n N_A_1084_115#_M1033_g 0.00419378f $X=7.937 $Y=2.482
+ $X2=7.685 $Y2=3.235
cc_694 N_SN_c_733_n N_A_1084_115#_M1033_g 0.0103641f $X=7.79 $Y=2.85 $X2=7.685
+ $Y2=3.235
cc_695 SN N_A_1084_115#_M1033_g 0.00222077f $X=7.94 $Y=2.845 $X2=7.685 $Y2=3.235
cc_696 N_SN_M1019_g N_A_1084_115#_c_1890_n 0.0610015f $X=8.115 $Y=3.235
+ $X2=7.685 $Y2=2.285
cc_697 N_SN_c_719_n N_A_1084_115#_c_1890_n 0.00419378f $X=7.937 $Y=2.395
+ $X2=7.685 $Y2=2.285
cc_698 N_SN_c_733_n N_A_1084_115#_c_1890_n 0.00208293f $X=7.79 $Y=2.85 $X2=7.685
+ $Y2=2.285
cc_699 N_SN_c_733_n N_A_1084_115#_c_1941_n 0.0259947f $X=7.79 $Y=2.85 $X2=5.475
+ $Y2=2.705
cc_700 N_SN_c_733_n N_A_1084_115#_c_1942_n 0.0139251f $X=7.79 $Y=2.85 $X2=5.15
+ $Y2=2.705
cc_701 N_SN_c_733_n N_A_1084_115#_c_1911_n 0.0334018f $X=7.79 $Y=2.85 $X2=5.645
+ $Y2=3.295
cc_702 N_SN_M1004_g N_A_1084_115#_c_1893_n 0.00226691f $X=8.045 $Y=0.85
+ $X2=7.595 $Y2=1.37
cc_703 N_SN_c_714_n N_A_1084_115#_c_1893_n 0.00139113f $X=8.02 $Y=1.775
+ $X2=7.595 $Y2=1.37
cc_704 N_SN_c_718_n N_A_1084_115#_c_1893_n 0.018479f $X=8.02 $Y=1.775 $X2=7.595
+ $Y2=1.37
cc_705 N_SN_c_719_n N_A_1084_115#_c_1893_n 0.0357198f $X=7.937 $Y=2.395
+ $X2=7.595 $Y2=1.37
cc_706 N_SN_c_733_n N_A_1084_115#_c_1893_n 0.00460427f $X=7.79 $Y=2.85 $X2=7.595
+ $Y2=1.37
cc_707 N_SN_M1004_g N_A_1084_115#_c_1904_n 0.00271237f $X=8.045 $Y=0.85
+ $X2=7.595 $Y2=1.37
cc_708 N_SN_c_732_n N_A_300_521#_M1000_d 0.00346218f $X=1.71 $Y=2.777 $X2=1.5
+ $Y2=2.605
cc_709 N_SN_c_733_n N_A_300_521#_M1027_d 0.00640134f $X=7.79 $Y=2.85 $X2=2.36
+ $Y2=2.605
cc_710 N_SN_M1024_g N_A_300_521#_c_2146_n 0.0135899f $X=1.855 $Y=3.235 $X2=2.415
+ $Y2=3.19
cc_711 N_SN_c_732_n N_A_300_521#_c_2146_n 0.0169389f $X=1.71 $Y=2.777 $X2=2.415
+ $Y2=3.19
cc_712 N_SN_c_733_n N_A_300_521#_c_2146_n 0.0164002f $X=7.79 $Y=2.85 $X2=2.415
+ $Y2=3.19
cc_713 N_SN_c_742_n N_A_300_521#_c_2146_n 0.00951546f $X=2.195 $Y=2.85 $X2=2.415
+ $Y2=3.19
cc_714 N_SN_c_732_n N_A_300_521#_c_2159_n 0.00659638f $X=1.71 $Y=2.777 $X2=1.725
+ $Y2=3.19
cc_715 N_SN_c_733_n A_662_521# 0.00813565f $X=7.79 $Y=2.85 $X2=3.31 $Y2=2.605
cc_716 N_SN_c_733_n A_854_521# 0.0162713f $X=7.79 $Y=2.85 $X2=4.27 $Y2=2.605
cc_717 N_SN_c_733_n A_1012_521# 0.00813565f $X=7.79 $Y=2.85 $X2=5.06 $Y2=2.605
cc_718 N_SN_c_733_n A_1204_521# 0.0157244f $X=7.79 $Y=2.85 $X2=6.02 $Y2=2.605
cc_719 N_SN_c_733_n N_A_1469_521#_M1033_s 0.00825332f $X=7.79 $Y=2.85 $X2=7.345
+ $Y2=2.605
cc_720 N_SN_M1019_g N_A_1469_521#_c_2174_n 0.0161914f $X=8.115 $Y=3.235
+ $X2=8.245 $Y2=3.185
cc_721 N_SN_c_730_n N_A_1469_521#_c_2174_n 0.00931248f $X=7.935 $Y=2.845
+ $X2=8.245 $Y2=3.185
cc_722 N_SN_c_733_n N_A_1469_521#_c_2174_n 0.00818864f $X=7.79 $Y=2.85 $X2=8.245
+ $Y2=3.185
cc_723 SN N_A_1469_521#_c_2174_n 0.010847f $X=7.94 $Y=2.845 $X2=8.245 $Y2=3.185
cc_724 N_SN_c_733_n N_A_1469_521#_c_2184_n 0.008614f $X=7.79 $Y=2.85 $X2=7.555
+ $Y2=3.185
cc_725 N_A_432_424#_c_902_n N_D_M1005_g 0.0123483f $X=3.71 $Y=1.285 $X2=3.235
+ $Y2=0.85
cc_726 N_A_432_424#_c_906_n N_D_M1028_g 0.00596171f $X=2.685 $Y=2.285 $X2=3.235
+ $Y2=3.235
cc_727 N_A_432_424#_c_907_n N_D_M1028_g 0.00737998f $X=2.77 $Y=2.62 $X2=3.235
+ $Y2=3.235
cc_728 N_A_432_424#_c_920_n N_D_M1028_g 0.0178646f $X=3.725 $Y=2.705 $X2=3.235
+ $Y2=3.235
cc_729 N_A_432_424#_c_902_n N_D_c_1010_n 0.00207628f $X=3.71 $Y=1.285 $X2=3.295
+ $Y2=1.74
cc_730 N_A_432_424#_c_902_n N_D_c_1011_n 0.0086486f $X=3.71 $Y=1.285 $X2=3.295
+ $Y2=1.74
cc_731 N_A_432_424#_c_902_n D 0.00200799f $X=3.71 $Y=1.285 $X2=3.295 $Y2=1.74
cc_732 N_A_432_424#_c_920_n N_CK_M1018_g 0.0141124f $X=3.725 $Y=2.705 $X2=3.595
+ $Y2=3.235
cc_733 N_A_432_424#_c_924_n N_CK_M1018_g 0.00642954f $X=3.895 $Y=2.955 $X2=3.595
+ $Y2=3.235
cc_734 N_A_432_424#_c_920_n N_CK_c_1045_n 0.00248712f $X=3.725 $Y=2.705
+ $X2=3.685 $Y2=2.285
cc_735 N_A_432_424#_c_902_n N_CK_c_1046_n 7.46335e-19 $X=3.71 $Y=1.285 $X2=4.135
+ $Y2=1.4
cc_736 N_A_432_424#_c_909_n N_CK_c_1046_n 0.00158678f $X=3.795 $Y=0.755
+ $X2=4.135 $Y2=1.4
cc_737 N_A_432_424#_c_902_n N_CK_c_1047_n 9.05754e-19 $X=3.71 $Y=1.285 $X2=4.135
+ $Y2=1.235
cc_738 N_A_432_424#_c_908_n N_CK_c_1047_n 0.00464203f $X=3.795 $Y=1.2 $X2=4.135
+ $Y2=1.235
cc_739 N_A_432_424#_c_909_n N_CK_c_1047_n 0.00243799f $X=3.795 $Y=0.755
+ $X2=4.135 $Y2=1.235
cc_740 N_A_432_424#_c_902_n N_CK_c_1061_n 0.00160862f $X=3.71 $Y=1.285 $X2=4.05
+ $Y2=2.11
cc_741 N_A_432_424#_c_920_n N_CK_c_1061_n 0.00810069f $X=3.725 $Y=2.705 $X2=4.05
+ $Y2=2.11
cc_742 N_A_432_424#_c_902_n N_CK_c_1062_n 0.00989572f $X=3.71 $Y=1.285 $X2=4.135
+ $Y2=1.4
cc_743 N_A_432_424#_c_909_n N_CK_c_1062_n 5.01691e-19 $X=3.795 $Y=0.755
+ $X2=4.135 $Y2=1.4
cc_744 N_A_432_424#_c_902_n N_CK_c_1067_n 0.00263105f $X=3.71 $Y=1.285 $X2=3.655
+ $Y2=2.11
cc_745 N_A_432_424#_c_920_n N_CK_c_1067_n 0.0102995f $X=3.725 $Y=2.705 $X2=3.655
+ $Y2=2.11
cc_746 N_A_432_424#_c_920_n N_CK_c_1069_n 0.00596172f $X=3.725 $Y=2.705 $X2=5.74
+ $Y2=2.11
cc_747 N_A_432_424#_c_920_n N_CK_c_1070_n 0.00225232f $X=3.725 $Y=2.705 $X2=3.8
+ $Y2=2.11
cc_748 N_A_432_424#_M1003_g N_A_217_521#_c_1312_n 8.95606e-19 $X=2.285 $Y=0.85
+ $X2=1.71 $Y2=0.755
cc_749 N_A_432_424#_c_901_n N_A_217_521#_c_1312_n 0.00949364f $X=2.295 $Y=2.2
+ $X2=1.71 $Y2=0.755
cc_750 N_A_432_424#_c_905_n N_A_217_521#_c_1312_n 0.00488587f $X=2.38 $Y=1.285
+ $X2=1.71 $Y2=0.755
cc_751 N_A_432_424#_M1003_g N_A_217_521#_c_1319_n 8.36391e-19 $X=2.285 $Y=0.85
+ $X2=4.49 $Y2=1.37
cc_752 N_A_432_424#_c_901_n N_A_217_521#_c_1319_n 0.0151086f $X=2.295 $Y=2.2
+ $X2=4.49 $Y2=1.37
cc_753 N_A_432_424#_c_902_n N_A_217_521#_c_1319_n 0.0579231f $X=3.71 $Y=1.285
+ $X2=4.49 $Y2=1.37
cc_754 N_A_432_424#_c_905_n N_A_217_521#_c_1319_n 0.00475107f $X=2.38 $Y=1.285
+ $X2=4.49 $Y2=1.37
cc_755 N_A_432_424#_c_909_n N_A_217_521#_c_1319_n 8.84716e-19 $X=3.795 $Y=0.755
+ $X2=4.49 $Y2=1.37
cc_756 N_A_432_424#_c_901_n N_A_217_521#_c_1320_n 6.43795e-19 $X=2.295 $Y=2.2
+ $X2=1.855 $Y2=1.37
cc_757 N_A_432_424#_c_905_n N_A_217_521#_c_1320_n 6.84883e-19 $X=2.38 $Y=1.285
+ $X2=1.855 $Y2=1.37
cc_758 N_A_432_424#_c_902_n N_A_704_89#_c_1460_n 0.0022787f $X=3.71 $Y=1.285
+ $X2=3.595 $Y2=1.205
cc_759 N_A_432_424#_c_908_n N_A_704_89#_c_1460_n 0.00432939f $X=3.795 $Y=1.2
+ $X2=3.595 $Y2=1.205
cc_760 N_A_432_424#_c_909_n N_A_704_89#_c_1460_n 0.00116801f $X=3.795 $Y=0.755
+ $X2=3.595 $Y2=1.205
cc_761 N_A_432_424#_c_902_n N_A_704_89#_c_1463_n 0.00333286f $X=3.71 $Y=1.285
+ $X2=3.715 $Y2=1.775
cc_762 N_A_432_424#_c_920_n N_A_704_89#_c_1464_n 6.56088e-19 $X=3.725 $Y=2.705
+ $X2=4.12 $Y2=1.85
cc_763 N_A_432_424#_c_920_n N_A_704_89#_M1014_g 0.0029243f $X=3.725 $Y=2.705
+ $X2=4.195 $Y2=3.235
cc_764 N_A_432_424#_c_924_n N_A_704_89#_M1014_g 0.00642954f $X=3.895 $Y=2.955
+ $X2=4.195 $Y2=3.235
cc_765 N_A_432_424#_c_902_n N_A_704_89#_c_1473_n 0.00993421f $X=3.71 $Y=1.285
+ $X2=3.715 $Y2=1.28
cc_766 N_A_432_424#_M1027_g N_A_300_521#_c_2146_n 0.014647f $X=2.285 $Y=3.235
+ $X2=2.415 $Y2=3.19
cc_767 N_A_432_424#_c_900_n N_A_300_521#_c_2146_n 3.89774e-19 $X=2.295 $Y=2.285
+ $X2=2.415 $Y2=3.19
cc_768 N_A_432_424#_c_901_n N_A_300_521#_c_2146_n 0.00153613f $X=2.295 $Y=2.2
+ $X2=2.415 $Y2=3.19
cc_769 N_A_432_424#_c_920_n A_662_521# 0.00529859f $X=3.725 $Y=2.705 $X2=3.31
+ $Y2=2.605
cc_770 N_D_M1028_g N_CK_c_1045_n 0.11342f $X=3.235 $Y=3.235 $X2=3.685 $Y2=2.285
cc_771 N_D_c_1011_n N_CK_c_1062_n 0.00479659f $X=3.295 $Y=1.74 $X2=4.135 $Y2=1.4
cc_772 D N_CK_c_1062_n 0.00555005f $X=3.295 $Y=1.74 $X2=4.135 $Y2=1.4
cc_773 N_D_M1028_g N_CK_c_1067_n 0.00566966f $X=3.235 $Y=3.235 $X2=3.655
+ $Y2=2.11
cc_774 N_D_M1028_g N_CK_c_1070_n 0.00542304f $X=3.235 $Y=3.235 $X2=3.8 $Y2=2.11
cc_775 D N_CK_c_1070_n 0.00375733f $X=3.295 $Y=1.74 $X2=3.8 $Y2=2.11
cc_776 N_D_M1005_g N_A_217_521#_c_1319_n 0.00303372f $X=3.235 $Y=0.85 $X2=4.49
+ $Y2=1.37
cc_777 N_D_c_1010_n N_A_217_521#_c_1319_n 7.9412e-19 $X=3.295 $Y=1.74 $X2=4.49
+ $Y2=1.37
cc_778 N_D_c_1011_n N_A_217_521#_c_1319_n 0.00111625f $X=3.295 $Y=1.74 $X2=4.49
+ $Y2=1.37
cc_779 D N_A_217_521#_c_1319_n 0.0353362f $X=3.295 $Y=1.74 $X2=4.49 $Y2=1.37
cc_780 N_D_M1005_g N_A_704_89#_c_1460_n 0.0567053f $X=3.235 $Y=0.85 $X2=3.595
+ $Y2=1.205
cc_781 N_D_M1005_g N_A_704_89#_c_1463_n 0.00932846f $X=3.235 $Y=0.85 $X2=3.715
+ $Y2=1.775
cc_782 N_D_c_1010_n N_A_704_89#_c_1463_n 0.0214858f $X=3.295 $Y=1.74 $X2=3.715
+ $Y2=1.775
cc_783 N_D_c_1011_n N_A_704_89#_c_1463_n 0.00166174f $X=3.295 $Y=1.74 $X2=3.715
+ $Y2=1.775
cc_784 D N_A_704_89#_c_1463_n 0.00338565f $X=3.295 $Y=1.74 $X2=3.715 $Y2=1.775
cc_785 N_D_M1028_g N_A_704_89#_c_1465_n 9.71193e-19 $X=3.235 $Y=3.235 $X2=3.79
+ $Y2=1.85
cc_786 D N_A_704_89#_c_1465_n 4.62757e-19 $X=3.295 $Y=1.74 $X2=3.79 $Y2=1.85
cc_787 N_CK_c_1047_n N_A_217_521#_M1020_g 0.0347751f $X=4.135 $Y=1.235 $X2=4.555
+ $Y2=0.85
cc_788 N_CK_c_1062_n N_A_217_521#_M1020_g 0.00109085f $X=4.135 $Y=1.4 $X2=4.555
+ $Y2=0.85
cc_789 N_CK_c_1050_n N_A_217_521#_c_1300_n 0.0343274f $X=5.405 $Y=1.4 $X2=4.91
+ $Y2=1.4
cc_790 N_CK_c_1046_n N_A_217_521#_c_1302_n 0.0347751f $X=4.135 $Y=1.4 $X2=4.63
+ $Y2=1.4
cc_791 N_CK_c_1069_n N_A_217_521#_c_1303_n 0.00765556f $X=5.74 $Y=2.11 $X2=4.91
+ $Y2=2.285
cc_792 N_CK_c_1069_n N_A_217_521#_c_1304_n 0.00673865f $X=5.74 $Y=2.11 $X2=4.63
+ $Y2=2.285
cc_793 N_CK_c_1051_n N_A_217_521#_M1023_g 0.0343274f $X=5.405 $Y=1.235 $X2=4.985
+ $Y2=0.85
cc_794 N_CK_c_1063_n N_A_217_521#_M1023_g 3.67139e-19 $X=5.405 $Y=1.4 $X2=4.985
+ $Y2=0.85
cc_795 N_CK_c_1046_n N_A_217_521#_c_1315_n 8.1208e-19 $X=4.135 $Y=1.4 $X2=4.725
+ $Y2=2.285
cc_796 N_CK_c_1061_n N_A_217_521#_c_1315_n 0.00402252f $X=4.05 $Y=2.11 $X2=4.725
+ $Y2=2.285
cc_797 N_CK_c_1062_n N_A_217_521#_c_1315_n 0.0202707f $X=4.135 $Y=1.4 $X2=4.725
+ $Y2=2.285
cc_798 N_CK_c_1069_n N_A_217_521#_c_1315_n 0.0206843f $X=5.74 $Y=2.11 $X2=4.725
+ $Y2=2.285
cc_799 N_CK_c_1046_n N_A_217_521#_c_1317_n 6.279e-19 $X=4.135 $Y=1.4 $X2=4.725
+ $Y2=1.4
cc_800 N_CK_c_1062_n N_A_217_521#_c_1317_n 0.00643639f $X=4.135 $Y=1.4 $X2=4.725
+ $Y2=1.4
cc_801 N_CK_c_1069_n N_A_217_521#_c_1317_n 0.00102309f $X=5.74 $Y=2.11 $X2=4.725
+ $Y2=1.4
cc_802 N_CK_c_1046_n N_A_217_521#_c_1319_n 0.00383333f $X=4.135 $Y=1.4 $X2=4.49
+ $Y2=1.37
cc_803 N_CK_c_1061_n N_A_217_521#_c_1319_n 0.0043165f $X=4.05 $Y=2.11 $X2=4.49
+ $Y2=1.37
cc_804 N_CK_c_1062_n N_A_217_521#_c_1319_n 0.0148598f $X=4.135 $Y=1.4 $X2=4.49
+ $Y2=1.37
cc_805 N_CK_c_1067_n N_A_217_521#_c_1319_n 8.37938e-19 $X=3.655 $Y=2.11 $X2=4.49
+ $Y2=1.37
cc_806 N_CK_c_1070_n N_A_217_521#_c_1319_n 0.0126162f $X=3.8 $Y=2.11 $X2=4.49
+ $Y2=1.37
cc_807 N_CK_c_1046_n N_A_217_521#_c_1372_n 3.26623e-19 $X=4.135 $Y=1.4 $X2=4.635
+ $Y2=1.37
cc_808 N_CK_c_1062_n N_A_217_521#_c_1372_n 0.00141649f $X=4.135 $Y=1.4 $X2=4.635
+ $Y2=1.37
cc_809 N_CK_c_1069_n N_A_217_521#_c_1372_n 0.0129652f $X=5.74 $Y=2.11 $X2=4.635
+ $Y2=1.37
cc_810 N_CK_c_1047_n N_A_704_89#_c_1460_n 0.01713f $X=4.135 $Y=1.235 $X2=3.595
+ $Y2=1.205
cc_811 N_CK_c_1062_n N_A_704_89#_c_1463_n 0.00602582f $X=4.135 $Y=1.4 $X2=3.715
+ $Y2=1.775
cc_812 N_CK_c_1046_n N_A_704_89#_c_1464_n 0.0183472f $X=4.135 $Y=1.4 $X2=4.12
+ $Y2=1.85
cc_813 N_CK_c_1062_n N_A_704_89#_c_1464_n 0.00665821f $X=4.135 $Y=1.4 $X2=4.12
+ $Y2=1.85
cc_814 N_CK_c_1069_n N_A_704_89#_c_1464_n 0.00549601f $X=5.74 $Y=2.11 $X2=4.12
+ $Y2=1.85
cc_815 N_CK_c_1045_n N_A_704_89#_c_1465_n 0.012591f $X=3.685 $Y=2.285 $X2=3.79
+ $Y2=1.85
cc_816 N_CK_c_1061_n N_A_704_89#_c_1465_n 0.00756374f $X=4.05 $Y=2.11 $X2=3.79
+ $Y2=1.85
cc_817 N_CK_c_1067_n N_A_704_89#_c_1465_n 0.00154604f $X=3.655 $Y=2.11 $X2=3.79
+ $Y2=1.85
cc_818 N_CK_c_1070_n N_A_704_89#_c_1465_n 0.00130179f $X=3.8 $Y=2.11 $X2=3.79
+ $Y2=1.85
cc_819 N_CK_M1018_g N_A_704_89#_M1014_g 0.0334679f $X=3.595 $Y=3.235 $X2=4.195
+ $Y2=3.235
cc_820 N_CK_c_1045_n N_A_704_89#_M1014_g 0.014942f $X=3.685 $Y=2.285 $X2=4.195
+ $Y2=3.235
cc_821 N_CK_c_1061_n N_A_704_89#_M1014_g 0.00849934f $X=4.05 $Y=2.11 $X2=4.195
+ $Y2=3.235
cc_822 N_CK_c_1062_n N_A_704_89#_M1014_g 0.00368559f $X=4.135 $Y=1.4 $X2=4.195
+ $Y2=3.235
cc_823 N_CK_c_1067_n N_A_704_89#_M1014_g 0.00148098f $X=3.655 $Y=2.11 $X2=4.195
+ $Y2=3.235
cc_824 N_CK_c_1069_n N_A_704_89#_M1014_g 0.00937774f $X=5.74 $Y=2.11 $X2=4.195
+ $Y2=3.235
cc_825 N_CK_c_1069_n N_A_704_89#_c_1467_n 0.00615595f $X=5.74 $Y=2.11 $X2=5.27
+ $Y2=1.85
cc_826 N_CK_M1002_g N_A_704_89#_M1010_g 0.0334711f $X=5.945 $Y=3.235 $X2=5.345
+ $Y2=3.235
cc_827 N_CK_c_1054_n N_A_704_89#_M1010_g 0.0138379f $X=5.855 $Y=2.285 $X2=5.345
+ $Y2=3.235
cc_828 N_CK_c_1063_n N_A_704_89#_M1010_g 0.00305863f $X=5.405 $Y=1.4 $X2=5.345
+ $Y2=3.235
cc_829 N_CK_c_1065_n N_A_704_89#_M1010_g 0.00692515f $X=5.49 $Y=2.11 $X2=5.345
+ $Y2=3.235
cc_830 N_CK_c_1068_n N_A_704_89#_M1010_g 8.92314e-19 $X=5.885 $Y=2.11 $X2=5.345
+ $Y2=3.235
cc_831 N_CK_c_1069_n N_A_704_89#_M1010_g 0.00496221f $X=5.74 $Y=2.11 $X2=5.345
+ $Y2=3.235
cc_832 N_CK_c_1054_n N_A_704_89#_c_1469_n 0.0199895f $X=5.855 $Y=2.285 $X2=5.75
+ $Y2=1.85
cc_833 N_CK_c_1063_n N_A_704_89#_c_1469_n 0.00748489f $X=5.405 $Y=1.4 $X2=5.75
+ $Y2=1.85
cc_834 N_CK_c_1064_n N_A_704_89#_c_1469_n 0.00733892f $X=5.77 $Y=2.11 $X2=5.75
+ $Y2=1.85
cc_835 N_CK_c_1069_n N_A_704_89#_c_1469_n 0.00525796f $X=5.74 $Y=2.11 $X2=5.75
+ $Y2=1.85
cc_836 N_CK_c_1072_n N_A_704_89#_c_1469_n 0.00130143f $X=6.03 $Y=2.11 $X2=5.75
+ $Y2=1.85
cc_837 N_CK_c_1050_n N_A_704_89#_M1017_g 0.0130327f $X=5.405 $Y=1.4 $X2=5.945
+ $Y2=0.85
cc_838 N_CK_c_1051_n N_A_704_89#_M1017_g 0.0176417f $X=5.405 $Y=1.235 $X2=5.945
+ $Y2=0.85
cc_839 N_CK_c_1063_n N_A_704_89#_M1017_g 9.23153e-19 $X=5.405 $Y=1.4 $X2=5.945
+ $Y2=0.85
cc_840 N_CK_c_1046_n N_A_704_89#_c_1473_n 0.0216996f $X=4.135 $Y=1.4 $X2=3.715
+ $Y2=1.28
cc_841 N_CK_c_1047_n N_A_704_89#_c_1473_n 9.76811e-19 $X=4.135 $Y=1.235
+ $X2=3.715 $Y2=1.28
cc_842 N_CK_c_1067_n N_A_704_89#_c_1473_n 2.43077e-19 $X=3.655 $Y=2.11 $X2=3.715
+ $Y2=1.28
cc_843 N_CK_c_1062_n N_A_704_89#_c_1474_n 0.00568091f $X=4.135 $Y=1.4 $X2=4.195
+ $Y2=1.85
cc_844 N_CK_c_1050_n N_A_704_89#_c_1475_n 0.0183472f $X=5.405 $Y=1.4 $X2=5.345
+ $Y2=1.85
cc_845 N_CK_c_1063_n N_A_704_89#_c_1475_n 0.00436024f $X=5.405 $Y=1.4 $X2=5.345
+ $Y2=1.85
cc_846 N_CK_c_1050_n N_A_704_89#_c_1476_n 3.30686e-19 $X=5.405 $Y=1.4 $X2=5.885
+ $Y2=1.725
cc_847 N_CK_c_1063_n N_A_704_89#_c_1476_n 0.00322821f $X=5.405 $Y=1.4 $X2=5.885
+ $Y2=1.725
cc_848 N_CK_c_1068_n N_A_704_89#_c_1476_n 0.00140833f $X=5.885 $Y=2.11 $X2=5.885
+ $Y2=1.725
cc_849 N_CK_c_1054_n N_A_704_89#_c_1477_n 7.52731e-19 $X=5.855 $Y=2.285
+ $X2=5.885 $Y2=1.725
cc_850 N_CK_c_1063_n N_A_704_89#_c_1477_n 0.00807959f $X=5.405 $Y=1.4 $X2=5.885
+ $Y2=1.725
cc_851 N_CK_c_1064_n N_A_704_89#_c_1477_n 0.0026204f $X=5.77 $Y=2.11 $X2=5.885
+ $Y2=1.725
cc_852 N_CK_c_1068_n N_A_704_89#_c_1477_n 0.0107916f $X=5.885 $Y=2.11 $X2=5.885
+ $Y2=1.725
cc_853 N_CK_c_1072_n N_A_704_89#_c_1477_n 0.00184909f $X=6.03 $Y=2.11 $X2=5.885
+ $Y2=1.725
cc_854 N_CK_c_1055_n N_A_704_89#_c_1478_n 0.00734472f $X=6.762 $Y=1.205 $X2=6.95
+ $Y2=0.755
cc_855 N_CK_c_1060_n N_A_704_89#_c_1478_n 0.0107024f $X=6.762 $Y=1.355 $X2=6.95
+ $Y2=0.755
cc_856 N_CK_M1031_g N_A_704_89#_c_1494_n 0.0016169f $X=6.735 $Y=3.235 $X2=6.95
+ $Y2=2.955
cc_857 N_CK_c_1043_n N_A_704_89#_c_1483_n 0.00262756f $X=6.735 $Y=2.45 $X2=7.22
+ $Y2=2.62
cc_858 N_CK_M1031_g N_A_704_89#_c_1483_n 0.00391574f $X=6.735 $Y=3.235 $X2=7.22
+ $Y2=2.62
cc_859 N_CK_c_1044_n N_A_704_89#_c_1483_n 0.00464589f $X=6.79 $Y=2.12 $X2=7.22
+ $Y2=2.62
cc_860 N_CK_c_1066_n N_A_704_89#_c_1483_n 0.0277276f $X=6.88 $Y=2.11 $X2=7.22
+ $Y2=2.62
cc_861 CK N_A_704_89#_c_1483_n 0.00253999f $X=6.88 $Y=2.11 $X2=7.22 $Y2=2.62
cc_862 N_CK_c_1043_n N_A_704_89#_c_1484_n 0.00161723f $X=6.735 $Y=2.45 $X2=7.22
+ $Y2=1.717
cc_863 N_CK_c_1044_n N_A_704_89#_c_1484_n 0.00277593f $X=6.79 $Y=2.12 $X2=7.22
+ $Y2=1.717
cc_864 N_CK_c_1066_n N_A_704_89#_c_1484_n 0.00565404f $X=6.88 $Y=2.11 $X2=7.22
+ $Y2=1.717
cc_865 CK N_A_704_89#_c_1484_n 7.89423e-19 $X=6.88 $Y=2.11 $X2=7.22 $Y2=1.717
cc_866 N_CK_c_1043_n N_A_704_89#_c_1499_n 0.00233394f $X=6.735 $Y=2.45 $X2=7.22
+ $Y2=2.705
cc_867 N_CK_M1031_g N_A_704_89#_c_1499_n 0.00289158f $X=6.735 $Y=3.235 $X2=7.22
+ $Y2=2.705
cc_868 N_CK_c_1066_n N_A_704_89#_c_1499_n 0.00601669f $X=6.88 $Y=2.11 $X2=7.22
+ $Y2=2.705
cc_869 N_CK_c_1044_n N_A_704_89#_c_1485_n 0.00341708f $X=6.79 $Y=2.12 $X2=6.835
+ $Y2=1.725
cc_870 N_CK_c_1060_n N_A_704_89#_c_1485_n 2.68475e-19 $X=6.762 $Y=1.355
+ $X2=6.835 $Y2=1.725
cc_871 N_CK_c_1066_n N_A_704_89#_c_1485_n 6.06587e-19 $X=6.88 $Y=2.11 $X2=6.835
+ $Y2=1.725
cc_872 N_CK_c_1071_n N_A_704_89#_c_1485_n 0.0547764f $X=6.735 $Y=2.11 $X2=6.835
+ $Y2=1.725
cc_873 CK N_A_704_89#_c_1485_n 0.00873337f $X=6.88 $Y=2.11 $X2=6.835 $Y2=1.725
cc_874 N_CK_c_1063_n N_A_704_89#_c_1486_n 0.00792502f $X=5.405 $Y=1.4 $X2=6.05
+ $Y2=1.725
cc_875 N_CK_c_1068_n N_A_704_89#_c_1486_n 5.96993e-19 $X=5.885 $Y=2.11 $X2=6.05
+ $Y2=1.725
cc_876 N_CK_c_1069_n N_A_704_89#_c_1486_n 0.00217458f $X=5.74 $Y=2.11 $X2=6.05
+ $Y2=1.725
cc_877 N_CK_c_1071_n N_A_704_89#_c_1486_n 0.00175935f $X=6.735 $Y=2.11 $X2=6.05
+ $Y2=1.725
cc_878 N_CK_c_1072_n N_A_704_89#_c_1486_n 0.0283385f $X=6.03 $Y=2.11 $X2=6.05
+ $Y2=1.725
cc_879 N_CK_c_1043_n N_A_704_89#_c_1487_n 2.37666e-19 $X=6.735 $Y=2.45 $X2=6.95
+ $Y2=1.725
cc_880 N_CK_c_1044_n N_A_704_89#_c_1487_n 0.00133063f $X=6.79 $Y=2.12 $X2=6.95
+ $Y2=1.725
cc_881 N_CK_c_1066_n N_A_704_89#_c_1487_n 8.21587e-19 $X=6.88 $Y=2.11 $X2=6.95
+ $Y2=1.725
cc_882 CK N_A_704_89#_c_1487_n 0.018764f $X=6.88 $Y=2.11 $X2=6.95 $Y2=1.725
cc_883 N_CK_c_1044_n N_A_1246_89#_M1006_g 0.00751867f $X=6.79 $Y=2.12 $X2=6.305
+ $Y2=0.85
cc_884 N_CK_c_1055_n N_A_1246_89#_M1006_g 0.0242212f $X=6.762 $Y=1.205 $X2=6.305
+ $Y2=0.85
cc_885 N_CK_c_1043_n N_A_1246_89#_M1029_g 0.041784f $X=6.735 $Y=2.45 $X2=6.305
+ $Y2=3.235
cc_886 N_CK_c_1044_n N_A_1246_89#_M1029_g 0.0149738f $X=6.79 $Y=2.12 $X2=6.305
+ $Y2=3.235
cc_887 N_CK_c_1054_n N_A_1246_89#_M1029_g 0.112607f $X=5.855 $Y=2.285 $X2=6.305
+ $Y2=3.235
cc_888 N_CK_c_1066_n N_A_1246_89#_M1029_g 5.92505e-19 $X=6.88 $Y=2.11 $X2=6.305
+ $Y2=3.235
cc_889 N_CK_c_1068_n N_A_1246_89#_M1029_g 0.0026293f $X=5.885 $Y=2.11 $X2=6.305
+ $Y2=3.235
cc_890 N_CK_c_1071_n N_A_1246_89#_M1029_g 0.00324541f $X=6.735 $Y=2.11 $X2=6.305
+ $Y2=3.235
cc_891 N_CK_c_1072_n N_A_1246_89#_M1029_g 0.00113587f $X=6.03 $Y=2.11 $X2=6.305
+ $Y2=3.235
cc_892 N_CK_c_1044_n N_A_1246_89#_c_1677_n 0.0208734f $X=6.79 $Y=2.12 $X2=6.365
+ $Y2=1.71
cc_893 N_CK_c_1071_n N_A_1246_89#_c_1677_n 7.95823e-19 $X=6.735 $Y=2.11
+ $X2=6.365 $Y2=1.71
cc_894 N_CK_c_1043_n N_A_1246_89#_c_1689_n 0.00273823f $X=6.735 $Y=2.45
+ $X2=6.365 $Y2=1.71
cc_895 N_CK_c_1044_n N_A_1246_89#_c_1689_n 0.00577586f $X=6.79 $Y=2.12 $X2=6.365
+ $Y2=1.71
cc_896 N_CK_c_1054_n N_A_1246_89#_c_1689_n 0.00220493f $X=5.855 $Y=2.285
+ $X2=6.365 $Y2=1.71
cc_897 N_CK_c_1066_n N_A_1246_89#_c_1689_n 0.0147163f $X=6.88 $Y=2.11 $X2=6.365
+ $Y2=1.71
cc_898 N_CK_c_1068_n N_A_1246_89#_c_1689_n 0.0145499f $X=5.885 $Y=2.11 $X2=6.365
+ $Y2=1.71
cc_899 N_CK_c_1071_n N_A_1246_89#_c_1689_n 0.0139276f $X=6.735 $Y=2.11 $X2=6.365
+ $Y2=1.71
cc_900 N_CK_c_1072_n N_A_1246_89#_c_1689_n 0.00207022f $X=6.03 $Y=2.11 $X2=6.365
+ $Y2=1.71
cc_901 CK N_A_1246_89#_c_1689_n 0.00189954f $X=6.88 $Y=2.11 $X2=6.365 $Y2=1.71
cc_902 N_CK_c_1043_n N_A_1246_89#_c_1696_n 0.00430818f $X=6.735 $Y=2.45
+ $X2=7.165 $Y2=2.482
cc_903 N_CK_M1031_g N_A_1246_89#_c_1696_n 0.00423375f $X=6.735 $Y=3.235
+ $X2=7.165 $Y2=2.482
cc_904 N_CK_c_1066_n N_A_1246_89#_c_1696_n 0.00649534f $X=6.88 $Y=2.11 $X2=7.165
+ $Y2=2.482
cc_905 N_CK_c_1071_n N_A_1246_89#_c_1696_n 0.018682f $X=6.735 $Y=2.11 $X2=7.165
+ $Y2=2.482
cc_906 CK N_A_1246_89#_c_1696_n 0.0251859f $X=6.88 $Y=2.11 $X2=7.165 $Y2=2.482
cc_907 N_CK_c_1066_n N_A_1246_89#_c_1697_n 0.00118692f $X=6.88 $Y=2.11 $X2=7.305
+ $Y2=2.39
cc_908 CK N_A_1246_89#_c_1697_n 0.0191038f $X=6.88 $Y=2.11 $X2=7.305 $Y2=2.39
cc_909 N_CK_c_1043_n N_A_1246_89#_c_1700_n 4.87662e-19 $X=6.735 $Y=2.45
+ $X2=6.515 $Y2=2.48
cc_910 N_CK_M1031_g N_A_1246_89#_c_1700_n 3.89642e-19 $X=6.735 $Y=3.235
+ $X2=6.515 $Y2=2.48
cc_911 N_CK_c_1054_n N_A_1246_89#_c_1700_n 0.00409438f $X=5.855 $Y=2.285
+ $X2=6.515 $Y2=2.48
cc_912 N_CK_c_1066_n N_A_1246_89#_c_1700_n 8.0542e-19 $X=6.88 $Y=2.11 $X2=6.515
+ $Y2=2.48
cc_913 N_CK_c_1068_n N_A_1246_89#_c_1700_n 0.00250499f $X=5.885 $Y=2.11
+ $X2=6.515 $Y2=2.48
cc_914 N_CK_c_1071_n N_A_1246_89#_c_1700_n 0.0257812f $X=6.735 $Y=2.11 $X2=6.515
+ $Y2=2.48
cc_915 N_CK_c_1043_n N_A_1084_115#_c_1883_n 0.00731225f $X=6.735 $Y=2.45
+ $X2=7.505 $Y2=2.15
cc_916 N_CK_c_1044_n N_A_1084_115#_c_1883_n 0.00724311f $X=6.79 $Y=2.12
+ $X2=7.505 $Y2=2.15
cc_917 N_CK_c_1043_n N_A_1084_115#_M1033_g 5.00344e-19 $X=6.735 $Y=2.45
+ $X2=7.685 $Y2=3.235
cc_918 N_CK_c_1060_n N_A_1084_115#_c_1888_n 0.00724311f $X=6.762 $Y=1.355
+ $X2=7.685 $Y2=1.29
cc_919 N_CK_c_1050_n N_A_1084_115#_c_1891_n 0.00215979f $X=5.405 $Y=1.4
+ $X2=5.065 $Y2=1.37
cc_920 N_CK_c_1063_n N_A_1084_115#_c_1891_n 0.0548695f $X=5.405 $Y=1.4 $X2=5.065
+ $Y2=1.37
cc_921 N_CK_c_1065_n N_A_1084_115#_c_1891_n 0.0116464f $X=5.49 $Y=2.11 $X2=5.065
+ $Y2=1.37
cc_922 N_CK_c_1068_n N_A_1084_115#_c_1891_n 0.00640739f $X=5.885 $Y=2.11
+ $X2=5.065 $Y2=1.37
cc_923 N_CK_c_1069_n N_A_1084_115#_c_1891_n 0.020359f $X=5.74 $Y=2.11 $X2=5.065
+ $Y2=1.37
cc_924 N_CK_c_1072_n N_A_1084_115#_c_1891_n 5.47744e-19 $X=6.03 $Y=2.11
+ $X2=5.065 $Y2=1.37
cc_925 N_CK_M1002_g N_A_1084_115#_c_1941_n 0.00130117f $X=5.945 $Y=3.235
+ $X2=5.475 $Y2=2.705
cc_926 N_CK_c_1054_n N_A_1084_115#_c_1941_n 0.00248712f $X=5.855 $Y=2.285
+ $X2=5.475 $Y2=2.705
cc_927 N_CK_c_1064_n N_A_1084_115#_c_1941_n 0.00748399f $X=5.77 $Y=2.11
+ $X2=5.475 $Y2=2.705
cc_928 N_CK_c_1065_n N_A_1084_115#_c_1941_n 0.00323798f $X=5.49 $Y=2.11
+ $X2=5.475 $Y2=2.705
cc_929 N_CK_c_1068_n N_A_1084_115#_c_1941_n 0.00329042f $X=5.885 $Y=2.11
+ $X2=5.475 $Y2=2.705
cc_930 N_CK_c_1069_n N_A_1084_115#_c_1941_n 0.0125804f $X=5.74 $Y=2.11 $X2=5.475
+ $Y2=2.705
cc_931 N_CK_c_1072_n N_A_1084_115#_c_1941_n 4.61668e-19 $X=6.03 $Y=2.11
+ $X2=5.475 $Y2=2.705
cc_932 N_CK_M1002_g N_A_1084_115#_c_1911_n 0.00774456f $X=5.945 $Y=3.235
+ $X2=5.645 $Y2=3.295
cc_933 N_CK_c_1050_n N_A_1084_115#_c_1892_n 0.00114703f $X=5.405 $Y=1.4
+ $X2=5.745 $Y2=1.34
cc_934 N_CK_c_1051_n N_A_1084_115#_c_1892_n 0.00378955f $X=5.405 $Y=1.235
+ $X2=5.745 $Y2=1.34
cc_935 N_CK_c_1063_n N_A_1084_115#_c_1892_n 0.0125904f $X=5.405 $Y=1.4 $X2=5.745
+ $Y2=1.34
cc_936 N_CK_c_1064_n N_A_1084_115#_c_1892_n 0.00103909f $X=5.77 $Y=2.11
+ $X2=5.745 $Y2=1.34
cc_937 N_CK_c_1069_n N_A_1084_115#_c_1892_n 8.69566e-19 $X=5.74 $Y=2.11
+ $X2=5.745 $Y2=1.34
cc_938 N_CK_c_1044_n N_A_1084_115#_c_1893_n 4.42019e-19 $X=6.79 $Y=2.12
+ $X2=7.595 $Y2=1.37
cc_939 N_CK_c_1050_n N_A_1084_115#_c_1895_n 0.00183284f $X=5.405 $Y=1.4
+ $X2=5.645 $Y2=0.755
cc_940 N_CK_c_1051_n N_A_1084_115#_c_1895_n 0.00389012f $X=5.405 $Y=1.235
+ $X2=5.645 $Y2=0.755
cc_941 N_CK_c_1063_n N_A_1084_115#_c_1895_n 7.53857e-19 $X=5.405 $Y=1.4
+ $X2=5.645 $Y2=0.755
cc_942 N_CK_c_1050_n N_A_1084_115#_c_1898_n 0.00421189f $X=5.405 $Y=1.4 $X2=5.6
+ $Y2=1.37
cc_943 N_CK_c_1063_n N_A_1084_115#_c_1898_n 0.0127625f $X=5.405 $Y=1.4 $X2=5.6
+ $Y2=1.37
cc_944 N_CK_c_1064_n N_A_1084_115#_c_1898_n 0.00386167f $X=5.77 $Y=2.11 $X2=5.6
+ $Y2=1.37
cc_945 N_CK_c_1050_n N_A_1084_115#_c_1899_n 6.81488e-19 $X=5.405 $Y=1.4 $X2=5.21
+ $Y2=1.37
cc_946 N_CK_c_1063_n N_A_1084_115#_c_1899_n 0.0012142f $X=5.405 $Y=1.4 $X2=5.21
+ $Y2=1.37
cc_947 N_CK_c_1069_n N_A_1084_115#_c_1899_n 0.0128239f $X=5.74 $Y=2.11 $X2=5.21
+ $Y2=1.37
cc_948 N_CK_c_1044_n N_A_1084_115#_c_1900_n 0.00329792f $X=6.79 $Y=2.12 $X2=7.45
+ $Y2=1.37
cc_949 N_CK_c_1060_n N_A_1084_115#_c_1900_n 0.00383994f $X=6.762 $Y=1.355
+ $X2=7.45 $Y2=1.37
cc_950 N_CK_c_1050_n N_A_1084_115#_c_1903_n 5.48392e-19 $X=5.405 $Y=1.4 $X2=5.89
+ $Y2=1.37
cc_951 N_CK_c_1063_n N_A_1084_115#_c_1903_n 8.69968e-19 $X=5.405 $Y=1.4 $X2=5.89
+ $Y2=1.37
cc_952 N_A_217_521#_c_1319_n N_A_704_89#_c_1463_n 0.00256992f $X=4.49 $Y=1.37
+ $X2=3.715 $Y2=1.775
cc_953 N_A_217_521#_c_1319_n N_A_704_89#_c_1464_n 0.00290011f $X=4.49 $Y=1.37
+ $X2=4.12 $Y2=1.85
cc_954 N_A_217_521#_c_1304_n N_A_704_89#_M1014_g 0.115227f $X=4.63 $Y=2.285
+ $X2=4.195 $Y2=3.235
cc_955 N_A_217_521#_c_1315_n N_A_704_89#_M1014_g 0.00435172f $X=4.725 $Y=2.285
+ $X2=4.195 $Y2=3.235
cc_956 N_A_217_521#_c_1302_n N_A_704_89#_c_1467_n 0.0342442f $X=4.63 $Y=1.4
+ $X2=5.27 $Y2=1.85
cc_957 N_A_217_521#_c_1304_n N_A_704_89#_c_1467_n 0.0355605f $X=4.63 $Y=2.285
+ $X2=5.27 $Y2=1.85
cc_958 N_A_217_521#_c_1315_n N_A_704_89#_c_1467_n 0.0111197f $X=4.725 $Y=2.285
+ $X2=5.27 $Y2=1.85
cc_959 N_A_217_521#_c_1317_n N_A_704_89#_c_1467_n 8.22237e-19 $X=4.725 $Y=1.4
+ $X2=5.27 $Y2=1.85
cc_960 N_A_217_521#_c_1319_n N_A_704_89#_c_1467_n 0.00477469f $X=4.49 $Y=1.37
+ $X2=5.27 $Y2=1.85
cc_961 N_A_217_521#_c_1372_n N_A_704_89#_c_1467_n 3.93645e-19 $X=4.635 $Y=1.37
+ $X2=5.27 $Y2=1.85
cc_962 N_A_217_521#_c_1303_n N_A_704_89#_M1010_g 0.111657f $X=4.91 $Y=2.285
+ $X2=5.345 $Y2=3.235
cc_963 N_A_217_521#_M1009_g N_A_1084_115#_c_1891_n 9.36754e-19 $X=4.555 $Y=3.235
+ $X2=5.065 $Y2=1.37
cc_964 N_A_217_521#_c_1300_n N_A_1084_115#_c_1891_n 0.00625851f $X=4.91 $Y=1.4
+ $X2=5.065 $Y2=1.37
cc_965 N_A_217_521#_c_1303_n N_A_1084_115#_c_1891_n 0.00729195f $X=4.91 $Y=2.285
+ $X2=5.065 $Y2=1.37
cc_966 N_A_217_521#_M1023_g N_A_1084_115#_c_1891_n 0.00190765f $X=4.985 $Y=0.85
+ $X2=5.065 $Y2=1.37
cc_967 N_A_217_521#_M1012_g N_A_1084_115#_c_1891_n 0.00479454f $X=4.985 $Y=3.235
+ $X2=5.065 $Y2=1.37
cc_968 N_A_217_521#_c_1315_n N_A_1084_115#_c_1891_n 0.0700092f $X=4.725 $Y=2.285
+ $X2=5.065 $Y2=1.37
cc_969 N_A_217_521#_c_1317_n N_A_1084_115#_c_1891_n 0.0137157f $X=4.725 $Y=1.4
+ $X2=5.065 $Y2=1.37
cc_970 N_A_217_521#_c_1372_n N_A_1084_115#_c_1891_n 4.17564e-19 $X=4.635 $Y=1.37
+ $X2=5.065 $Y2=1.37
cc_971 N_A_217_521#_M1009_g N_A_1084_115#_c_1942_n 0.00100689f $X=4.555 $Y=3.235
+ $X2=5.15 $Y2=2.705
cc_972 N_A_217_521#_M1012_g N_A_1084_115#_c_1942_n 0.00751605f $X=4.985 $Y=3.235
+ $X2=5.15 $Y2=2.705
cc_973 N_A_217_521#_c_1300_n N_A_1084_115#_c_1899_n 0.00167673f $X=4.91 $Y=1.4
+ $X2=5.21 $Y2=1.37
cc_974 N_A_217_521#_M1023_g N_A_1084_115#_c_1899_n 5.96517e-19 $X=4.985 $Y=0.85
+ $X2=5.21 $Y2=1.37
cc_975 N_A_217_521#_c_1317_n N_A_1084_115#_c_1899_n 0.00121185f $X=4.725 $Y=1.4
+ $X2=5.21 $Y2=1.37
cc_976 N_A_217_521#_c_1372_n N_A_1084_115#_c_1899_n 0.0241344f $X=4.635 $Y=1.37
+ $X2=5.21 $Y2=1.37
cc_977 N_A_704_89#_M1017_g N_A_1246_89#_M1006_g 0.0477253f $X=5.945 $Y=0.85
+ $X2=6.305 $Y2=0.85
cc_978 N_A_704_89#_c_1476_n N_A_1246_89#_c_1677_n 0.0477253f $X=5.885 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_979 N_A_704_89#_c_1477_n N_A_1246_89#_c_1677_n 7.65216e-19 $X=5.885 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_980 N_A_704_89#_c_1484_n N_A_1246_89#_c_1677_n 5.63779e-19 $X=7.22 $Y=1.717
+ $X2=6.365 $Y2=1.71
cc_981 N_A_704_89#_c_1485_n N_A_1246_89#_c_1677_n 0.0032375f $X=6.835 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_982 N_A_704_89#_c_1486_n N_A_1246_89#_c_1677_n 9.33997e-19 $X=6.05 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_983 N_A_704_89#_c_1487_n N_A_1246_89#_c_1677_n 2.8797e-19 $X=6.95 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_984 N_A_704_89#_M1017_g N_A_1246_89#_c_1689_n 5.76765e-19 $X=5.945 $Y=0.85
+ $X2=6.365 $Y2=1.71
cc_985 N_A_704_89#_c_1476_n N_A_1246_89#_c_1689_n 0.0010529f $X=5.885 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_986 N_A_704_89#_c_1477_n N_A_1246_89#_c_1689_n 0.00843011f $X=5.885 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_987 N_A_704_89#_c_1478_n N_A_1246_89#_c_1689_n 0.00274567f $X=6.95 $Y=0.755
+ $X2=6.365 $Y2=1.71
cc_988 N_A_704_89#_c_1484_n N_A_1246_89#_c_1689_n 0.00391882f $X=7.22 $Y=1.717
+ $X2=6.365 $Y2=1.71
cc_989 N_A_704_89#_c_1485_n N_A_1246_89#_c_1689_n 0.012602f $X=6.835 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_990 N_A_704_89#_c_1486_n N_A_1246_89#_c_1689_n 0.0025776f $X=6.05 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_991 N_A_704_89#_c_1487_n N_A_1246_89#_c_1689_n 0.00157515f $X=6.95 $Y=1.725
+ $X2=6.365 $Y2=1.71
cc_992 N_A_704_89#_c_1483_n N_A_1246_89#_c_1696_n 0.0130526f $X=7.22 $Y=2.62
+ $X2=7.165 $Y2=2.482
cc_993 N_A_704_89#_c_1484_n N_A_1246_89#_c_1696_n 0.001994f $X=7.22 $Y=1.717
+ $X2=7.165 $Y2=2.482
cc_994 N_A_704_89#_c_1499_n N_A_1246_89#_c_1696_n 0.00626008f $X=7.22 $Y=2.705
+ $X2=7.165 $Y2=2.482
cc_995 N_A_704_89#_c_1487_n N_A_1246_89#_c_1696_n 0.00354883f $X=6.95 $Y=1.725
+ $X2=7.165 $Y2=2.482
cc_996 N_A_704_89#_c_1483_n N_A_1246_89#_c_1697_n 0.0150687f $X=7.22 $Y=2.62
+ $X2=7.305 $Y2=2.39
cc_997 N_A_704_89#_c_1484_n N_A_1246_89#_c_1697_n 3.31865e-19 $X=7.22 $Y=1.717
+ $X2=7.305 $Y2=2.39
cc_998 N_A_704_89#_c_1484_n N_A_1246_89#_c_1699_n 0.00676543f $X=7.22 $Y=1.717
+ $X2=7.375 $Y2=1.71
cc_999 N_A_704_89#_c_1487_n N_A_1246_89#_c_1699_n 0.0215891f $X=6.95 $Y=1.725
+ $X2=7.375 $Y2=1.71
cc_1000 N_A_704_89#_c_1483_n N_A_1084_115#_c_1883_n 0.00526325f $X=7.22 $Y=2.62
+ $X2=7.505 $Y2=2.15
cc_1001 N_A_704_89#_c_1484_n N_A_1084_115#_c_1883_n 0.00148649f $X=7.22 $Y=1.717
+ $X2=7.505 $Y2=2.15
cc_1002 N_A_704_89#_c_1487_n N_A_1084_115#_c_1883_n 2.21095e-19 $X=6.95 $Y=1.725
+ $X2=7.505 $Y2=2.15
cc_1003 N_A_704_89#_c_1478_n N_A_1084_115#_c_1884_n 0.00540908f $X=6.95 $Y=0.755
+ $X2=7.685 $Y2=1.21
cc_1004 N_A_704_89#_c_1494_n N_A_1084_115#_M1033_g 0.00491855f $X=6.95 $Y=2.955
+ $X2=7.685 $Y2=3.235
cc_1005 N_A_704_89#_c_1483_n N_A_1084_115#_M1033_g 0.00320908f $X=7.22 $Y=2.62
+ $X2=7.685 $Y2=3.235
cc_1006 N_A_704_89#_c_1499_n N_A_1084_115#_M1033_g 0.00330729f $X=7.22 $Y=2.705
+ $X2=7.685 $Y2=3.235
cc_1007 N_A_704_89#_c_1478_n N_A_1084_115#_c_1888_n 0.00358178f $X=6.95 $Y=0.755
+ $X2=7.685 $Y2=1.29
cc_1008 N_A_704_89#_c_1467_n N_A_1084_115#_c_1891_n 0.012215f $X=5.27 $Y=1.85
+ $X2=5.065 $Y2=1.37
cc_1009 N_A_704_89#_M1010_g N_A_1084_115#_c_1891_n 0.0104621f $X=5.345 $Y=3.235
+ $X2=5.065 $Y2=1.37
cc_1010 N_A_704_89#_c_1467_n N_A_1084_115#_c_1941_n 5.88705e-19 $X=5.27 $Y=1.85
+ $X2=5.475 $Y2=2.705
cc_1011 N_A_704_89#_M1010_g N_A_1084_115#_c_1941_n 0.0132272f $X=5.345 $Y=3.235
+ $X2=5.475 $Y2=2.705
cc_1012 N_A_704_89#_c_1469_n N_A_1084_115#_c_1941_n 6.306e-19 $X=5.75 $Y=1.85
+ $X2=5.475 $Y2=2.705
cc_1013 N_A_704_89#_M1010_g N_A_1084_115#_c_1911_n 0.00795444f $X=5.345 $Y=3.235
+ $X2=5.645 $Y2=3.295
cc_1014 N_A_704_89#_c_1476_n N_A_1084_115#_c_1892_n 0.00192187f $X=5.885
+ $Y=1.725 $X2=5.745 $Y2=1.34
cc_1015 N_A_704_89#_c_1477_n N_A_1084_115#_c_1892_n 0.00603136f $X=5.885
+ $Y=1.725 $X2=5.745 $Y2=1.34
cc_1016 N_A_704_89#_c_1486_n N_A_1084_115#_c_1892_n 3.56744e-19 $X=6.05 $Y=1.725
+ $X2=5.745 $Y2=1.34
cc_1017 N_A_704_89#_c_1478_n N_A_1084_115#_c_1893_n 0.00850247f $X=6.95 $Y=0.755
+ $X2=7.595 $Y2=1.37
cc_1018 N_A_704_89#_c_1483_n N_A_1084_115#_c_1893_n 0.0325734f $X=7.22 $Y=2.62
+ $X2=7.595 $Y2=1.37
cc_1019 N_A_704_89#_c_1484_n N_A_1084_115#_c_1893_n 0.0103463f $X=7.22 $Y=1.717
+ $X2=7.595 $Y2=1.37
cc_1020 N_A_704_89#_c_1487_n N_A_1084_115#_c_1893_n 5.67824e-19 $X=6.95 $Y=1.725
+ $X2=7.595 $Y2=1.37
cc_1021 N_A_704_89#_M1017_g N_A_1084_115#_c_1895_n 0.0118283f $X=5.945 $Y=0.85
+ $X2=5.645 $Y2=0.755
cc_1022 N_A_704_89#_c_1467_n N_A_1084_115#_c_1898_n 0.0015396f $X=5.27 $Y=1.85
+ $X2=5.6 $Y2=1.37
cc_1023 N_A_704_89#_c_1469_n N_A_1084_115#_c_1898_n 0.00243388f $X=5.75 $Y=1.85
+ $X2=5.6 $Y2=1.37
cc_1024 N_A_704_89#_c_1475_n N_A_1084_115#_c_1898_n 5.01668e-19 $X=5.345 $Y=1.85
+ $X2=5.6 $Y2=1.37
cc_1025 N_A_704_89#_c_1467_n N_A_1084_115#_c_1899_n 0.00117411f $X=5.27 $Y=1.85
+ $X2=5.21 $Y2=1.37
cc_1026 N_A_704_89#_M1017_g N_A_1084_115#_c_1900_n 0.00354979f $X=5.945 $Y=0.85
+ $X2=7.45 $Y2=1.37
cc_1027 N_A_704_89#_c_1478_n N_A_1084_115#_c_1900_n 0.017327f $X=6.95 $Y=0.755
+ $X2=7.45 $Y2=1.37
cc_1028 N_A_704_89#_c_1484_n N_A_1084_115#_c_1900_n 0.00762396f $X=7.22 $Y=1.717
+ $X2=7.45 $Y2=1.37
cc_1029 N_A_704_89#_c_1485_n N_A_1084_115#_c_1900_n 0.0680549f $X=6.835 $Y=1.725
+ $X2=7.45 $Y2=1.37
cc_1030 N_A_704_89#_c_1487_n N_A_1084_115#_c_1900_n 0.0234074f $X=6.95 $Y=1.725
+ $X2=7.45 $Y2=1.37
cc_1031 N_A_704_89#_M1017_g N_A_1084_115#_c_1903_n 0.00265988f $X=5.945 $Y=0.85
+ $X2=5.89 $Y2=1.37
cc_1032 N_A_704_89#_c_1476_n N_A_1084_115#_c_1903_n 0.00194236f $X=5.885
+ $Y=1.725 $X2=5.89 $Y2=1.37
cc_1033 N_A_704_89#_c_1477_n N_A_1084_115#_c_1903_n 0.00337066f $X=5.885
+ $Y=1.725 $X2=5.89 $Y2=1.37
cc_1034 N_A_704_89#_c_1486_n N_A_1084_115#_c_1903_n 0.0323443f $X=6.05 $Y=1.725
+ $X2=5.89 $Y2=1.37
cc_1035 N_A_704_89#_c_1478_n N_A_1084_115#_c_1904_n 0.00168079f $X=6.95 $Y=0.755
+ $X2=7.595 $Y2=1.37
cc_1036 N_A_704_89#_c_1494_n N_A_1469_521#_c_2171_n 0.0253961f $X=6.95 $Y=2.955
+ $X2=7.47 $Y2=3.295
cc_1037 N_A_704_89#_c_1494_n N_A_1469_521#_c_2184_n 0.00961556f $X=6.95 $Y=2.955
+ $X2=7.555 $Y2=3.185
cc_1038 N_A_1246_89#_c_1697_n N_A_1084_115#_c_1883_n 0.00498349f $X=7.305
+ $Y=2.39 $X2=7.505 $Y2=2.15
cc_1039 N_A_1246_89#_c_1698_n N_A_1084_115#_c_1883_n 0.00499408f $X=9.235
+ $Y=1.71 $X2=7.505 $Y2=2.15
cc_1040 N_A_1246_89#_c_1696_n N_A_1084_115#_M1033_g 0.00324314f $X=7.165
+ $Y=2.482 $X2=7.685 $Y2=3.235
cc_1041 N_A_1246_89#_c_1698_n N_A_1084_115#_c_1888_n 6.8924e-19 $X=9.235 $Y=1.71
+ $X2=7.685 $Y2=1.29
cc_1042 N_A_1246_89#_c_1696_n N_A_1084_115#_c_1890_n 0.00498349f $X=7.165
+ $Y=2.482 $X2=7.685 $Y2=2.285
cc_1043 N_A_1246_89#_c_1698_n N_A_1084_115#_c_1890_n 0.00207076f $X=9.235
+ $Y=1.71 $X2=7.685 $Y2=2.285
cc_1044 N_A_1246_89#_c_1690_n N_A_1084_115#_c_1893_n 0.0010677f $X=8.26 $Y=0.755
+ $X2=7.595 $Y2=1.37
cc_1045 N_A_1246_89#_c_1694_n N_A_1084_115#_c_1893_n 0.00830619f $X=8.845
+ $Y=1.71 $X2=7.595 $Y2=1.37
cc_1046 N_A_1246_89#_c_1697_n N_A_1084_115#_c_1893_n 0.0176387f $X=7.305 $Y=2.39
+ $X2=7.595 $Y2=1.37
cc_1047 N_A_1246_89#_c_1698_n N_A_1084_115#_c_1893_n 0.01645f $X=9.235 $Y=1.71
+ $X2=7.595 $Y2=1.37
cc_1048 N_A_1246_89#_M1006_g N_A_1084_115#_c_1900_n 0.00571159f $X=6.305 $Y=0.85
+ $X2=7.45 $Y2=1.37
cc_1049 N_A_1246_89#_c_1677_n N_A_1084_115#_c_1900_n 8.17219e-19 $X=6.365
+ $Y=1.71 $X2=7.45 $Y2=1.37
cc_1050 N_A_1246_89#_c_1689_n N_A_1084_115#_c_1900_n 0.00519268f $X=6.365
+ $Y=1.71 $X2=7.45 $Y2=1.37
cc_1051 N_A_1246_89#_c_1699_n N_A_1084_115#_c_1900_n 0.0206868f $X=7.375 $Y=1.71
+ $X2=7.45 $Y2=1.37
cc_1052 N_A_1246_89#_c_1690_n N_A_1084_115#_c_1904_n 0.00247064f $X=8.26
+ $Y=0.755 $X2=7.595 $Y2=1.37
cc_1053 N_A_1246_89#_c_1694_n N_A_1084_115#_c_1904_n 0.00385209f $X=8.845
+ $Y=1.71 $X2=7.595 $Y2=1.37
cc_1054 N_A_1246_89#_c_1698_n N_A_1084_115#_c_1904_n 0.027605f $X=9.235 $Y=1.71
+ $X2=7.595 $Y2=1.37
cc_1055 N_A_1246_89#_c_1680_n N_QN_M1008_g 0.0131322f $X=9.382 $Y=1.545
+ $X2=9.925 $Y2=0.85
cc_1056 N_A_1246_89#_c_1681_n N_QN_M1008_g 0.0230653f $X=9.47 $Y=1.23 $X2=9.925
+ $Y2=0.85
cc_1057 N_A_1246_89#_c_1695_n N_QN_M1008_g 4.79563e-19 $X=9.38 $Y=1.71 $X2=9.925
+ $Y2=0.85
cc_1058 N_A_1246_89#_c_1687_n N_QN_M1032_g 0.0102953f $X=9.47 $Y=2.375 $X2=9.925
+ $Y2=3.235
cc_1059 N_A_1246_89#_c_1688_n N_QN_M1032_g 0.021932f $X=9.47 $Y=2.525 $X2=9.925
+ $Y2=3.235
cc_1060 N_A_1246_89#_c_1679_n N_QN_c_2064_n 0.021196f $X=9.38 $Y=1.71 $X2=9.865
+ $Y2=1.915
cc_1061 N_A_1246_89#_c_1695_n N_QN_c_2064_n 3.0115e-19 $X=9.38 $Y=1.71 $X2=9.865
+ $Y2=1.915
cc_1062 N_A_1246_89#_c_1701_n N_QN_c_2064_n 4.60229e-19 $X=9.38 $Y=1.71
+ $X2=9.865 $Y2=1.915
cc_1063 N_A_1246_89#_c_1681_n N_QN_c_2065_n 0.00575865f $X=9.47 $Y=1.23 $X2=9.28
+ $Y2=0.755
cc_1064 N_A_1246_89#_c_1686_n N_QN_c_2065_n 0.00147419f $X=9.47 $Y=1.38 $X2=9.28
+ $Y2=0.755
cc_1065 N_A_1246_89#_c_1687_n N_QN_c_2069_n 0.00521938f $X=9.47 $Y=2.375
+ $X2=9.28 $Y2=2.48
cc_1066 N_A_1246_89#_c_1688_n N_QN_c_2069_n 0.00631458f $X=9.47 $Y=2.525
+ $X2=9.28 $Y2=2.48
cc_1067 N_A_1246_89#_c_1693_n N_QN_c_2069_n 0.0610685f $X=8.76 $Y=3.295 $X2=9.28
+ $Y2=2.48
cc_1068 N_A_1246_89#_c_1680_n N_QN_c_2070_n 0.00473974f $X=9.382 $Y=1.545
+ $X2=9.78 $Y2=1.37
cc_1069 N_A_1246_89#_c_1686_n N_QN_c_2070_n 0.0130902f $X=9.47 $Y=1.38 $X2=9.78
+ $Y2=1.37
cc_1070 N_A_1246_89#_c_1695_n N_QN_c_2070_n 0.0110497f $X=9.38 $Y=1.71 $X2=9.78
+ $Y2=1.37
cc_1071 N_A_1246_89#_c_1701_n N_QN_c_2070_n 0.00387586f $X=9.38 $Y=1.71 $X2=9.78
+ $Y2=1.37
cc_1072 N_A_1246_89#_c_1679_n N_QN_c_2072_n 0.00308111f $X=9.38 $Y=1.71
+ $X2=9.365 $Y2=1.37
cc_1073 N_A_1246_89#_c_1695_n N_QN_c_2072_n 0.0120703f $X=9.38 $Y=1.71 $X2=9.365
+ $Y2=1.37
cc_1074 N_A_1246_89#_c_1698_n N_QN_c_2072_n 0.0010572f $X=9.235 $Y=1.71
+ $X2=9.365 $Y2=1.37
cc_1075 N_A_1246_89#_c_1701_n N_QN_c_2072_n 0.00336135f $X=9.38 $Y=1.71
+ $X2=9.365 $Y2=1.37
cc_1076 N_A_1246_89#_c_1687_n N_QN_c_2073_n 0.0152835f $X=9.47 $Y=2.375 $X2=9.78
+ $Y2=2.285
cc_1077 N_A_1246_89#_c_1688_n N_QN_c_2073_n 0.00248624f $X=9.47 $Y=2.525
+ $X2=9.78 $Y2=2.285
cc_1078 N_A_1246_89#_c_1695_n N_QN_c_2073_n 0.00426371f $X=9.38 $Y=1.71 $X2=9.78
+ $Y2=2.285
cc_1079 N_A_1246_89#_c_1701_n N_QN_c_2073_n 0.00253233f $X=9.38 $Y=1.71 $X2=9.78
+ $Y2=2.285
cc_1080 N_A_1246_89#_c_1679_n N_QN_c_2074_n 0.00265611f $X=9.38 $Y=1.71
+ $X2=9.365 $Y2=2.285
cc_1081 N_A_1246_89#_c_1693_n N_QN_c_2074_n 0.00826781f $X=8.76 $Y=3.295
+ $X2=9.365 $Y2=2.285
cc_1082 N_A_1246_89#_c_1695_n N_QN_c_2074_n 0.00471962f $X=9.38 $Y=1.71
+ $X2=9.365 $Y2=2.285
cc_1083 N_A_1246_89#_c_1698_n N_QN_c_2074_n 9.40773e-19 $X=9.235 $Y=1.71
+ $X2=9.365 $Y2=2.285
cc_1084 N_A_1246_89#_c_1701_n N_QN_c_2074_n 0.00140341f $X=9.38 $Y=1.71
+ $X2=9.365 $Y2=2.285
cc_1085 N_A_1246_89#_c_1679_n N_QN_c_2075_n 0.00216137f $X=9.38 $Y=1.71
+ $X2=9.865 $Y2=1.915
cc_1086 N_A_1246_89#_c_1680_n N_QN_c_2075_n 0.00323473f $X=9.382 $Y=1.545
+ $X2=9.865 $Y2=1.915
cc_1087 N_A_1246_89#_c_1687_n N_QN_c_2075_n 0.00226435f $X=9.47 $Y=2.375
+ $X2=9.865 $Y2=1.915
cc_1088 N_A_1246_89#_c_1695_n N_QN_c_2075_n 0.00987106f $X=9.38 $Y=1.71
+ $X2=9.865 $Y2=1.915
cc_1089 N_A_1246_89#_c_1701_n N_QN_c_2075_n 0.00377439f $X=9.38 $Y=1.71
+ $X2=9.865 $Y2=1.915
cc_1090 N_A_1246_89#_c_1688_n QN 0.00718989f $X=9.47 $Y=2.525 $X2=9.285 $Y2=2.48
cc_1091 N_A_1246_89#_c_1693_n QN 0.00721908f $X=8.76 $Y=3.295 $X2=9.285 $Y2=2.48
cc_1092 N_A_1246_89#_c_1695_n QN 0.00359685f $X=9.38 $Y=1.71 $X2=9.285 $Y2=2.48
cc_1093 N_A_1246_89#_c_1701_n QN 0.00842298f $X=9.38 $Y=1.71 $X2=9.285 $Y2=2.48
cc_1094 N_A_1084_115#_c_1941_n A_1012_521# 0.00185532f $X=5.475 $Y=2.705
+ $X2=5.06 $Y2=2.605
cc_1095 N_A_1084_115#_c_1942_n A_1012_521# 5.47801e-19 $X=5.15 $Y=2.705 $X2=5.06
+ $Y2=2.605
cc_1096 N_A_1084_115#_M1033_g N_A_1469_521#_c_2174_n 0.0138653f $X=7.685
+ $Y=3.235 $X2=8.245 $Y2=3.185
cc_1097 N_A_1084_115#_c_1893_n N_A_1469_521#_c_2174_n 0.00107647f $X=7.595
+ $Y=1.37 $X2=8.245 $Y2=3.185
cc_1098 N_A_1084_115#_c_1890_n N_A_1469_521#_c_2184_n 0.00265163f $X=7.685
+ $Y=2.285 $X2=7.555 $Y2=3.185
cc_1099 N_A_1084_115#_c_1893_n N_A_1469_521#_c_2184_n 6.20558e-19 $X=7.595
+ $Y=1.37 $X2=7.555 $Y2=3.185
cc_1100 N_QN_M1032_g N_Q_c_2195_n 0.00224668f $X=9.925 $Y=3.235 $X2=10.14
+ $Y2=2.85
cc_1101 N_QN_M1008_g N_Q_c_2193_n 0.0330655f $X=9.925 $Y=0.85 $X2=10.255
+ $Y2=2.525
cc_1102 N_QN_c_2070_n N_Q_c_2193_n 0.0111776f $X=9.78 $Y=1.37 $X2=10.255
+ $Y2=2.525
cc_1103 N_QN_c_2073_n N_Q_c_2193_n 0.0111776f $X=9.78 $Y=2.285 $X2=10.255
+ $Y2=2.525
cc_1104 N_QN_c_2075_n N_Q_c_2193_n 0.0438362f $X=9.865 $Y=1.915 $X2=10.255
+ $Y2=2.525
cc_1105 N_QN_M1032_g N_Q_c_2199_n 0.00495318f $X=9.925 $Y=3.235 $X2=10.255
+ $Y2=2.61
cc_1106 N_QN_M1032_g Q 0.0101636f $X=9.925 $Y=3.235 $X2=10.14 $Y2=2.85
cc_1107 N_QN_c_2073_n Q 0.00228117f $X=9.78 $Y=2.285 $X2=10.14 $Y2=2.85
