* File: sky130_osu_sc_18T_ms__nand2_1.pex.spice
* Created: Thu Oct 29 17:30:30 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_1%GND 1 12 14 21 24 27
r25 24 27 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r26 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r27 12 19 4.26217 $w=1.7e-07 $l=2.14243e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=1.05 $Y2=0.305
r28 12 14 3.29607 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=0.965 $Y2=0.152
r29 12 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r30 12 14 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r31 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_1%VDD 1 2 13 17 23 30 32 35
r20 35 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r21 32 35 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r22 30 39 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r23 27 39 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r24 27 29 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r25 23 26 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r26 21 30 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.035 $Y2=6.507
r27 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r28 17 20 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r29 15 29 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r30 15 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r31 13 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r32 13 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r33 2 26 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r34 2 23 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r35 1 20 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r36 1 17 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_1%A 3 7 10 15 16
r31 16 18 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.685
+ $X2=0.367 $Y2=2.85
r32 16 17 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.685
+ $X2=0.367 $Y2=2.52
r33 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.685 $X2=0.32 $Y2=2.685
r34 12 15 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=2.685
r35 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r36 7 18 889.649 $w=1.5e-07 $l=1.735e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.85
r37 3 17 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.52
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_1%B 3 7 11 13 17 19
c38 3 0 1.57512e-19 $X=0.835 $Y=1.075
r39 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.06 $Y=2.96
+ $X2=1.06 $Y2=2.96
r40 14 19 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.06 $Y=2.305
+ $X2=1.06 $Y2=2.96
r41 13 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=2.22
+ $X2=1.06 $Y2=2.305
r42 11 22 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.055
r43 10 13 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.915 $Y=2.22
+ $X2=1.06 $Y2=2.22
r44 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=2.22 $X2=0.915 $Y2=2.22
r45 5 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.385
+ $X2=0.905 $Y2=2.22
r46 5 7 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.905 $Y=2.385
+ $X2=0.905 $Y2=4.585
r47 3 22 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__NAND2_1%Y 1 2 7 8 12 19 20 23
c41 12 0 4.69618e-20 $X=0.68 $Y=2.35
c42 8 0 1.57512e-19 $X=0.405 $Y=1.48
r43 30 32 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r44 20 30 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=0.69 $Y=2.59
+ $X2=0.69 $Y2=3.455
r45 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.59
+ $X2=0.69 $Y2=2.59
r46 16 23 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.26 $Y=1.48
+ $X2=0.26 $Y2=0.825
r47 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.48
+ $X2=0.26 $Y2=1.48
r48 10 19 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.475
+ $X2=0.69 $Y2=2.59
r49 10 12 0.12036 $w=1.7e-07 $l=1.25e-07 $layer=MET1_cond $X=0.69 $Y=2.475
+ $X2=0.69 $Y2=2.35
r50 9 12 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=0.69 $Y=1.565
+ $X2=0.69 $Y2=2.35
r51 8 15 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=1.48
+ $X2=0.26 $Y2=1.48
r52 7 9 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=1.48
+ $X2=0.69 $Y2=1.565
r53 7 8 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=1.48 $X2=0.405
+ $Y2=1.48
r54 2 32 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r55 2 30 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r56 1 23 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

