* File: sky130_osu_sc_15T_ms__inv_10.pex.spice
* Created: Fri Nov 12 14:43:46 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__INV_10%GND 1 2 3 4 5 6 67 71 73 80 82 89 91 98
+ 100 107 109 117 132 134
r138 132 134 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r139 115 117 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.56 $Y2=0.865
r140 109 115 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.475
+ $Y=0.152 $X2=4.56 $Y2=0.305
r141 105 107 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.865
r142 101 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r143 96 125 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r144 96 98 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.865
r145 92 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r146 91 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r147 87 124 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r148 87 89 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.865
r149 83 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r150 82 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r151 78 123 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r152 78 80 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.865
r153 73 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r154 69 71 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r155 67 134 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r156 67 132 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r157 67 105 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.7 $Y2=0.305
r158 67 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.615 $Y2=0.152
r159 67 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.785 $Y2=0.152
r160 67 69 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r161 67 74 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r162 67 109 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.475 $Y2=0.152
r163 67 110 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=3.785 $Y2=0.152
r164 67 100 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r165 67 101 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r166 67 91 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r167 67 92 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r168 67 82 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r169 67 83 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r170 67 73 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r171 67 74 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r172 6 117 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.575 $X2=4.56 $Y2=0.865
r173 5 107 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.865
r174 4 98 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.865
r175 3 89 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.865
r176 2 80 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r177 1 71 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__INV_10%VDD 1 2 3 4 5 6 53 57 61 67 71 77 81 87
+ 91 97 101 108 121 125
r96 121 125 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=4.42 $Y2=5.397
r97 113 121 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r98 108 111 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.56 $Y=3.205
+ $X2=4.56 $Y2=4.565
r99 106 111 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.56 $Y=5.245
+ $X2=4.56 $Y2=4.565
r100 104 125 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=5.36
+ $X2=4.42 $Y2=5.36
r101 102 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=5.397
+ $X2=3.7 $Y2=5.397
r102 102 104 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=5.397
+ $X2=4.42 $Y2=5.397
r103 101 106 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.475 $Y=5.397
+ $X2=4.56 $Y2=5.245
r104 101 104 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.475 $Y=5.397
+ $X2=4.42 $Y2=5.397
r105 97 100 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.7 $Y=3.205
+ $X2=3.7 $Y2=4.565
r106 95 119 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.7 $Y=5.245
+ $X2=3.7 $Y2=5.397
r107 95 100 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=5.245
+ $X2=3.7 $Y2=4.565
r108 92 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=2.84 $Y2=5.397
r109 92 94 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=3.06 $Y2=5.397
r110 91 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.7 $Y2=5.397
r111 91 94 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.06 $Y2=5.397
r112 87 90 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.205
+ $X2=2.84 $Y2=4.565
r113 85 117 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=5.397
r114 85 90 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.565
r115 82 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r116 82 84 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r117 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.397
r118 81 84 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r119 77 80 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.205
+ $X2=1.98 $Y2=4.565
r120 75 116 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r121 75 80 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.565
r122 72 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r123 72 74 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r124 71 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r125 71 74 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r126 67 70 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=3.205
+ $X2=1.12 $Y2=4.565
r127 65 115 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r128 65 70 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r129 62 113 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r130 62 64 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r131 61 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r132 61 64 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r133 57 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r134 55 113 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r135 55 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r136 53 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=5.245 $X2=4.42 $Y2=5.33
r137 53 119 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r138 53 94 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r139 53 84 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r140 53 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r141 53 64 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r142 53 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r143 6 111 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.825 $X2=4.56 $Y2=4.565
r144 6 108 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.825 $X2=4.56 $Y2=3.205
r145 5 100 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=4.565
r146 5 97 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=3.205
r147 4 90 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.565
r148 4 87 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.205
r149 3 80 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.565
r150 3 77 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.205
r151 2 70 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r152 2 67 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.205
r153 1 60 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r154 1 57 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__INV_10%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 45 47 49 50 52 53 55 57 59 60 62 63 65 67 69
+ 70 72 73 75 77 79 80 82 83 85 87 89 90 92 93 95 97 99 100 102 103 105 106 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 127 129 131
+ 134
c289 90 0 1.33323e-19 $X=3.915 $Y=2.7
c290 87 0 1.33323e-19 $X=3.915 $Y=1.44
c291 80 0 1.33323e-19 $X=3.485 $Y=2.7
c292 77 0 1.33323e-19 $X=3.485 $Y=1.44
c293 70 0 1.33323e-19 $X=3.055 $Y=2.7
c294 67 0 1.33323e-19 $X=3.055 $Y=1.44
c295 60 0 1.33323e-19 $X=2.625 $Y=2.7
c296 57 0 1.33323e-19 $X=2.625 $Y=1.44
c297 50 0 1.33323e-19 $X=2.195 $Y=2.7
c298 45 0 1.33323e-19 $X=2.195 $Y=1.44
c299 38 0 1.33323e-19 $X=1.765 $Y=2.7
c300 35 0 1.33323e-19 $X=1.765 $Y=1.44
c301 28 0 1.33323e-19 $X=1.335 $Y=2.7
c302 25 0 1.33323e-19 $X=1.335 $Y=1.44
c303 18 0 1.33323e-19 $X=0.905 $Y=2.7
c304 15 0 1.33323e-19 $X=0.905 $Y=1.44
r305 134 137 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=3.065
+ $X2=0.405 $Y2=3.07
r306 129 131 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.045
+ $X2=0.535 $Y2=2.045
r307 127 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r308 125 129 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.405 $Y2=2.045
r309 125 127 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.32 $Y2=3.07
r310 105 131 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.045 $X2=0.535 $Y2=2.045
r311 105 107 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=2.21
r312 105 106 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=1.88
r313 100 102 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=4.345 $Y=2.7
+ $X2=4.345 $Y2=3.825
r314 97 99 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.345 $Y=1.44
+ $X2=4.345 $Y2=0.945
r315 96 124 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=2.625
+ $X2=3.915 $Y2=2.625
r316 95 100 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=2.625
+ $X2=4.345 $Y2=2.7
r317 95 96 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=2.625
+ $X2=3.99 $Y2=2.625
r318 94 123 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.515
+ $X2=3.915 $Y2=1.515
r319 93 97 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=1.515
+ $X2=4.345 $Y2=1.44
r320 93 94 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.515
+ $X2=3.99 $Y2=1.515
r321 90 124 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=2.7
+ $X2=3.915 $Y2=2.625
r322 90 92 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.915 $Y=2.7
+ $X2=3.915 $Y2=3.825
r323 87 123 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=1.44
+ $X2=3.915 $Y2=1.515
r324 87 89 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.915 $Y=1.44
+ $X2=3.915 $Y2=0.945
r325 86 122 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.625
+ $X2=3.485 $Y2=2.625
r326 85 124 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.625
+ $X2=3.915 $Y2=2.625
r327 85 86 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.625
+ $X2=3.56 $Y2=2.625
r328 84 121 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.515
+ $X2=3.485 $Y2=1.515
r329 83 123 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.515
+ $X2=3.915 $Y2=1.515
r330 83 84 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.515
+ $X2=3.56 $Y2=1.515
r331 80 122 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=2.625
r332 80 82 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=3.825
r333 77 121 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.485 $Y2=1.515
r334 77 79 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.485 $Y2=0.945
r335 76 120 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.625
+ $X2=3.055 $Y2=2.625
r336 75 122 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.485 $Y2=2.625
r337 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.13 $Y2=2.625
r338 74 119 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.055 $Y2=1.515
r339 73 121 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.515
+ $X2=3.485 $Y2=1.515
r340 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.515
+ $X2=3.13 $Y2=1.515
r341 70 120 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=2.625
r342 70 72 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=3.825
r343 67 119 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=1.515
r344 67 69 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=0.945
r345 66 118 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.625
+ $X2=2.625 $Y2=2.625
r346 65 120 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=3.055 $Y2=2.625
r347 65 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=2.7 $Y2=2.625
r348 64 117 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.625 $Y2=1.515
r349 63 119 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=3.055 $Y2=1.515
r350 63 64 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=2.7 $Y2=1.515
r351 60 118 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=2.625
r352 60 62 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r353 57 117 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=1.515
r354 57 59 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=0.945
r355 56 116 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r356 55 118 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.625
r357 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r358 54 115 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.515
+ $X2=2.195 $Y2=1.515
r359 53 117 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.625 $Y2=1.515
r360 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.27 $Y2=1.515
r361 50 116 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=2.625
r362 50 52 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r363 49 116 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.55
+ $X2=2.195 $Y2=2.625
r364 48 115 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.59
+ $X2=2.195 $Y2=1.515
r365 48 49 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.59
+ $X2=2.195 $Y2=2.55
r366 45 115 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.44
+ $X2=2.195 $Y2=1.515
r367 45 47 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.195 $Y=1.44
+ $X2=2.195 $Y2=0.945
r368 44 114 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r369 43 116 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r370 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r371 42 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.515
+ $X2=1.765 $Y2=1.515
r372 41 115 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.515
+ $X2=2.195 $Y2=1.515
r373 41 42 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.515
+ $X2=1.84 $Y2=1.515
r374 38 114 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r375 38 40 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r376 35 113 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.44
+ $X2=1.765 $Y2=1.515
r377 35 37 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.765 $Y=1.44
+ $X2=1.765 $Y2=0.945
r378 34 112 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.625
+ $X2=1.335 $Y2=2.625
r379 33 114 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r380 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.41 $Y2=2.625
r381 32 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.335 $Y2=1.515
r382 31 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.765 $Y2=1.515
r383 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.41 $Y2=1.515
r384 28 112 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=2.625
r385 28 30 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r386 25 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.44
+ $X2=1.335 $Y2=1.515
r387 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.335 $Y=1.44
+ $X2=1.335 $Y2=0.945
r388 24 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.625
+ $X2=0.905 $Y2=2.625
r389 23 112 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.625
+ $X2=1.335 $Y2=2.625
r390 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.625
+ $X2=0.98 $Y2=2.625
r391 22 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.515
+ $X2=0.905 $Y2=1.515
r392 21 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=1.335 $Y2=1.515
r393 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=0.98 $Y2=1.515
r394 18 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.7
+ $X2=0.905 $Y2=2.625
r395 18 20 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=2.7
+ $X2=0.905 $Y2=3.825
r396 15 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.44
+ $X2=0.905 $Y2=1.515
r397 15 17 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.905 $Y=1.44
+ $X2=0.905 $Y2=0.945
r398 14 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.625
+ $X2=0.475 $Y2=2.625
r399 13 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.625
+ $X2=0.905 $Y2=2.625
r400 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.625
+ $X2=0.55 $Y2=2.625
r401 12 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.515
+ $X2=0.475 $Y2=1.515
r402 11 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.515
+ $X2=0.905 $Y2=1.515
r403 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.515
+ $X2=0.55 $Y2=1.515
r404 8 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.7
+ $X2=0.475 $Y2=2.625
r405 8 10 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.475 $Y=2.7
+ $X2=0.475 $Y2=3.825
r406 7 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.55
+ $X2=0.475 $Y2=2.625
r407 7 107 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.55
+ $X2=0.475 $Y2=2.21
r408 4 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.59
+ $X2=0.475 $Y2=1.515
r409 4 106 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.59
+ $X2=0.475 $Y2=1.88
r410 1 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=1.515
r411 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__INV_10%Y 1 2 3 4 5 11 12 13 14 15 42 48 56 62
+ 70 76 84 90 98 104 111 112 114 116 118 121 122 123 124 125 127 128 129 130 131
+ 133 134 135 136 137 138 139
c213 139 0 1.33323e-19 $X=4.13 $Y=2.585
c214 138 0 1.33323e-19 $X=4.13 $Y=1.335
c215 137 0 2.66647e-19 $X=3.415 $Y=2.7
c216 135 0 2.66647e-19 $X=3.415 $Y=1.22
c217 131 0 2.66647e-19 $X=2.555 $Y=2.7
c218 129 0 2.66647e-19 $X=2.555 $Y=1.22
c219 125 0 2.66647e-19 $X=1.695 $Y=2.7
c220 123 0 2.66647e-19 $X=1.695 $Y=1.22
c221 112 0 1.33323e-19 $X=0.69 $Y=2.585
c222 111 0 1.33323e-19 $X=0.69 $Y=1.335
r223 139 159 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=2.585
+ $X2=4.13 $Y2=2.7
r224 138 157 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.335
+ $X2=4.13 $Y2=1.22
r225 138 139 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=4.13 $Y=1.335
+ $X2=4.13 $Y2=2.585
r226 137 155 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=2.7
+ $X2=3.27 $Y2=2.7
r227 136 159 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=2.7
+ $X2=4.13 $Y2=2.7
r228 136 137 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=2.7
+ $X2=3.415 $Y2=2.7
r229 135 153 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=1.22
+ $X2=3.27 $Y2=1.22
r230 134 157 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=1.22
+ $X2=4.13 $Y2=1.22
r231 134 135 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=1.22
+ $X2=3.415 $Y2=1.22
r232 133 155 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.585
+ $X2=3.27 $Y2=2.7
r233 132 153 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=1.22
r234 132 133 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=2.585
r235 131 151 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.7
+ $X2=2.41 $Y2=2.7
r236 130 155 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.7
+ $X2=3.27 $Y2=2.7
r237 130 131 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.7
+ $X2=2.555 $Y2=2.7
r238 129 149 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.22
+ $X2=2.41 $Y2=1.22
r239 128 153 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=3.27 $Y2=1.22
r240 128 129 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=2.555 $Y2=1.22
r241 127 151 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.585
+ $X2=2.41 $Y2=2.7
r242 126 149 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r243 126 127 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.585
r244 125 147 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.7
+ $X2=1.55 $Y2=2.7
r245 124 151 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.7
+ $X2=2.41 $Y2=2.7
r246 124 125 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.7
+ $X2=1.695 $Y2=2.7
r247 123 145 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r248 122 149 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r249 122 123 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r250 121 147 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.585
+ $X2=1.55 $Y2=2.7
r251 120 145 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r252 120 121 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=2.585
r253 119 143 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.7
+ $X2=0.69 $Y2=2.7
r254 118 147 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.7
+ $X2=1.55 $Y2=2.7
r255 118 119 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.7
+ $X2=0.835 $Y2=2.7
r256 117 141 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.22
+ $X2=0.69 $Y2=1.22
r257 116 145 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.22
+ $X2=1.55 $Y2=1.22
r258 116 117 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.22
+ $X2=0.835 $Y2=1.22
r259 112 143 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=2.7
r260 112 114 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=1.94
r261 111 141 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.22
r262 111 114 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.94
r263 107 109 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.13 $Y=3.205
+ $X2=4.13 $Y2=4.565
r264 104 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=2.7
+ $X2=4.13 $Y2=2.7
r265 104 107 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.13 $Y=2.7
+ $X2=4.13 $Y2=3.205
r266 101 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=1.22
+ $X2=4.13 $Y2=1.22
r267 98 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.13 $Y=0.865
+ $X2=4.13 $Y2=1.22
r268 93 95 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.27 $Y=3.205
+ $X2=3.27 $Y2=4.565
r269 90 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.7
+ $X2=3.27 $Y2=2.7
r270 90 93 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.27 $Y=2.7
+ $X2=3.27 $Y2=3.205
r271 87 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.22
+ $X2=3.27 $Y2=1.22
r272 84 87 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.27 $Y=0.865
+ $X2=3.27 $Y2=1.22
r273 79 81 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.205
+ $X2=2.41 $Y2=4.565
r274 76 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.7
+ $X2=2.41 $Y2=2.7
r275 76 79 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.41 $Y=2.7
+ $X2=2.41 $Y2=3.205
r276 73 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r277 70 73 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.41 $Y=0.865
+ $X2=2.41 $Y2=1.22
r278 65 67 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.205
+ $X2=1.55 $Y2=4.565
r279 62 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.7
+ $X2=1.55 $Y2=2.7
r280 62 65 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.55 $Y=2.7
+ $X2=1.55 $Y2=3.205
r281 59 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r282 56 59 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.55 $Y=0.865
+ $X2=1.55 $Y2=1.22
r283 51 53 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r284 48 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=2.7
r285 48 51 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=3.205
r286 45 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.22
+ $X2=0.69 $Y2=1.22
r287 42 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.69 $Y=0.865
+ $X2=0.69 $Y2=1.22
r288 15 109 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.825 $X2=4.13 $Y2=4.565
r289 15 107 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.825 $X2=4.13 $Y2=3.205
r290 14 95 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=4.565
r291 14 93 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=3.205
r292 13 81 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.565
r293 13 79 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.205
r294 12 67 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.565
r295 12 65 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.205
r296 11 53 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r297 11 51 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r298 5 98 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.865
r299 4 84 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.865
r300 3 70 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.865
r301 2 56 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.865
r302 1 42 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

