* File: sky130_osu_sc_15T_ls__tbufi_1.pex.spice
* Created: Fri Nov 12 14:59:54 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__TBUFI_1%GND 1 17 19 26 35 38
r38 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r39 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r40 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r41 24 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.865
r42 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r43 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r44 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r45 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r46 1 26 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TBUFI_1%VDD 1 13 15 21 27 31 34
r21 31 34 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r22 27 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r23 25 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r24 25 27 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397 $X2=1.02
+ $Y2=5.397
r25 21 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=3.545
+ $X2=0.69 $Y2=4.565
r26 19 29 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r27 19 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.565
r28 15 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r29 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r30 13 27 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r31 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r32 1 24 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r33 1 21 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.545
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TBUFI_1%OE 2 3 5 6 8 9 11 14 19 22 29 32
c65 29 0 2.60266e-19 $X=0.69 $Y=1.59
r66 26 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.705
+ $X2=0.69 $Y2=1.59
r67 26 32 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=0.69 $Y=1.705
+ $X2=0.69 $Y2=2.585
r68 22 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.59
+ $X2=0.69 $Y2=1.59
r69 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.59 $X2=0.69 $Y2=1.59
r70 12 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.675
+ $X2=0.475 $Y2=2.675
r71 9 19 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.905 $Y=1.39
+ $X2=0.69 $Y2=1.572
r72 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.905 $Y=1.39
+ $X2=0.905 $Y2=0.945
r73 6 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=2.675
r74 6 8 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=3.825
r75 3 19 46.4709 $w=2.23e-07 $l=2.92156e-07 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.69 $Y2=1.572
r76 3 5 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.475 $Y=1.39
+ $X2=0.475 $Y2=0.945
r77 2 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.6 $X2=0.27
+ $Y2=2.675
r78 1 3 44.3094 $w=2.23e-07 $l=2.69768e-07 $layer=POLY_cond $X=0.27 $Y=1.54
+ $X2=0.475 $Y2=1.39
r79 1 2 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.54 $X2=0.27
+ $Y2=2.6
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TBUFI_1%A_27_115# 1 3 11 16 20 24 28 30 33
r50 29 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.22
+ $X2=0.26 $Y2=2.22
r51 28 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.22
+ $X2=0.8 $Y2=2.22
r52 28 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=2.22
+ $X2=0.345 $Y2=2.22
r53 24 26 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.205
+ $X2=0.26 $Y2=4.565
r54 22 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.305
+ $X2=0.26 $Y2=2.22
r55 22 24 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=0.26 $Y=2.305 $X2=0.26
+ $Y2=3.205
r56 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.135
+ $X2=0.26 $Y2=2.22
r57 18 20 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=0.26 $Y=2.135
+ $X2=0.26 $Y2=0.865
r58 14 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=2.22 $X2=0.8 $Y2=2.22
r59 14 16 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.8 $Y=2.22
+ $X2=0.905 $Y2=2.22
r60 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.385
+ $X2=0.905 $Y2=2.22
r61 9 11 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=0.905 $Y=2.385
+ $X2=0.905 $Y2=3.825
r62 3 26 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r63 3 24 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.205
r64 1 20 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TBUFI_1%A 3 7 10 15 20 23
c47 10 0 1.90743e-19 $X=1.325 $Y=1.83
c48 3 0 6.95226e-20 $X=1.265 $Y=0.945
r49 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.83
+ $X2=1.325 $Y2=1.83
r50 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=3.07
+ $X2=1.14 $Y2=3.07
r51 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.915
+ $X2=1.14 $Y2=1.83
r52 13 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=1.915
+ $X2=1.14 $Y2=3.07
r53 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.83 $X2=1.325 $Y2=1.83
r54 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.83
+ $X2=1.325 $Y2=1.995
r55 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.83
+ $X2=1.325 $Y2=1.665
r56 7 12 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=1.265 $Y=3.825
+ $X2=1.265 $Y2=1.995
r57 3 11 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.265 $Y=0.945
+ $X2=1.265 $Y2=1.665
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__TBUFI_1%Y 1 3 10 16 26 29 32
r35 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=2.215
+ $X2=1.48 $Y2=2.33
r36 24 26 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=2.215
+ $X2=1.48 $Y2=1.56
r37 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.335
+ $X2=1.48 $Y2=1.22
r38 23 26 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.335
+ $X2=1.48 $Y2=1.56
r39 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.48 $Y=3.205
+ $X2=1.48 $Y2=4.565
r40 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.33
+ $X2=1.48 $Y2=2.33
r41 16 19 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.48 $Y=2.33
+ $X2=1.48 $Y2=3.205
r42 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1.22
+ $X2=1.48 $Y2=1.22
r43 10 13 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.48 $Y=0.865
+ $X2=1.48 $Y2=1.22
r44 3 21 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.48 $Y2=4.565
r45 3 19 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=2.825 $X2=1.48 $Y2=3.205
r46 1 10 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.48 $Y2=0.865
.ends

