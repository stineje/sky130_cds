* File: sky130_osu_sc_12T_ms__buf_4.pxi.spice
* Created: Fri Nov 12 15:21:45 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__BUF_4%GND N_GND_M1003_d N_GND_M1001_s N_GND_M1009_s
+ N_GND_M1003_b N_GND_c_2_p N_GND_c_12_p N_GND_c_21_p N_GND_c_3_p N_GND_c_27_p
+ GND N_GND_c_22_p PM_SKY130_OSU_SC_12T_MS__BUF_4%GND
x_PM_SKY130_OSU_SC_12T_MS__BUF_4%VDD N_VDD_M1002_d N_VDD_M1005_s N_VDD_M1007_s
+ N_VDD_M1002_b N_VDD_c_63_p N_VDD_c_64_p N_VDD_c_73_p N_VDD_c_78_p N_VDD_c_85_p
+ N_VDD_c_90_p VDD N_VDD_c_65_p PM_SKY130_OSU_SC_12T_MS__BUF_4%VDD
x_PM_SKY130_OSU_SC_12T_MS__BUF_4%A N_A_M1003_g N_A_M1002_g N_A_c_110_n
+ N_A_c_111_n A PM_SKY130_OSU_SC_12T_MS__BUF_4%A
x_PM_SKY130_OSU_SC_12T_MS__BUF_4%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1002_s N_A_27_115#_M1000_g N_A_27_115#_c_177_n
+ N_A_27_115#_M1004_g N_A_27_115#_c_148_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_181_n N_A_27_115#_M1005_g N_A_27_115#_c_152_n
+ N_A_27_115#_c_154_n N_A_27_115#_c_155_n N_A_27_115#_c_156_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_189_n N_A_27_115#_M1006_g
+ N_A_27_115#_c_161_n N_A_27_115#_c_162_n N_A_27_115#_M1009_g
+ N_A_27_115#_c_194_n N_A_27_115#_M1007_g N_A_27_115#_c_167_n
+ N_A_27_115#_c_168_n N_A_27_115#_c_169_n N_A_27_115#_c_172_n
+ N_A_27_115#_c_173_n N_A_27_115#_c_175_n N_A_27_115#_c_176_n
+ PM_SKY130_OSU_SC_12T_MS__BUF_4%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__BUF_4%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1004_d
+ N_Y_M1006_d N_Y_c_263_n N_Y_c_286_n N_Y_c_267_n N_Y_c_289_n N_Y_c_271_n
+ N_Y_c_275_n Y N_Y_c_277_n N_Y_c_293_n N_Y_c_281_n N_Y_c_285_n
+ PM_SKY130_OSU_SC_12T_MS__BUF_4%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.0588895f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1003_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_A_M1003_g 0.00607478f $X=1.635 $Y=0.152 $X2=0.475 $Y2=0.835
cc_4 N_GND_M1003_b N_A_M1002_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_5 N_GND_M1003_b N_A_c_110_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_6 N_GND_M1003_b N_A_c_111_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_7 N_GND_M1003_b N_A_27_115#_M1000_g 0.0207482f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.835
cc_8 N_GND_c_2_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.905
+ $Y2=0.835
cc_9 N_GND_c_3_p N_A_27_115#_M1000_g 0.00607478f $X=1.635 $Y=0.152 $X2=0.905
+ $Y2=0.835
cc_10 N_GND_M1003_b N_A_27_115#_c_148_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.38
cc_11 N_GND_M1003_b N_A_27_115#_M1001_g 0.0202101f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.835
cc_12 N_GND_c_12_p N_A_27_115#_M1001_g 0.00311745f $X=1.55 $Y=0.755 $X2=1.335
+ $Y2=0.835
cc_13 N_GND_c_3_p N_A_27_115#_M1001_g 0.00607478f $X=1.635 $Y=0.152 $X2=1.335
+ $Y2=0.835
cc_14 N_GND_M1003_b N_A_27_115#_c_152_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.365
cc_15 N_GND_c_12_p N_A_27_115#_c_152_n 0.00256938f $X=1.55 $Y=0.755 $X2=1.69
+ $Y2=1.365
cc_16 N_GND_M1003_b N_A_27_115#_c_154_n 0.0479019f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.365
cc_17 N_GND_M1003_b N_A_27_115#_c_155_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.455
cc_18 N_GND_M1003_b N_A_27_115#_c_156_n 0.0244408f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.455
cc_19 N_GND_M1003_b N_A_27_115#_M1008_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.835
cc_20 N_GND_c_12_p N_A_27_115#_M1008_g 0.00311745f $X=1.55 $Y=0.755 $X2=1.765
+ $Y2=0.835
cc_21 N_GND_c_21_p N_A_27_115#_M1008_g 0.00606474f $X=2.325 $Y=0.152 $X2=1.765
+ $Y2=0.835
cc_22 N_GND_c_22_p N_A_27_115#_M1008_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.765
+ $Y2=0.835
cc_23 N_GND_M1003_b N_A_27_115#_c_161_n 0.0385034f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.365
cc_24 N_GND_M1003_b N_A_27_115#_c_162_n 0.0221499f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.455
cc_25 N_GND_M1003_b N_A_27_115#_M1009_g 0.0264941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.835
cc_26 N_GND_c_21_p N_A_27_115#_M1009_g 0.00606474f $X=2.325 $Y=0.152 $X2=2.195
+ $Y2=0.835
cc_27 N_GND_c_27_p N_A_27_115#_M1009_g 0.00502587f $X=2.41 $Y=0.755 $X2=2.195
+ $Y2=0.835
cc_28 N_GND_c_22_p N_A_27_115#_M1009_g 0.00468827f $X=1.7 $Y=0.19 $X2=2.195
+ $Y2=0.835
cc_29 N_GND_M1003_b N_A_27_115#_c_167_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.365
cc_30 N_GND_M1003_b N_A_27_115#_c_168_n 0.00890086f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.455
cc_31 N_GND_M1003_b N_A_27_115#_c_169_n 0.0142137f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_32 N_GND_c_3_p N_A_27_115#_c_169_n 0.00895373f $X=1.635 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_33 N_GND_c_22_p N_A_27_115#_c_169_n 0.00136847f $X=1.7 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_34 N_GND_M1003_b N_A_27_115#_c_172_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.955
cc_35 N_GND_M1003_b N_A_27_115#_c_173_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.455
cc_36 N_GND_c_2_p N_A_27_115#_c_173_n 0.00702738f $X=0.69 $Y=0.755 $X2=0.88
+ $Y2=1.455
cc_37 N_GND_M1003_b N_A_27_115#_c_175_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.455
cc_38 N_GND_M1003_b N_A_27_115#_c_176_n 0.00592383f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.455
cc_39 N_GND_M1003_b N_Y_c_263_n 0.00153033f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.755
cc_40 N_GND_c_12_p N_Y_c_263_n 8.14297e-19 $X=1.55 $Y=0.755 $X2=1.12 $Y2=0.755
cc_41 N_GND_c_3_p N_Y_c_263_n 0.00800299f $X=1.635 $Y=0.152 $X2=1.12 $Y2=0.755
cc_42 N_GND_c_22_p N_Y_c_263_n 0.00132073f $X=1.7 $Y=0.19 $X2=1.12 $Y2=0.755
cc_43 N_GND_M1003_b N_Y_c_267_n 0.00154299f $X=-0.045 $Y=0 $X2=1.98 $Y2=0.755
cc_44 N_GND_c_12_p N_Y_c_267_n 8.14297e-19 $X=1.55 $Y=0.755 $X2=1.98 $Y2=0.755
cc_45 N_GND_c_21_p N_Y_c_267_n 0.00738926f $X=2.325 $Y=0.152 $X2=1.98 $Y2=0.755
cc_46 N_GND_c_22_p N_Y_c_267_n 0.0047139f $X=1.7 $Y=0.19 $X2=1.98 $Y2=0.755
cc_47 N_GND_M1003_b N_Y_c_271_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.115
cc_48 N_GND_c_2_p N_Y_c_271_n 0.00134236f $X=0.69 $Y=0.755 $X2=1.12 $Y2=1.115
cc_49 N_GND_c_12_p N_Y_c_271_n 7.53951e-19 $X=1.55 $Y=0.755 $X2=1.12 $Y2=1.115
cc_50 N_GND_c_3_p N_Y_c_271_n 0.00282311f $X=1.635 $Y=0.152 $X2=1.12 $Y2=1.115
cc_51 N_GND_M1003_b N_Y_c_275_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.365
cc_52 N_GND_M1003_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=1.79
cc_53 N_GND_M1001_s N_Y_c_277_n 0.0100321f $X=1.41 $Y=0.575 $X2=1.835 $Y2=1
cc_54 N_GND_c_12_p N_Y_c_277_n 0.0142303f $X=1.55 $Y=0.755 $X2=1.835 $Y2=1
cc_55 N_GND_c_21_p N_Y_c_277_n 0.0028844f $X=2.325 $Y=0.152 $X2=1.835 $Y2=1
cc_56 N_GND_c_3_p N_Y_c_277_n 0.00288904f $X=1.635 $Y=0.152 $X2=1.835 $Y2=1
cc_57 N_GND_M1003_b N_Y_c_281_n 0.00409378f $X=-0.045 $Y=0 $X2=1.98 $Y2=1.115
cc_58 N_GND_c_12_p N_Y_c_281_n 7.53951e-19 $X=1.55 $Y=0.755 $X2=1.98 $Y2=1.115
cc_59 N_GND_c_21_p N_Y_c_281_n 0.00245319f $X=2.325 $Y=0.152 $X2=1.98 $Y2=1.115
cc_60 N_GND_c_27_p N_Y_c_281_n 0.00134236f $X=2.41 $Y=0.755 $X2=1.98 $Y2=1.115
cc_61 N_GND_M1003_b N_Y_c_285_n 0.0651512f $X=-0.045 $Y=0 $X2=1.98 $Y2=2.365
cc_62 N_VDD_M1002_b N_A_M1002_g 0.0245629f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_63 N_VDD_c_63_p N_A_M1002_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=3.235
cc_64 N_VDD_c_64_p N_A_M1002_g 0.00337744f $X=0.69 $Y=3.635 $X2=0.475 $Y2=3.235
cc_65 N_VDD_c_65_p N_A_M1002_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.475 $Y2=3.235
cc_66 N_VDD_M1002_d N_A_c_111_n 0.00628533f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2
cc_67 N_VDD_M1002_b N_A_c_111_n 0.00328912f $X=-0.045 $Y=2.425 $X2=0.635 $Y2=2
cc_68 N_VDD_c_64_p N_A_c_111_n 0.00264661f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2
cc_69 N_VDD_M1002_d A 0.00797576f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2.85
cc_70 N_VDD_c_64_p A 0.00510982f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2.85
cc_71 N_VDD_M1002_b N_A_27_115#_c_177_n 0.014249f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.53
cc_72 N_VDD_c_64_p N_A_27_115#_c_177_n 0.00337744f $X=0.69 $Y=3.635 $X2=0.905
+ $Y2=2.53
cc_73 N_VDD_c_73_p N_A_27_115#_c_177_n 0.00606474f $X=1.465 $Y=4.287 $X2=0.905
+ $Y2=2.53
cc_74 N_VDD_c_65_p N_A_27_115#_c_177_n 0.00468827f $X=1.7 $Y=4.25 $X2=0.905
+ $Y2=2.53
cc_75 N_VDD_M1002_b N_A_27_115#_c_181_n 0.0141063f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.53
cc_76 N_VDD_c_64_p N_A_27_115#_c_181_n 3.67508e-19 $X=0.69 $Y=3.635 $X2=1.335
+ $Y2=2.53
cc_77 N_VDD_c_73_p N_A_27_115#_c_181_n 0.00610567f $X=1.465 $Y=4.287 $X2=1.335
+ $Y2=2.53
cc_78 N_VDD_c_78_p N_A_27_115#_c_181_n 0.0035715f $X=1.55 $Y=2.955 $X2=1.335
+ $Y2=2.53
cc_79 N_VDD_c_65_p N_A_27_115#_c_181_n 0.00470215f $X=1.7 $Y=4.25 $X2=1.335
+ $Y2=2.53
cc_80 N_VDD_M1002_b N_A_27_115#_c_155_n 0.00647677f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.455
cc_81 N_VDD_c_78_p N_A_27_115#_c_155_n 0.00364479f $X=1.55 $Y=2.955 $X2=1.69
+ $Y2=2.455
cc_82 N_VDD_M1002_b N_A_27_115#_c_156_n 0.0113915f $X=-0.045 $Y=2.425 $X2=1.41
+ $Y2=2.455
cc_83 N_VDD_M1002_b N_A_27_115#_c_189_n 0.0137901f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.53
cc_84 N_VDD_c_78_p N_A_27_115#_c_189_n 0.00337744f $X=1.55 $Y=2.955 $X2=1.765
+ $Y2=2.53
cc_85 N_VDD_c_85_p N_A_27_115#_c_189_n 0.00606474f $X=2.325 $Y=4.287 $X2=1.765
+ $Y2=2.53
cc_86 N_VDD_c_65_p N_A_27_115#_c_189_n 0.00468827f $X=1.7 $Y=4.25 $X2=1.765
+ $Y2=2.53
cc_87 N_VDD_M1002_b N_A_27_115#_c_162_n 0.0134369f $X=-0.045 $Y=2.425 $X2=2.12
+ $Y2=2.455
cc_88 N_VDD_M1002_b N_A_27_115#_c_194_n 0.0166569f $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.53
cc_89 N_VDD_c_85_p N_A_27_115#_c_194_n 0.00606474f $X=2.325 $Y=4.287 $X2=2.195
+ $Y2=2.53
cc_90 N_VDD_c_90_p N_A_27_115#_c_194_n 0.00636672f $X=2.41 $Y=2.955 $X2=2.195
+ $Y2=2.53
cc_91 N_VDD_c_65_p N_A_27_115#_c_194_n 0.00468827f $X=1.7 $Y=4.25 $X2=2.195
+ $Y2=2.53
cc_92 N_VDD_M1002_b N_A_27_115#_c_168_n 0.00167153f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.455
cc_93 N_VDD_M1002_b N_A_27_115#_c_172_n 0.00996008f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=2.955
cc_94 N_VDD_c_63_p N_A_27_115#_c_172_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=2.955
cc_95 N_VDD_c_65_p N_A_27_115#_c_172_n 0.00476261f $X=1.7 $Y=4.25 $X2=0.26
+ $Y2=2.955
cc_96 N_VDD_M1002_b N_Y_c_286_n 0.00290209f $X=-0.045 $Y=2.425 $X2=1.12 $Y2=2.48
cc_97 N_VDD_c_73_p N_Y_c_286_n 0.00734006f $X=1.465 $Y=4.287 $X2=1.12 $Y2=2.48
cc_98 N_VDD_c_65_p N_Y_c_286_n 0.00475776f $X=1.7 $Y=4.25 $X2=1.12 $Y2=2.48
cc_99 N_VDD_M1002_b N_Y_c_289_n 0.00337919f $X=-0.045 $Y=2.425 $X2=1.98 $Y2=2.48
cc_100 N_VDD_c_85_p N_Y_c_289_n 0.00754406f $X=2.325 $Y=4.287 $X2=1.98 $Y2=2.48
cc_101 N_VDD_c_65_p N_Y_c_289_n 0.00475776f $X=1.7 $Y=4.25 $X2=1.98 $Y2=2.48
cc_102 N_VDD_M1002_b N_Y_c_275_n 0.00409378f $X=-0.045 $Y=2.425 $X2=1.12
+ $Y2=2.365
cc_103 N_VDD_M1002_b N_Y_c_293_n 0.00520877f $X=-0.045 $Y=2.425 $X2=1.835
+ $Y2=2.48
cc_104 N_VDD_c_78_p N_Y_c_293_n 0.0090257f $X=1.55 $Y=2.955 $X2=1.835 $Y2=2.48
cc_105 N_VDD_M1002_b N_Y_c_285_n 0.00409378f $X=-0.045 $Y=2.425 $X2=1.98
+ $Y2=2.365
cc_106 A N_A_27_115#_M1002_s 0.00410657f $X=0.635 $Y=2.85 $X2=0.135 $Y2=2.605
cc_107 N_A_M1003_g N_A_27_115#_M1000_g 0.0342527f $X=0.475 $Y=0.835 $X2=0.905
+ $Y2=0.835
cc_108 A N_A_27_115#_c_177_n 0.00419145f $X=0.635 $Y=2.85 $X2=0.905 $Y2=2.53
cc_109 N_A_M1003_g N_A_27_115#_c_148_n 0.00260138f $X=0.475 $Y=0.835 $X2=1.18
+ $Y2=2.38
cc_110 N_A_M1002_g N_A_27_115#_c_148_n 0.00209773f $X=0.475 $Y=3.235 $X2=1.18
+ $Y2=2.38
cc_111 N_A_c_110_n N_A_27_115#_c_148_n 0.0139096f $X=0.635 $Y=2 $X2=1.18
+ $Y2=2.38
cc_112 N_A_c_111_n N_A_27_115#_c_148_n 0.00361737f $X=0.635 $Y=2 $X2=1.18
+ $Y2=2.38
cc_113 N_A_M1002_g N_A_27_115#_c_156_n 0.0485392f $X=0.475 $Y=3.235 $X2=1.41
+ $Y2=2.455
cc_114 N_A_c_111_n N_A_27_115#_c_156_n 0.00477416f $X=0.635 $Y=2 $X2=1.41
+ $Y2=2.455
cc_115 N_A_M1003_g N_A_27_115#_c_169_n 0.0124465f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.755
cc_116 N_A_M1003_g N_A_27_115#_c_172_n 0.0330322f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=2.955
cc_117 N_A_c_111_n N_A_27_115#_c_172_n 0.0548951f $X=0.635 $Y=2 $X2=0.26
+ $Y2=2.955
cc_118 A N_A_27_115#_c_172_n 0.0155137f $X=0.635 $Y=2.85 $X2=0.26 $Y2=2.955
cc_119 N_A_M1003_g N_A_27_115#_c_173_n 0.0207696f $X=0.475 $Y=0.835 $X2=0.88
+ $Y2=1.455
cc_120 N_A_c_110_n N_A_27_115#_c_173_n 0.00273049f $X=0.635 $Y=2 $X2=0.88
+ $Y2=1.455
cc_121 N_A_c_111_n N_A_27_115#_c_173_n 0.00886797f $X=0.635 $Y=2 $X2=0.88
+ $Y2=1.455
cc_122 N_A_M1003_g N_A_27_115#_c_176_n 6.59135e-19 $X=0.475 $Y=0.835 $X2=0.965
+ $Y2=1.455
cc_123 N_A_c_111_n N_Y_c_286_n 0.0135622f $X=0.635 $Y=2 $X2=1.12 $Y2=2.48
cc_124 A N_Y_c_286_n 0.00731851f $X=0.635 $Y=2.85 $X2=1.12 $Y2=2.48
cc_125 N_A_M1003_g N_Y_c_271_n 8.01483e-19 $X=0.475 $Y=0.835 $X2=1.12 $Y2=1.115
cc_126 N_A_c_111_n N_Y_c_275_n 0.00677552f $X=0.635 $Y=2 $X2=1.12 $Y2=2.365
cc_127 N_A_M1003_g Y 0.00310306f $X=0.475 $Y=0.835 $X2=1.055 $Y2=1.79
cc_128 N_A_c_110_n Y 0.00441844f $X=0.635 $Y=2 $X2=1.055 $Y2=1.79
cc_129 N_A_c_111_n Y 0.0200396f $X=0.635 $Y=2 $X2=1.055 $Y2=1.79
cc_130 N_A_27_115#_M1000_g N_Y_c_263_n 0.00182852f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_131 N_A_27_115#_M1001_g N_Y_c_263_n 0.00182852f $X=1.335 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_132 N_A_27_115#_c_154_n N_Y_c_263_n 0.00296072f $X=1.41 $Y=1.365 $X2=1.12
+ $Y2=0.755
cc_133 N_A_27_115#_c_176_n N_Y_c_263_n 7.29965e-19 $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=0.755
cc_134 N_A_27_115#_c_177_n N_Y_c_286_n 0.00138273f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_135 N_A_27_115#_c_181_n N_Y_c_286_n 0.00233646f $X=1.335 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_136 N_A_27_115#_c_156_n N_Y_c_286_n 0.0126676f $X=1.41 $Y=2.455 $X2=1.12
+ $Y2=2.48
cc_137 N_A_27_115#_M1008_g N_Y_c_267_n 0.00182852f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=0.755
cc_138 N_A_27_115#_c_161_n N_Y_c_267_n 0.00274041f $X=2.12 $Y=1.365 $X2=1.98
+ $Y2=0.755
cc_139 N_A_27_115#_M1009_g N_Y_c_267_n 0.00182852f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=0.755
cc_140 N_A_27_115#_c_189_n N_Y_c_289_n 0.00233646f $X=1.765 $Y=2.53 $X2=1.98
+ $Y2=2.48
cc_141 N_A_27_115#_c_162_n N_Y_c_289_n 0.013404f $X=2.12 $Y=2.455 $X2=1.98
+ $Y2=2.48
cc_142 N_A_27_115#_c_194_n N_Y_c_289_n 0.00233646f $X=2.195 $Y=2.53 $X2=1.98
+ $Y2=2.48
cc_143 N_A_27_115#_M1000_g N_Y_c_271_n 0.00480694f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=1.115
cc_144 N_A_27_115#_M1001_g N_Y_c_271_n 0.00198614f $X=1.335 $Y=0.835 $X2=1.12
+ $Y2=1.115
cc_145 N_A_27_115#_c_176_n N_Y_c_271_n 0.00278861f $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=1.115
cc_146 N_A_27_115#_c_177_n N_Y_c_275_n 0.00120715f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.365
cc_147 N_A_27_115#_c_148_n N_Y_c_275_n 0.00215118f $X=1.18 $Y=2.38 $X2=1.12
+ $Y2=2.365
cc_148 N_A_27_115#_c_181_n N_Y_c_275_n 0.00113627f $X=1.335 $Y=2.53 $X2=1.12
+ $Y2=2.365
cc_149 N_A_27_115#_c_156_n N_Y_c_275_n 0.0038035f $X=1.41 $Y=2.455 $X2=1.12
+ $Y2=2.365
cc_150 N_A_27_115#_M1000_g Y 0.00251111f $X=0.905 $Y=0.835 $X2=1.055 $Y2=1.79
cc_151 N_A_27_115#_c_148_n Y 0.0314621f $X=1.18 $Y=2.38 $X2=1.055 $Y2=1.79
cc_152 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=0.835 $X2=1.055 $Y2=1.79
cc_153 N_A_27_115#_c_154_n Y 0.0166018f $X=1.41 $Y=1.365 $X2=1.055 $Y2=1.79
cc_154 N_A_27_115#_c_173_n Y 8.73078e-19 $X=0.88 $Y=1.455 $X2=1.055 $Y2=1.79
cc_155 N_A_27_115#_c_176_n Y 0.0121742f $X=0.965 $Y=1.455 $X2=1.055 $Y2=1.79
cc_156 N_A_27_115#_M1001_g N_Y_c_277_n 0.00872983f $X=1.335 $Y=0.835 $X2=1.835
+ $Y2=1
cc_157 N_A_27_115#_c_152_n N_Y_c_277_n 0.00213861f $X=1.69 $Y=1.365 $X2=1.835
+ $Y2=1
cc_158 N_A_27_115#_M1008_g N_Y_c_277_n 0.00873177f $X=1.765 $Y=0.835 $X2=1.835
+ $Y2=1
cc_159 N_A_27_115#_c_181_n N_Y_c_293_n 0.00639369f $X=1.335 $Y=2.53 $X2=1.835
+ $Y2=2.48
cc_160 N_A_27_115#_c_155_n N_Y_c_293_n 0.0125005f $X=1.69 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_161 N_A_27_115#_c_156_n N_Y_c_293_n 0.00580646f $X=1.41 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_162 N_A_27_115#_c_189_n N_Y_c_293_n 0.00639369f $X=1.765 $Y=2.53 $X2=1.835
+ $Y2=2.48
cc_163 N_A_27_115#_c_168_n N_Y_c_293_n 0.00580646f $X=1.765 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_164 N_A_27_115#_M1008_g N_Y_c_281_n 0.00198614f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=1.115
cc_165 N_A_27_115#_M1009_g N_Y_c_281_n 0.00878256f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=1.115
cc_166 N_A_27_115#_c_154_n N_Y_c_285_n 0.013329f $X=1.41 $Y=1.365 $X2=1.98
+ $Y2=2.365
cc_167 N_A_27_115#_M1008_g N_Y_c_285_n 0.00251111f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=2.365
cc_168 N_A_27_115#_c_189_n N_Y_c_285_n 0.00113627f $X=1.765 $Y=2.53 $X2=1.98
+ $Y2=2.365
cc_169 N_A_27_115#_c_161_n N_Y_c_285_n 0.0170354f $X=2.12 $Y=1.365 $X2=1.98
+ $Y2=2.365
cc_170 N_A_27_115#_c_162_n N_Y_c_285_n 0.00966211f $X=2.12 $Y=2.455 $X2=1.98
+ $Y2=2.365
cc_171 N_A_27_115#_M1009_g N_Y_c_285_n 0.00251111f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=2.365
cc_172 N_A_27_115#_c_194_n N_Y_c_285_n 0.0031083f $X=2.195 $Y=2.53 $X2=1.98
+ $Y2=2.365
cc_173 N_A_27_115#_c_168_n N_Y_c_285_n 6.99501e-19 $X=1.765 $Y=2.455 $X2=1.98
+ $Y2=2.365
