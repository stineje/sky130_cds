* File: sky130_osu_sc_12T_hs__aoi22_l.pxi.spice
* Created: Fri Nov 12 15:07:55 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%GND N_GND_M1004_s N_GND_M1007_d N_GND_M1004_b
+ N_GND_c_3_p N_GND_c_4_p N_GND_c_28_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_12T_HS__AOI22_L%GND
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%VDD N_VDD_M1000_d N_VDD_M1000_b N_VDD_c_48_p
+ N_VDD_c_49_p N_VDD_c_54_p VDD N_VDD_c_50_p
+ PM_SKY130_OSU_SC_12T_HS__AOI22_L%VDD
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%A0 N_A0_c_76_n N_A0_c_77_n N_A0_M1004_g
+ N_A0_M1000_g N_A0_c_81_n N_A0_c_83_n N_A0_c_84_n A0
+ PM_SKY130_OSU_SC_12T_HS__AOI22_L%A0
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%A1 N_A1_M1002_g N_A1_c_112_n N_A1_M1005_g
+ N_A1_c_114_n A1 PM_SKY130_OSU_SC_12T_HS__AOI22_L%A1
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%B0 N_B0_M1001_g N_B0_M1006_g N_B0_c_157_n
+ N_B0_c_158_n N_B0_c_159_n B0 PM_SKY130_OSU_SC_12T_HS__AOI22_L%B0
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%B1 N_B1_M1007_g N_B1_M1003_g N_B1_c_200_n
+ N_B1_c_202_n B1 PM_SKY130_OSU_SC_12T_HS__AOI22_L%B1
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%A_27_521# N_A_27_521#_M1000_s
+ N_A_27_521#_M1005_d N_A_27_521#_M1003_d N_A_27_521#_c_221_n
+ N_A_27_521#_c_223_n N_A_27_521#_c_234_n N_A_27_521#_c_225_n
+ N_A_27_521#_c_228_n PM_SKY130_OSU_SC_12T_HS__AOI22_L%A_27_521#
x_PM_SKY130_OSU_SC_12T_HS__AOI22_L%Y N_Y_M1002_d N_Y_M1006_d N_Y_c_244_n
+ N_Y_c_282_n N_Y_c_247_n N_Y_c_248_n N_Y_c_250_n Y N_Y_c_254_n
+ PM_SKY130_OSU_SC_12T_HS__AOI22_L%Y
cc_1 N_GND_M1004_b N_A0_c_76_n 0.0639487f $X=-0.045 $Y=0 $X2=0.295 $Y2=2.15
cc_2 N_GND_M1004_b N_A0_c_77_n 0.0174934f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.21
cc_3 N_GND_c_3_p N_A0_c_77_n 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=1.21
cc_4 N_GND_c_4_p N_A0_c_77_n 0.00606474f $X=1.825 $Y=0.152 $X2=0.475 $Y2=1.21
cc_5 N_GND_c_5_p N_A0_c_77_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=1.21
cc_6 N_GND_M1004_b N_A0_c_81_n 0.0299632f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.29
cc_7 N_GND_c_3_p N_A0_c_81_n 0.00534003f $X=0.26 $Y=0.755 $X2=0.475 $Y2=1.29
cc_8 N_GND_M1004_b N_A0_c_83_n 0.0395437f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.285
cc_9 N_GND_M1004_b N_A0_c_84_n 0.0018756f $X=-0.045 $Y=0 $X2=0.385 $Y2=2.11
cc_10 N_GND_M1004_b A0 0.00797389f $X=-0.045 $Y=0 $X2=0.385 $Y2=2.11
cc_11 N_GND_M1004_b N_A1_M1002_g 0.036803f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.85
cc_12 N_GND_c_4_p N_A1_M1002_g 0.00606474f $X=1.825 $Y=0.152 $X2=0.835 $Y2=0.85
cc_13 N_GND_c_5_p N_A1_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.835 $Y2=0.85
cc_14 N_GND_M1004_b N_A1_c_112_n 0.0514426f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.09
cc_15 N_GND_M1004_b N_A1_M1005_g 0.01783f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_16 N_GND_M1004_b N_A1_c_114_n 0.011098f $X=-0.045 $Y=0 $X2=0.725 $Y2=1.775
cc_17 N_GND_M1004_b A1 0.00153071f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.48
cc_18 N_GND_M1004_b N_B0_M1001_g 0.0178475f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.85
cc_19 N_GND_c_4_p N_B0_M1001_g 0.00606474f $X=1.825 $Y=0.152 $X2=1.335 $Y2=0.85
cc_20 N_GND_c_5_p N_B0_M1001_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335 $Y2=0.85
cc_21 N_GND_M1004_b N_B0_M1006_g 0.0435719f $X=-0.045 $Y=0 $X2=1.335 $Y2=3.235
cc_22 N_GND_M1004_b N_B0_c_157_n 0.0272094f $X=-0.045 $Y=0 $X2=1.255 $Y2=1.42
cc_23 N_GND_M1004_b N_B0_c_158_n 0.0123234f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.11
cc_24 N_GND_M1004_b N_B0_c_159_n 0.00417976f $X=-0.045 $Y=0 $X2=1.165 $Y2=1.42
cc_25 N_GND_M1004_b B0 0.0143696f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.11
cc_26 N_GND_M1004_b N_B1_M1007_g 0.0412241f $X=-0.045 $Y=0 $X2=1.695 $Y2=0.85
cc_27 N_GND_c_4_p N_B1_M1007_g 0.00606474f $X=1.825 $Y=0.152 $X2=1.695 $Y2=0.85
cc_28 N_GND_c_28_p N_B1_M1007_g 0.00502587f $X=1.91 $Y=0.755 $X2=1.695 $Y2=0.85
cc_29 N_GND_c_5_p N_B1_M1007_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.695 $Y2=0.85
cc_30 N_GND_M1004_b N_B1_M1003_g 0.0424628f $X=-0.045 $Y=0 $X2=1.765 $Y2=3.235
cc_31 N_GND_M1004_b N_B1_c_200_n 0.0574006f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.722
cc_32 N_GND_c_28_p N_B1_c_200_n 0.00159696f $X=1.91 $Y=0.755 $X2=1.765 $Y2=1.722
cc_33 N_GND_M1004_b N_B1_c_202_n 0.00957801f $X=-0.045 $Y=0 $X2=1.935 $Y2=1.74
cc_34 N_GND_c_28_p N_B1_c_202_n 0.00415495f $X=1.91 $Y=0.755 $X2=1.935 $Y2=1.74
cc_35 N_GND_M1004_b B1 0.0102463f $X=-0.045 $Y=0 $X2=1.935 $Y2=1.74
cc_36 N_GND_M1004_b N_Y_c_244_n 0.00156158f $X=-0.045 $Y=0 $X2=1.085 $Y2=0.755
cc_37 N_GND_c_4_p N_Y_c_244_n 0.00722805f $X=1.825 $Y=0.152 $X2=1.085 $Y2=0.755
cc_38 N_GND_c_5_p N_Y_c_244_n 0.00472308f $X=1.7 $Y=0.19 $X2=1.085 $Y2=0.755
cc_39 N_GND_M1004_b N_Y_c_247_n 0.0173617f $X=-0.045 $Y=0 $X2=1.595 $Y2=1.37
cc_40 N_GND_c_4_p N_Y_c_248_n 0.00774628f $X=1.825 $Y=0.152 $X2=1.52 $Y2=1
cc_41 N_GND_c_28_p N_Y_c_248_n 7.45493e-19 $X=1.91 $Y=0.755 $X2=1.52 $Y2=1
cc_42 N_GND_c_3_p N_Y_c_250_n 0.00115996f $X=0.26 $Y=0.755 $X2=1.23 $Y2=1
cc_43 N_GND_c_4_p N_Y_c_250_n 0.00263877f $X=1.825 $Y=0.152 $X2=1.23 $Y2=1
cc_44 N_GND_c_28_p N_Y_c_250_n 6.58722e-19 $X=1.91 $Y=0.755 $X2=1.23 $Y2=1
cc_45 N_GND_M1004_b Y 0.00182066f $X=-0.045 $Y=0 $X2=1.605 $Y2=1.22
cc_46 N_GND_M1004_b N_Y_c_254_n 0.00421975f $X=-0.045 $Y=0 $X2=1.595 $Y2=1.37
cc_47 N_VDD_M1000_b N_A0_M1000_g 0.0287852f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_48 N_VDD_c_48_p N_A0_M1000_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_49 N_VDD_c_49_p N_A0_M1000_g 0.00339848f $X=0.69 $Y=3.655 $X2=0.475 $Y2=3.235
cc_50 N_VDD_c_50_p N_A0_M1000_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.475 $Y2=3.235
cc_51 N_VDD_M1000_b N_A0_c_84_n 0.0024763f $X=-0.045 $Y=2.425 $X2=0.385 $Y2=2.11
cc_52 N_VDD_M1000_b N_A1_M1005_g 0.0189661f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_53 N_VDD_c_49_p N_A1_M1005_g 0.00271216f $X=0.69 $Y=3.655 $X2=0.905 $Y2=3.235
cc_54 N_VDD_c_54_p N_A1_M1005_g 0.00606474f $X=1.7 $Y=4.22 $X2=0.905 $Y2=3.235
cc_55 N_VDD_c_50_p N_A1_M1005_g 0.00468827f $X=1.7 $Y=4.25 $X2=0.905 $Y2=3.235
cc_56 N_VDD_M1000_b N_A1_c_114_n 0.00550561f $X=-0.045 $Y=2.425 $X2=0.725
+ $Y2=1.775
cc_57 N_VDD_M1000_b A1 0.00660952f $X=-0.045 $Y=2.425 $X2=0.725 $Y2=2.48
cc_58 N_VDD_M1000_b N_B0_M1006_g 0.0200589f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=3.235
cc_59 N_VDD_c_54_p N_B0_M1006_g 0.00413449f $X=1.7 $Y=4.22 $X2=1.335 $Y2=3.235
cc_60 N_VDD_c_50_p N_B0_M1006_g 0.00468827f $X=1.7 $Y=4.25 $X2=1.335 $Y2=3.235
cc_61 N_VDD_M1000_b N_B1_M1003_g 0.028148f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=3.235
cc_62 N_VDD_c_54_p N_B1_M1003_g 0.00413449f $X=1.7 $Y=4.22 $X2=1.765 $Y2=3.235
cc_63 N_VDD_c_50_p N_B1_M1003_g 0.00468827f $X=1.7 $Y=4.25 $X2=1.765 $Y2=3.235
cc_64 N_VDD_c_48_p N_A_27_521#_c_221_n 0.00485776f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=3.485
cc_65 N_VDD_c_50_p N_A_27_521#_c_221_n 0.00442406f $X=1.7 $Y=4.25 $X2=0.26
+ $Y2=3.485
cc_66 N_VDD_M1000_d N_A_27_521#_c_223_n 0.00460359f $X=0.55 $Y=2.605 $X2=1.035
+ $Y2=3.145
cc_67 N_VDD_c_49_p N_A_27_521#_c_223_n 0.0135055f $X=0.69 $Y=3.655 $X2=1.035
+ $Y2=3.145
cc_68 N_VDD_M1000_b N_A_27_521#_c_225_n 0.00659135f $X=-0.045 $Y=2.425 $X2=1.895
+ $Y2=3.825
cc_69 N_VDD_c_54_p N_A_27_521#_c_225_n 0.0427205f $X=1.7 $Y=4.22 $X2=1.895
+ $Y2=3.825
cc_70 N_VDD_c_50_p N_A_27_521#_c_225_n 0.0240576f $X=1.7 $Y=4.25 $X2=1.895
+ $Y2=3.825
cc_71 N_VDD_M1000_b N_A_27_521#_c_228_n 0.00182934f $X=-0.045 $Y=2.425 $X2=1.205
+ $Y2=3.825
cc_72 N_VDD_c_49_p N_A_27_521#_c_228_n 0.00275564f $X=0.69 $Y=3.655 $X2=1.205
+ $Y2=3.825
cc_73 N_VDD_c_54_p N_A_27_521#_c_228_n 0.00928857f $X=1.7 $Y=4.22 $X2=1.205
+ $Y2=3.825
cc_74 N_VDD_c_50_p N_A_27_521#_c_228_n 0.00493883f $X=1.7 $Y=4.25 $X2=1.205
+ $Y2=3.825
cc_75 N_VDD_M1000_b N_Y_c_247_n 0.00371086f $X=-0.045 $Y=2.425 $X2=1.595
+ $Y2=1.37
cc_76 N_A0_c_76_n N_A1_M1002_g 0.00899556f $X=0.295 $Y=2.15 $X2=0.835 $Y2=0.85
cc_77 N_A0_c_77_n N_A1_M1002_g 0.0575985f $X=0.475 $Y=1.21 $X2=0.835 $Y2=0.85
cc_78 N_A0_c_76_n N_A1_c_112_n 0.0256414f $X=0.295 $Y=2.15 $X2=0.905 $Y2=2.09
cc_79 A0 N_A1_c_112_n 0.00143344f $X=0.385 $Y=2.11 $X2=0.905 $Y2=2.09
cc_80 N_A0_c_76_n N_A1_M1005_g 0.00113657f $X=0.295 $Y=2.15 $X2=0.905 $Y2=3.235
cc_81 N_A0_c_83_n N_A1_M1005_g 0.063953f $X=0.475 $Y=2.285 $X2=0.905 $Y2=3.235
cc_82 N_A0_c_76_n N_A1_c_114_n 0.00388024f $X=0.295 $Y=2.15 $X2=0.725 $Y2=1.775
cc_83 N_A0_c_83_n N_A1_c_114_n 0.00432627f $X=0.475 $Y=2.285 $X2=0.725 $Y2=1.775
cc_84 N_A0_c_84_n N_A1_c_114_n 0.0279492f $X=0.385 $Y=2.11 $X2=0.725 $Y2=1.775
cc_85 A0 N_A1_c_114_n 0.00370699f $X=0.385 $Y=2.11 $X2=0.725 $Y2=1.775
cc_86 N_A0_c_83_n A1 0.00417236f $X=0.475 $Y=2.285 $X2=0.725 $Y2=2.48
cc_87 N_A0_c_84_n A1 0.00265232f $X=0.385 $Y=2.11 $X2=0.725 $Y2=2.48
cc_88 A0 A1 0.00516633f $X=0.385 $Y=2.11 $X2=0.725 $Y2=2.48
cc_89 A0 B0 0.0147019f $X=0.385 $Y=2.11 $X2=1.165 $Y2=2.11
cc_90 N_A0_M1000_g N_A_27_521#_c_223_n 0.0196156f $X=0.475 $Y=3.235 $X2=1.035
+ $Y2=3.145
cc_91 N_A0_c_84_n N_A_27_521#_c_223_n 0.00272894f $X=0.385 $Y=2.11 $X2=1.035
+ $Y2=3.145
cc_92 N_A0_c_83_n N_A_27_521#_c_234_n 0.00264631f $X=0.475 $Y=2.285 $X2=0.345
+ $Y2=3.145
cc_93 N_A0_c_84_n N_A_27_521#_c_234_n 0.00150818f $X=0.385 $Y=2.11 $X2=0.345
+ $Y2=3.145
cc_94 N_A1_M1002_g N_B0_M1001_g 0.0163064f $X=0.835 $Y=0.85 $X2=1.335 $Y2=0.85
cc_95 N_A1_M1002_g N_B0_M1006_g 0.00961043f $X=0.835 $Y=0.85 $X2=1.335 $Y2=3.235
cc_96 N_A1_c_112_n N_B0_M1006_g 0.0716045f $X=0.905 $Y=2.09 $X2=1.335 $Y2=3.235
cc_97 A1 N_B0_M1006_g 0.0011808f $X=0.725 $Y=2.48 $X2=1.335 $Y2=3.235
cc_98 N_A1_M1002_g N_B0_c_157_n 0.0198874f $X=0.835 $Y=0.85 $X2=1.255 $Y2=1.42
cc_99 N_A1_M1002_g N_B0_c_158_n 0.0032219f $X=0.835 $Y=0.85 $X2=1.165 $Y2=2.11
cc_100 N_A1_c_112_n N_B0_c_158_n 0.00187204f $X=0.905 $Y=2.09 $X2=1.165 $Y2=2.11
cc_101 N_A1_c_114_n N_B0_c_158_n 0.0273961f $X=0.725 $Y=1.775 $X2=1.165 $Y2=2.11
cc_102 N_A1_M1002_g N_B0_c_159_n 0.00591675f $X=0.835 $Y=0.85 $X2=1.165 $Y2=1.42
cc_103 N_A1_c_112_n B0 0.00170611f $X=0.905 $Y=2.09 $X2=1.165 $Y2=2.11
cc_104 N_A1_c_114_n B0 0.00301508f $X=0.725 $Y=1.775 $X2=1.165 $Y2=2.11
cc_105 N_A1_M1005_g N_A_27_521#_c_223_n 0.0157671f $X=0.905 $Y=3.235 $X2=1.035
+ $Y2=3.145
cc_106 N_A1_c_114_n N_A_27_521#_c_223_n 0.00326229f $X=0.725 $Y=1.775 $X2=1.035
+ $Y2=3.145
cc_107 A1 N_A_27_521#_c_223_n 0.0109287f $X=0.725 $Y=2.48 $X2=1.035 $Y2=3.145
cc_108 N_A1_M1005_g N_A_27_521#_c_228_n 9.6635e-19 $X=0.905 $Y=3.235 $X2=1.205
+ $Y2=3.825
cc_109 N_A1_M1002_g N_Y_c_244_n 0.00585218f $X=0.835 $Y=0.85 $X2=1.085 $Y2=0.755
cc_110 A1 N_Y_c_247_n 0.00544969f $X=0.725 $Y=2.48 $X2=1.595 $Y2=1.37
cc_111 N_A1_M1002_g N_Y_c_250_n 0.00458957f $X=0.835 $Y=0.85 $X2=1.23 $Y2=1
cc_112 N_B0_M1001_g N_B1_M1007_g 0.0387476f $X=1.335 $Y=0.85 $X2=1.695 $Y2=0.85
cc_113 N_B0_c_159_n N_B1_M1007_g 4.28925e-19 $X=1.165 $Y=1.42 $X2=1.695 $Y2=0.85
cc_114 N_B0_M1006_g N_B1_c_200_n 0.0738942f $X=1.335 $Y=3.235 $X2=1.765
+ $Y2=1.722
cc_115 N_B0_c_157_n N_B1_c_200_n 0.0387476f $X=1.255 $Y=1.42 $X2=1.765 $Y2=1.722
cc_116 N_B0_M1006_g N_A_27_521#_c_225_n 0.0137697f $X=1.335 $Y=3.235 $X2=1.895
+ $Y2=3.825
cc_117 N_B0_M1001_g N_Y_c_244_n 0.00574971f $X=1.335 $Y=0.85 $X2=1.085 $Y2=0.755
cc_118 N_B0_c_157_n N_Y_c_244_n 0.00112933f $X=1.255 $Y=1.42 $X2=1.085 $Y2=0.755
cc_119 N_B0_c_159_n N_Y_c_244_n 0.00419353f $X=1.165 $Y=1.42 $X2=1.085 $Y2=0.755
cc_120 N_B0_c_157_n N_Y_c_247_n 0.0170201f $X=1.255 $Y=1.42 $X2=1.595 $Y2=1.37
cc_121 N_B0_c_158_n N_Y_c_247_n 0.0298961f $X=1.165 $Y=2.11 $X2=1.595 $Y2=1.37
cc_122 N_B0_c_159_n N_Y_c_247_n 0.0201907f $X=1.165 $Y=1.42 $X2=1.595 $Y2=1.37
cc_123 B0 N_Y_c_247_n 0.00795799f $X=1.165 $Y=2.11 $X2=1.595 $Y2=1.37
cc_124 N_B0_M1001_g N_Y_c_248_n 0.00821935f $X=1.335 $Y=0.85 $X2=1.52 $Y2=1
cc_125 N_B0_c_159_n N_Y_c_248_n 0.00477495f $X=1.165 $Y=1.42 $X2=1.52 $Y2=1
cc_126 N_B0_c_157_n N_Y_c_250_n 0.00131678f $X=1.255 $Y=1.42 $X2=1.23 $Y2=1
cc_127 N_B0_c_159_n N_Y_c_250_n 0.00568984f $X=1.165 $Y=1.42 $X2=1.23 $Y2=1
cc_128 N_B0_M1001_g Y 0.0019765f $X=1.335 $Y=0.85 $X2=1.605 $Y2=1.22
cc_129 N_B0_c_157_n N_Y_c_254_n 0.00382225f $X=1.255 $Y=1.42 $X2=1.595 $Y2=1.37
cc_130 N_B0_c_159_n N_Y_c_254_n 0.00751098f $X=1.165 $Y=1.42 $X2=1.595 $Y2=1.37
cc_131 N_B1_M1003_g N_A_27_521#_c_225_n 0.0154131f $X=1.765 $Y=3.235 $X2=1.895
+ $Y2=3.825
cc_132 N_B1_M1007_g N_Y_c_247_n 0.0097422f $X=1.695 $Y=0.85 $X2=1.595 $Y2=1.37
cc_133 N_B1_c_200_n N_Y_c_247_n 0.0264294f $X=1.765 $Y=1.722 $X2=1.595 $Y2=1.37
cc_134 N_B1_c_202_n N_Y_c_247_n 0.0209729f $X=1.935 $Y=1.74 $X2=1.595 $Y2=1.37
cc_135 B1 N_Y_c_247_n 0.00767175f $X=1.935 $Y=1.74 $X2=1.595 $Y2=1.37
cc_136 N_B1_M1007_g N_Y_c_248_n 0.00855008f $X=1.695 $Y=0.85 $X2=1.52 $Y2=1
cc_137 N_B1_M1007_g Y 0.00642782f $X=1.695 $Y=0.85 $X2=1.605 $Y2=1.22
cc_138 N_B1_M1007_g N_Y_c_254_n 0.011371f $X=1.695 $Y=0.85 $X2=1.595 $Y2=1.37
cc_139 B1 N_Y_c_254_n 0.00552429f $X=1.935 $Y=1.74 $X2=1.595 $Y2=1.37
cc_140 N_A_27_521#_c_225_n N_Y_M1006_d 0.00176461f $X=1.895 $Y=3.825 $X2=1.41
+ $Y2=2.605
cc_141 N_A_27_521#_c_225_n N_Y_c_282_n 0.013096f $X=1.895 $Y=3.825 $X2=1.55
+ $Y2=3.315
cc_142 N_Y_c_248_n A_282_115# 0.0049062f $X=1.52 $Y=1 $X2=1.41 $Y2=0.575
cc_143 Y A_282_115# 3.49194e-19 $X=1.605 $Y=1.22 $X2=1.41 $Y2=0.575
