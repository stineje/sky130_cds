* File: sky130_osu_sc_18T_ms__inv_3.pex.spice
* Created: Fri Nov 12 14:04:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%GND 1 2 21 25 27 35 42 44 47
r45 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r46 33 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r47 33 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r48 27 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r49 23 25 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r50 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r51 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r52 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r53 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r54 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r55 2 35 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r56 1 25 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%VDD 1 2 17 21 25 32 40 42 45
r33 42 45 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r34 32 35 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r35 30 40 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r36 30 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r37 28 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r38 26 39 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r39 26 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r40 25 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r41 25 28 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r42 21 24 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r43 19 39 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r44 19 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r45 17 28 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r46 17 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r47 2 35 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r48 2 32 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r49 1 24 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r50 1 21 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 34 36 37 38 41 43 45 48
c96 33 0 1.5442e-19 $X=0.535 $Y=2.305
c97 28 0 1.33323e-19 $X=1.335 $Y=2.96
c98 25 0 1.33323e-19 $X=1.335 $Y=1.7
c99 18 0 1.33323e-19 $X=0.905 $Y=2.96
c100 15 0 1.33323e-19 $X=0.905 $Y=1.7
r101 48 51 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=3.325
+ $X2=0.405 $Y2=3.33
r102 43 45 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.305
+ $X2=0.535 $Y2=2.305
r103 41 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r104 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=2.39
+ $X2=0.405 $Y2=2.305
r105 39 41 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.39
+ $X2=0.32 $Y2=3.33
r106 33 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.305 $X2=0.535 $Y2=2.305
r107 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.47
r108 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.14
r109 28 30 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r110 25 27 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.335 $Y=1.7
+ $X2=1.335 $Y2=1.075
r111 24 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.885
+ $X2=0.905 $Y2=2.885
r112 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=1.335 $Y2=2.96
r113 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=0.98 $Y2=2.885
r114 22 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.775
+ $X2=0.905 $Y2=1.775
r115 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=1.335 $Y2=1.7
r116 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=0.98 $Y2=1.775
r117 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=2.885
r118 18 20 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=4.585
r119 15 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.775
r120 15 17 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.075
r121 14 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.885
+ $X2=0.475 $Y2=2.885
r122 13 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.905 $Y2=2.885
r123 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.55 $Y2=2.885
r124 12 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.775
+ $X2=0.475 $Y2=1.775
r125 11 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.905 $Y2=1.775
r126 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.55 $Y2=1.775
r127 8 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=2.885
r128 8 10 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=4.585
r129 7 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.885
r130 7 35 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.47
r131 4 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=1.775
r132 4 34 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=2.14
r133 1 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.775
r134 1 3 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c74 55 0 1.33323e-19 $X=1.55 $Y=2.845
c75 54 0 1.33323e-19 $X=1.55 $Y=1.595
c76 46 0 1.33323e-19 $X=0.69 $Y=2.845
c77 45 0 1.33323e-19 $X=0.69 $Y=1.595
c78 18 0 1.5442e-19 $X=0.69 $Y=0.825
r79 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.845
+ $X2=1.55 $Y2=2.96
r80 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r81 54 55 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.845
r82 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.96
+ $X2=0.69 $Y2=2.96
r83 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=1.55 $Y2=2.96
r84 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=0.835 $Y2=2.96
r85 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.48
+ $X2=0.69 $Y2=1.48
r86 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=1.55 $Y2=1.48
r87 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=0.835 $Y2=1.48
r88 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.96
r89 46 48 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.2
r90 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.48
r91 45 48 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=2.2
r92 41 43 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r93 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=2.96
r94 38 41 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=3.455
r95 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r96 32 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r97 27 29 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r98 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=2.96
r99 24 27 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=3.455
r100 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.48
r101 18 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.69 $Y=0.825
+ $X2=0.69 $Y2=1.48
r102 6 43 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r103 6 41 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r104 5 29 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r105 5 27 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r106 2 32 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r107 1 18 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

