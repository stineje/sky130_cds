* File: sky130_osu_sc_15T_ms__and2_8.pxi.spice
* Created: Fri Nov 12 14:40:36 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__AND2_8%GND N_GND_M1003_d N_GND_M1008_s N_GND_M1012_s
+ N_GND_M1015_s N_GND_M1017_s N_GND_M1007_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p
+ N_GND_c_22_p N_GND_c_30_p N_GND_c_36_p N_GND_c_43_p N_GND_c_50_p N_GND_c_57_p
+ N_GND_c_63_p GND N_GND_c_3_p PM_SKY130_OSU_SC_15T_MS__AND2_8%GND
x_PM_SKY130_OSU_SC_15T_MS__AND2_8%VDD N_VDD_M1010_s N_VDD_M1005_d N_VDD_M1001_d
+ N_VDD_M1006_d N_VDD_M1013_d N_VDD_M1019_d N_VDD_M1010_b N_VDD_c_138_p
+ N_VDD_c_139_p N_VDD_c_150_p N_VDD_c_157_p N_VDD_c_163_p N_VDD_c_169_p
+ N_VDD_c_174_p N_VDD_c_180_p N_VDD_c_185_p N_VDD_c_191_p N_VDD_c_196_p VDD
+ N_VDD_c_140_p PM_SKY130_OSU_SC_15T_MS__AND2_8%VDD
x_PM_SKY130_OSU_SC_15T_MS__AND2_8%A N_A_M1007_g N_A_M1010_g N_A_c_227_n
+ N_A_c_228_n A PM_SKY130_OSU_SC_15T_MS__AND2_8%A
x_PM_SKY130_OSU_SC_15T_MS__AND2_8%B N_B_M1003_g N_B_M1005_g N_B_c_261_n
+ N_B_c_262_n B PM_SKY130_OSU_SC_15T_MS__AND2_8%B
x_PM_SKY130_OSU_SC_15T_MS__AND2_8%A_27_115# N_A_27_115#_M1007_s
+ N_A_27_115#_M1010_d N_A_27_115#_M1002_g N_A_27_115#_c_369_n
+ N_A_27_115#_M1000_g N_A_27_115#_c_301_n N_A_27_115#_c_302_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_374_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_307_n N_A_27_115#_c_309_n N_A_27_115#_c_310_n
+ N_A_27_115#_M1009_g N_A_27_115#_c_381_n N_A_27_115#_M1004_g
+ N_A_27_115#_c_315_n N_A_27_115#_c_316_n N_A_27_115#_M1012_g
+ N_A_27_115#_c_386_n N_A_27_115#_M1006_g N_A_27_115#_c_321_n
+ N_A_27_115#_c_323_n N_A_27_115#_M1014_g N_A_27_115#_c_328_n
+ N_A_27_115#_c_392_n N_A_27_115#_M1011_g N_A_27_115#_c_329_n
+ N_A_27_115#_c_330_n N_A_27_115#_M1015_g N_A_27_115#_c_397_n
+ N_A_27_115#_M1013_g N_A_27_115#_c_335_n N_A_27_115#_c_337_n
+ N_A_27_115#_M1016_g N_A_27_115#_c_403_n N_A_27_115#_M1018_g
+ N_A_27_115#_c_342_n N_A_27_115#_c_343_n N_A_27_115#_M1017_g
+ N_A_27_115#_c_408_n N_A_27_115#_M1019_g N_A_27_115#_c_348_n
+ N_A_27_115#_c_349_n N_A_27_115#_c_350_n N_A_27_115#_c_351_n
+ N_A_27_115#_c_352_n N_A_27_115#_c_353_n N_A_27_115#_c_354_n
+ N_A_27_115#_c_355_n N_A_27_115#_c_356_n N_A_27_115#_c_357_n
+ N_A_27_115#_c_358_n N_A_27_115#_c_359_n N_A_27_115#_c_360_n
+ N_A_27_115#_c_363_n N_A_27_115#_c_364_n N_A_27_115#_c_419_n
+ N_A_27_115#_c_365_n N_A_27_115#_c_367_n N_A_27_115#_c_368_n
+ N_A_27_115#_c_435_n PM_SKY130_OSU_SC_15T_MS__AND2_8%A_27_115#
x_PM_SKY130_OSU_SC_15T_MS__AND2_8%Y N_Y_M1002_d N_Y_M1009_d N_Y_M1014_d
+ N_Y_M1016_d N_Y_M1000_s N_Y_M1004_s N_Y_M1011_s N_Y_M1018_s N_Y_c_538_n
+ N_Y_c_543_n N_Y_c_544_n N_Y_c_549_n N_Y_c_550_n N_Y_c_555_n N_Y_c_556_n
+ N_Y_c_560_n N_Y_c_561_n N_Y_c_564_n Y N_Y_c_566_n N_Y_c_568_n N_Y_c_569_n
+ N_Y_c_570_n N_Y_c_572_n N_Y_c_575_n N_Y_c_576_n N_Y_c_577_n N_Y_c_580_n
+ N_Y_c_581_n N_Y_c_582_n N_Y_c_583_n N_Y_c_586_n N_Y_c_587_n
+ PM_SKY130_OSU_SC_15T_MS__AND2_8%Y
cc_1 N_GND_M1007_b N_A_M1007_g 0.0806078f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1007_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_A_M1007_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1007_b N_A_c_227_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.505
cc_5 N_GND_M1007_b N_A_c_228_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.505
cc_6 N_GND_M1007_b N_B_M1003_g 0.0460664f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_7 N_GND_c_2_p N_B_M1003_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.945
cc_8 N_GND_c_8_p N_B_M1003_g 0.00319969f $X=1.05 $Y=0.74 $X2=0.835 $Y2=0.945
cc_9 N_GND_c_3_p N_B_M1003_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.835 $Y2=0.945
cc_10 N_GND_M1007_b N_B_M1005_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_11 N_GND_M1007_b N_B_c_261_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.165
cc_12 N_GND_M1007_b N_B_c_262_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.165
cc_13 N_GND_M1007_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.7
cc_14 N_GND_M1007_b N_A_27_115#_M1002_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.945
cc_15 N_GND_c_8_p N_A_27_115#_M1002_g 0.00883341f $X=1.05 $Y=0.74 $X2=1.335
+ $Y2=0.945
cc_16 N_GND_c_16_p N_A_27_115#_M1002_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.945
cc_17 N_GND_c_3_p N_A_27_115#_M1002_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.335
+ $Y2=0.945
cc_18 N_GND_M1007_b N_A_27_115#_c_301_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.55
cc_19 N_GND_M1007_b N_A_27_115#_c_302_n 0.00727817f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.625
cc_20 N_GND_M1007_b N_A_27_115#_M1008_g 0.0202142f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.945
cc_21 N_GND_c_16_p N_A_27_115#_M1008_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.945
cc_22 N_GND_c_22_p N_A_27_115#_M1008_g 0.00327323f $X=1.98 $Y=0.74 $X2=1.765
+ $Y2=0.945
cc_23 N_GND_c_3_p N_A_27_115#_M1008_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.765
+ $Y2=0.945
cc_24 N_GND_M1007_b N_A_27_115#_c_307_n 0.0179436f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_25 N_GND_c_22_p N_A_27_115#_c_307_n 0.00291042f $X=1.98 $Y=0.74 $X2=2.12
+ $Y2=1.585
cc_26 N_GND_M1007_b N_A_27_115#_c_309_n 0.0456099f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.585
cc_27 N_GND_M1007_b N_A_27_115#_c_310_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.625
cc_28 N_GND_M1007_b N_A_27_115#_M1009_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.945
cc_29 N_GND_c_22_p N_A_27_115#_M1009_g 0.00327323f $X=1.98 $Y=0.74 $X2=2.195
+ $Y2=0.945
cc_30 N_GND_c_30_p N_A_27_115#_M1009_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.945
cc_31 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=4.42 $Y=0.19 $X2=2.195
+ $Y2=0.945
cc_32 N_GND_M1007_b N_A_27_115#_c_315_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.585
cc_33 N_GND_M1007_b N_A_27_115#_c_316_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.625
cc_34 N_GND_M1007_b N_A_27_115#_M1012_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.945
cc_35 N_GND_c_30_p N_A_27_115#_M1012_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.945
cc_36 N_GND_c_36_p N_A_27_115#_M1012_g 0.00327323f $X=2.84 $Y=0.74 $X2=2.625
+ $Y2=0.945
cc_37 N_GND_c_3_p N_A_27_115#_M1012_g 0.00468827f $X=4.42 $Y=0.19 $X2=2.625
+ $Y2=0.945
cc_38 N_GND_M1007_b N_A_27_115#_c_321_n 0.0179436f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.585
cc_39 N_GND_c_36_p N_A_27_115#_c_321_n 0.00291042f $X=2.84 $Y=0.74 $X2=2.98
+ $Y2=1.585
cc_40 N_GND_M1007_b N_A_27_115#_c_323_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.625
cc_41 N_GND_M1007_b N_A_27_115#_M1014_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.945
cc_42 N_GND_c_36_p N_A_27_115#_M1014_g 0.00327323f $X=2.84 $Y=0.74 $X2=3.055
+ $Y2=0.945
cc_43 N_GND_c_43_p N_A_27_115#_M1014_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.055
+ $Y2=0.945
cc_44 N_GND_c_3_p N_A_27_115#_M1014_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.055
+ $Y2=0.945
cc_45 N_GND_M1007_b N_A_27_115#_c_328_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.55
cc_46 N_GND_M1007_b N_A_27_115#_c_329_n 0.0180386f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.585
cc_47 N_GND_M1007_b N_A_27_115#_c_330_n 0.0118833f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.625
cc_48 N_GND_M1007_b N_A_27_115#_M1015_g 0.020212f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=0.945
cc_49 N_GND_c_43_p N_A_27_115#_M1015_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.485
+ $Y2=0.945
cc_50 N_GND_c_50_p N_A_27_115#_M1015_g 0.00327323f $X=3.7 $Y=0.74 $X2=3.485
+ $Y2=0.945
cc_51 N_GND_c_3_p N_A_27_115#_M1015_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.485
+ $Y2=0.945
cc_52 N_GND_M1007_b N_A_27_115#_c_335_n 0.0179436f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.585
cc_53 N_GND_c_50_p N_A_27_115#_c_335_n 0.00291042f $X=3.7 $Y=0.74 $X2=3.84
+ $Y2=1.585
cc_54 N_GND_M1007_b N_A_27_115#_c_337_n 0.013058f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.625
cc_55 N_GND_M1007_b N_A_27_115#_M1016_g 0.020212f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=0.945
cc_56 N_GND_c_50_p N_A_27_115#_M1016_g 0.00327323f $X=3.7 $Y=0.74 $X2=3.915
+ $Y2=0.945
cc_57 N_GND_c_57_p N_A_27_115#_M1016_g 0.00606474f $X=4.475 $Y=0.152 $X2=3.915
+ $Y2=0.945
cc_58 N_GND_c_3_p N_A_27_115#_M1016_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.915
+ $Y2=0.945
cc_59 N_GND_M1007_b N_A_27_115#_c_342_n 0.0369419f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=1.585
cc_60 N_GND_M1007_b N_A_27_115#_c_343_n 0.0268552f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=2.625
cc_61 N_GND_M1007_b N_A_27_115#_M1017_g 0.0264941f $X=-0.045 $Y=0 $X2=4.345
+ $Y2=0.945
cc_62 N_GND_c_57_p N_A_27_115#_M1017_g 0.00606474f $X=4.475 $Y=0.152 $X2=4.345
+ $Y2=0.945
cc_63 N_GND_c_63_p N_A_27_115#_M1017_g 0.00502587f $X=4.56 $Y=0.74 $X2=4.345
+ $Y2=0.945
cc_64 N_GND_c_3_p N_A_27_115#_M1017_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.345
+ $Y2=0.945
cc_65 N_GND_M1007_b N_A_27_115#_c_348_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.625
cc_66 N_GND_M1007_b N_A_27_115#_c_349_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.625
cc_67 N_GND_M1007_b N_A_27_115#_c_350_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.585
cc_68 N_GND_M1007_b N_A_27_115#_c_351_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.625
cc_69 N_GND_M1007_b N_A_27_115#_c_352_n 0.00873941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.585
cc_70 N_GND_M1007_b N_A_27_115#_c_353_n 0.00735657f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.625
cc_71 N_GND_M1007_b N_A_27_115#_c_354_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.585
cc_72 N_GND_M1007_b N_A_27_115#_c_355_n 0.00151234f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.625
cc_73 N_GND_M1007_b N_A_27_115#_c_356_n 0.00873941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.585
cc_74 N_GND_M1007_b N_A_27_115#_c_357_n 0.00735657f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.625
cc_75 N_GND_M1007_b N_A_27_115#_c_358_n 0.00873941f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=1.585
cc_76 N_GND_M1007_b N_A_27_115#_c_359_n 0.00735657f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=2.625
cc_77 N_GND_M1007_b N_A_27_115#_c_360_n 0.0143389f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_78 N_GND_c_2_p N_A_27_115#_c_360_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_79 N_GND_c_3_p N_A_27_115#_c_360_n 0.00476261f $X=4.42 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_80 N_GND_M1007_b N_A_27_115#_c_363_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.675
cc_81 N_GND_M1007_b N_A_27_115#_c_364_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.675
cc_82 N_GND_M1007_b N_A_27_115#_c_365_n 0.0227928f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_83 N_GND_c_8_p N_A_27_115#_c_365_n 0.00833003f $X=1.05 $Y=0.74 $X2=1.43
+ $Y2=1.675
cc_84 N_GND_M1007_b N_A_27_115#_c_367_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.675
cc_85 N_GND_M1007_b N_A_27_115#_c_368_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.305
cc_86 N_GND_M1007_b N_Y_c_538_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.74
cc_87 N_GND_c_8_p N_Y_c_538_n 0.0150458f $X=1.05 $Y=0.74 $X2=1.55 $Y2=0.74
cc_88 N_GND_c_16_p N_Y_c_538_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.74
cc_89 N_GND_c_22_p N_Y_c_538_n 0.0029082f $X=1.98 $Y=0.74 $X2=1.55 $Y2=0.74
cc_90 N_GND_c_3_p N_Y_c_538_n 0.00475776f $X=4.42 $Y=0.19 $X2=1.55 $Y2=0.74
cc_91 N_GND_M1007_b N_Y_c_543_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_92 N_GND_M1007_b N_Y_c_544_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.74
cc_93 N_GND_c_22_p N_Y_c_544_n 0.0029082f $X=1.98 $Y=0.74 $X2=2.41 $Y2=0.74
cc_94 N_GND_c_30_p N_Y_c_544_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.74
cc_95 N_GND_c_36_p N_Y_c_544_n 0.0029082f $X=2.84 $Y=0.74 $X2=2.41 $Y2=0.74
cc_96 N_GND_c_3_p N_Y_c_544_n 0.00475776f $X=4.42 $Y=0.19 $X2=2.41 $Y2=0.74
cc_97 N_GND_M1007_b N_Y_c_549_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.33
cc_98 N_GND_M1007_b N_Y_c_550_n 0.00155118f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.74
cc_99 N_GND_c_36_p N_Y_c_550_n 0.0029082f $X=2.84 $Y=0.74 $X2=3.27 $Y2=0.74
cc_100 N_GND_c_43_p N_Y_c_550_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.74
cc_101 N_GND_c_50_p N_Y_c_550_n 0.0029082f $X=3.7 $Y=0.74 $X2=3.27 $Y2=0.74
cc_102 N_GND_c_3_p N_Y_c_550_n 0.00475776f $X=4.42 $Y=0.19 $X2=3.27 $Y2=0.74
cc_103 N_GND_M1007_b N_Y_c_555_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.33
cc_104 N_GND_M1007_b N_Y_c_556_n 0.00155118f $X=-0.045 $Y=0 $X2=4.13 $Y2=0.74
cc_105 N_GND_c_50_p N_Y_c_556_n 0.0029082f $X=3.7 $Y=0.74 $X2=4.13 $Y2=0.74
cc_106 N_GND_c_57_p N_Y_c_556_n 0.0075556f $X=4.475 $Y=0.152 $X2=4.13 $Y2=0.74
cc_107 N_GND_c_3_p N_Y_c_556_n 0.00475776f $X=4.42 $Y=0.19 $X2=4.13 $Y2=0.74
cc_108 N_GND_M1007_b N_Y_c_560_n 0.0152877f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.33
cc_109 N_GND_M1007_b N_Y_c_561_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.335
cc_110 N_GND_c_8_p N_Y_c_561_n 0.00377613f $X=1.05 $Y=0.74 $X2=1.55 $Y2=1.335
cc_111 N_GND_c_22_p N_Y_c_561_n 7.53951e-19 $X=1.98 $Y=0.74 $X2=1.55 $Y2=1.335
cc_112 N_GND_M1007_b N_Y_c_564_n 0.00509006f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.215
cc_113 N_GND_M1007_b Y 0.0306813f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.96
cc_114 N_GND_M1008_s N_Y_c_566_n 0.0127109f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.22
cc_115 N_GND_c_22_p N_Y_c_566_n 0.0175563f $X=1.98 $Y=0.74 $X2=2.265 $Y2=1.22
cc_116 N_GND_M1007_b N_Y_c_568_n 0.0188475f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.33
cc_117 N_GND_M1007_b N_Y_c_569_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.215
cc_118 N_GND_M1012_s N_Y_c_570_n 0.0127109f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.22
cc_119 N_GND_c_36_p N_Y_c_570_n 0.0175563f $X=2.84 $Y=0.74 $X2=3.125 $Y2=1.22
cc_120 N_GND_M1007_b N_Y_c_572_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.22
cc_121 N_GND_c_22_p N_Y_c_572_n 7.53951e-19 $X=1.98 $Y=0.74 $X2=2.555 $Y2=1.22
cc_122 N_GND_c_36_p N_Y_c_572_n 7.53951e-19 $X=2.84 $Y=0.74 $X2=2.555 $Y2=1.22
cc_123 N_GND_M1007_b N_Y_c_575_n 0.0144616f $X=-0.045 $Y=0 $X2=3.125 $Y2=2.33
cc_124 N_GND_M1007_b N_Y_c_576_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.33
cc_125 N_GND_M1007_b N_Y_c_577_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.335
cc_126 N_GND_c_36_p N_Y_c_577_n 7.53951e-19 $X=2.84 $Y=0.74 $X2=3.27 $Y2=1.335
cc_127 N_GND_c_50_p N_Y_c_577_n 0.00113348f $X=3.7 $Y=0.74 $X2=3.27 $Y2=1.335
cc_128 N_GND_M1007_b N_Y_c_580_n 0.0358528f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.215
cc_129 N_GND_M1007_b N_Y_c_581_n 0.0188475f $X=-0.045 $Y=0 $X2=3.985 $Y2=2.33
cc_130 N_GND_M1007_b N_Y_c_582_n 0.00584404f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.33
cc_131 N_GND_M1007_b N_Y_c_583_n 0.00409378f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.335
cc_132 N_GND_c_50_p N_Y_c_583_n 7.53951e-19 $X=3.7 $Y=0.74 $X2=4.13 $Y2=1.335
cc_133 N_GND_c_63_p N_Y_c_583_n 0.00402079f $X=4.56 $Y=0.74 $X2=4.13 $Y2=1.335
cc_134 N_GND_M1007_b N_Y_c_586_n 0.06145f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.215
cc_135 N_GND_M1015_s N_Y_c_587_n 0.0127109f $X=3.56 $Y=0.575 $X2=4.13 $Y2=1.22
cc_136 N_GND_c_50_p N_Y_c_587_n 0.0166405f $X=3.7 $Y=0.74 $X2=4.13 $Y2=1.22
cc_137 N_VDD_M1010_b N_A_M1010_g 0.0193382f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_138 N_VDD_c_138_p N_A_M1010_g 0.00713292f $X=0.26 $Y=3.895 $X2=0.475
+ $Y2=3.825
cc_139 N_VDD_c_139_p N_A_M1010_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_140 N_VDD_c_140_p N_A_M1010_g 0.00429146f $X=4.42 $Y=5.36 $X2=0.475 $Y2=3.825
cc_141 N_VDD_M1010_b N_A_c_227_n 0.0111025f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=2.505
cc_142 N_VDD_M1010_s N_A_c_228_n 0.0127742f $X=0.135 $Y=2.825 $X2=0.27 $Y2=2.505
cc_143 N_VDD_M1010_b N_A_c_228_n 0.00612103f $X=-0.045 $Y=2.645 $X2=0.27
+ $Y2=2.505
cc_144 N_VDD_c_138_p N_A_c_228_n 0.00352433f $X=0.26 $Y=3.895 $X2=0.27 $Y2=2.505
cc_145 N_VDD_M1010_s A 0.00746694f $X=0.135 $Y=2.825 $X2=0.275 $Y2=3.07
cc_146 N_VDD_M1010_b A 0.00970321f $X=-0.045 $Y=2.645 $X2=0.275 $Y2=3.07
cc_147 N_VDD_c_138_p A 0.00428937f $X=0.26 $Y=3.895 $X2=0.275 $Y2=3.07
cc_148 N_VDD_M1010_b N_B_M1005_g 0.0191387f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_149 N_VDD_c_139_p N_B_M1005_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905
+ $Y2=3.825
cc_150 N_VDD_c_150_p N_B_M1005_g 0.00354579f $X=1.12 $Y=3.555 $X2=0.905
+ $Y2=3.825
cc_151 N_VDD_c_140_p N_B_M1005_g 0.00429146f $X=4.42 $Y=5.36 $X2=0.905 $Y2=3.825
cc_152 N_VDD_M1010_b N_B_c_262_n 0.00170274f $X=-0.045 $Y=2.645 $X2=0.95
+ $Y2=2.165
cc_153 N_VDD_M1010_b B 0.00860092f $X=-0.045 $Y=2.645 $X2=0.955 $Y2=2.7
cc_154 N_VDD_c_150_p B 0.00236322f $X=1.12 $Y=3.555 $X2=0.955 $Y2=2.7
cc_155 N_VDD_M1010_b N_A_27_115#_c_369_n 0.0174951f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.7
cc_156 N_VDD_c_150_p N_A_27_115#_c_369_n 0.00354579f $X=1.12 $Y=3.555 $X2=1.335
+ $Y2=2.7
cc_157 N_VDD_c_157_p N_A_27_115#_c_369_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335
+ $Y2=2.7
cc_158 N_VDD_c_140_p N_A_27_115#_c_369_n 0.00429146f $X=4.42 $Y=5.36 $X2=1.335
+ $Y2=2.7
cc_159 N_VDD_M1010_b N_A_27_115#_c_302_n 0.00427883f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_160 N_VDD_M1010_b N_A_27_115#_c_374_n 0.0173909f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.7
cc_161 N_VDD_c_150_p N_A_27_115#_c_374_n 3.67508e-19 $X=1.12 $Y=3.555 $X2=1.765
+ $Y2=2.7
cc_162 N_VDD_c_157_p N_A_27_115#_c_374_n 0.00500229f $X=1.895 $Y=5.397 $X2=1.765
+ $Y2=2.7
cc_163 N_VDD_c_163_p N_A_27_115#_c_374_n 0.00373985f $X=1.98 $Y=3.215 $X2=1.765
+ $Y2=2.7
cc_164 N_VDD_c_140_p N_A_27_115#_c_374_n 0.00430409f $X=4.42 $Y=5.36 $X2=1.765
+ $Y2=2.7
cc_165 N_VDD_M1010_b N_A_27_115#_c_310_n 0.00399373f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.625
cc_166 N_VDD_c_163_p N_A_27_115#_c_310_n 0.0037128f $X=1.98 $Y=3.215 $X2=2.12
+ $Y2=2.625
cc_167 N_VDD_M1010_b N_A_27_115#_c_381_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.7
cc_168 N_VDD_c_163_p N_A_27_115#_c_381_n 0.00354579f $X=1.98 $Y=3.215 $X2=2.195
+ $Y2=2.7
cc_169 N_VDD_c_169_p N_A_27_115#_c_381_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.195
+ $Y2=2.7
cc_170 N_VDD_c_140_p N_A_27_115#_c_381_n 0.00429146f $X=4.42 $Y=5.36 $X2=2.195
+ $Y2=2.7
cc_171 N_VDD_M1010_b N_A_27_115#_c_316_n 0.00448664f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.625
cc_172 N_VDD_M1010_b N_A_27_115#_c_386_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.7
cc_173 N_VDD_c_169_p N_A_27_115#_c_386_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.625
+ $Y2=2.7
cc_174 N_VDD_c_174_p N_A_27_115#_c_386_n 0.00354579f $X=2.84 $Y=3.215 $X2=2.625
+ $Y2=2.7
cc_175 N_VDD_c_140_p N_A_27_115#_c_386_n 0.00429146f $X=4.42 $Y=5.36 $X2=2.625
+ $Y2=2.7
cc_176 N_VDD_M1010_b N_A_27_115#_c_323_n 0.00399373f $X=-0.045 $Y=2.645 $X2=2.98
+ $Y2=2.625
cc_177 N_VDD_c_174_p N_A_27_115#_c_323_n 0.0037128f $X=2.84 $Y=3.215 $X2=2.98
+ $Y2=2.625
cc_178 N_VDD_M1010_b N_A_27_115#_c_392_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.055
+ $Y2=2.7
cc_179 N_VDD_c_174_p N_A_27_115#_c_392_n 0.00354579f $X=2.84 $Y=3.215 $X2=3.055
+ $Y2=2.7
cc_180 N_VDD_c_180_p N_A_27_115#_c_392_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.055
+ $Y2=2.7
cc_181 N_VDD_c_140_p N_A_27_115#_c_392_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.055
+ $Y2=2.7
cc_182 N_VDD_M1010_b N_A_27_115#_c_330_n 0.00448664f $X=-0.045 $Y=2.645 $X2=3.41
+ $Y2=2.625
cc_183 N_VDD_M1010_b N_A_27_115#_c_397_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.485
+ $Y2=2.7
cc_184 N_VDD_c_180_p N_A_27_115#_c_397_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.485
+ $Y2=2.7
cc_185 N_VDD_c_185_p N_A_27_115#_c_397_n 0.00354579f $X=3.7 $Y=3.215 $X2=3.485
+ $Y2=2.7
cc_186 N_VDD_c_140_p N_A_27_115#_c_397_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.485
+ $Y2=2.7
cc_187 N_VDD_M1010_b N_A_27_115#_c_337_n 0.00399373f $X=-0.045 $Y=2.645 $X2=3.84
+ $Y2=2.625
cc_188 N_VDD_c_185_p N_A_27_115#_c_337_n 0.0037128f $X=3.7 $Y=3.215 $X2=3.84
+ $Y2=2.625
cc_189 N_VDD_M1010_b N_A_27_115#_c_403_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.915
+ $Y2=2.7
cc_190 N_VDD_c_185_p N_A_27_115#_c_403_n 0.00354579f $X=3.7 $Y=3.215 $X2=3.915
+ $Y2=2.7
cc_191 N_VDD_c_191_p N_A_27_115#_c_403_n 0.00496961f $X=4.475 $Y=5.397 $X2=3.915
+ $Y2=2.7
cc_192 N_VDD_c_140_p N_A_27_115#_c_403_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.915
+ $Y2=2.7
cc_193 N_VDD_M1010_b N_A_27_115#_c_343_n 0.00840215f $X=-0.045 $Y=2.645 $X2=4.27
+ $Y2=2.625
cc_194 N_VDD_M1010_b N_A_27_115#_c_408_n 0.0212947f $X=-0.045 $Y=2.645 $X2=4.345
+ $Y2=2.7
cc_195 N_VDD_c_191_p N_A_27_115#_c_408_n 0.00496961f $X=4.475 $Y=5.397 $X2=4.345
+ $Y2=2.7
cc_196 N_VDD_c_196_p N_A_27_115#_c_408_n 0.00713292f $X=4.56 $Y=3.215 $X2=4.345
+ $Y2=2.7
cc_197 N_VDD_c_140_p N_A_27_115#_c_408_n 0.00429146f $X=4.42 $Y=5.36 $X2=4.345
+ $Y2=2.7
cc_198 N_VDD_M1010_b N_A_27_115#_c_348_n 0.0021704f $X=-0.045 $Y=2.645 $X2=1.352
+ $Y2=2.625
cc_199 N_VDD_M1010_b N_A_27_115#_c_349_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=1.765 $Y2=2.625
cc_200 N_VDD_M1010_b N_A_27_115#_c_351_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.195 $Y2=2.625
cc_201 N_VDD_M1010_b N_A_27_115#_c_353_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.625 $Y2=2.625
cc_202 N_VDD_M1010_b N_A_27_115#_c_355_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.055 $Y2=2.625
cc_203 N_VDD_M1010_b N_A_27_115#_c_357_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.485 $Y2=2.625
cc_204 N_VDD_M1010_b N_A_27_115#_c_359_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.915 $Y2=2.625
cc_205 N_VDD_M1010_b N_A_27_115#_c_419_n 0.00198641f $X=-0.045 $Y=2.645 $X2=0.69
+ $Y2=3.555
cc_206 N_VDD_c_139_p N_A_27_115#_c_419_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69
+ $Y2=3.555
cc_207 N_VDD_c_140_p N_A_27_115#_c_419_n 0.00434939f $X=4.42 $Y=5.36 $X2=0.69
+ $Y2=3.555
cc_208 N_VDD_M1010_b N_A_27_115#_c_368_n 8.22047e-19 $X=-0.045 $Y=2.645 $X2=0.65
+ $Y2=3.305
cc_209 N_VDD_M1010_b N_Y_c_543_n 0.00388477f $X=-0.045 $Y=2.645 $X2=1.55
+ $Y2=2.33
cc_210 N_VDD_c_157_p N_Y_c_543_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.33
cc_211 N_VDD_c_140_p N_Y_c_543_n 0.00434939f $X=4.42 $Y=5.36 $X2=1.55 $Y2=2.33
cc_212 N_VDD_M1010_b N_Y_c_549_n 0.0042387f $X=-0.045 $Y=2.645 $X2=2.41 $Y2=2.33
cc_213 N_VDD_c_169_p N_Y_c_549_n 0.0045126f $X=2.755 $Y=5.397 $X2=2.41 $Y2=2.33
cc_214 N_VDD_c_140_p N_Y_c_549_n 0.00434939f $X=4.42 $Y=5.36 $X2=2.41 $Y2=2.33
cc_215 N_VDD_M1010_b N_Y_c_555_n 0.0042387f $X=-0.045 $Y=2.645 $X2=3.27 $Y2=2.33
cc_216 N_VDD_c_180_p N_Y_c_555_n 0.00464147f $X=3.615 $Y=5.397 $X2=3.27 $Y2=2.33
cc_217 N_VDD_c_140_p N_Y_c_555_n 0.00434939f $X=4.42 $Y=5.36 $X2=3.27 $Y2=2.33
cc_218 N_VDD_M1010_b N_Y_c_560_n 0.0042387f $X=-0.045 $Y=2.645 $X2=4.13 $Y2=2.33
cc_219 N_VDD_c_191_p N_Y_c_560_n 0.00475585f $X=4.475 $Y=5.397 $X2=4.13 $Y2=2.33
cc_220 N_VDD_c_140_p N_Y_c_560_n 0.00434939f $X=4.42 $Y=5.36 $X2=4.13 $Y2=2.33
cc_221 N_VDD_c_163_p N_Y_c_568_n 0.00622932f $X=1.98 $Y=3.215 $X2=2.265 $Y2=2.33
cc_222 N_VDD_c_174_p N_Y_c_575_n 0.00622932f $X=2.84 $Y=3.215 $X2=3.125 $Y2=2.33
cc_223 N_VDD_c_185_p N_Y_c_581_n 0.00622932f $X=3.7 $Y=3.215 $X2=3.985 $Y2=2.33
cc_224 N_A_M1007_g N_B_M1003_g 0.113664f $X=0.475 $Y=0.945 $X2=0.835 $Y2=0.945
cc_225 N_A_M1007_g N_B_M1005_g 0.0506107f $X=0.475 $Y=0.945 $X2=0.905 $Y2=3.825
cc_226 N_A_M1007_g N_B_c_262_n 7.8234e-19 $X=0.475 $Y=0.945 $X2=0.95 $Y2=2.165
cc_227 N_A_M1007_g N_A_27_115#_c_360_n 0.0114001f $X=0.475 $Y=0.945 $X2=0.26
+ $Y2=0.74
cc_228 N_A_M1007_g N_A_27_115#_c_363_n 0.0160984f $X=0.475 $Y=0.945 $X2=0.525
+ $Y2=1.675
cc_229 N_A_c_227_n N_A_27_115#_c_363_n 0.00117122f $X=0.475 $Y=2.505 $X2=0.525
+ $Y2=1.675
cc_230 N_A_c_228_n N_A_27_115#_c_363_n 2.65873e-19 $X=0.27 $Y=2.505 $X2=0.525
+ $Y2=1.675
cc_231 N_A_c_227_n N_A_27_115#_c_364_n 0.00133457f $X=0.475 $Y=2.505 $X2=0.345
+ $Y2=1.675
cc_232 N_A_c_228_n N_A_27_115#_c_364_n 0.0055861f $X=0.27 $Y=2.505 $X2=0.345
+ $Y2=1.675
cc_233 N_A_M1007_g N_A_27_115#_c_367_n 0.00322084f $X=0.475 $Y=0.945 $X2=0.61
+ $Y2=1.675
cc_234 N_A_M1007_g N_A_27_115#_c_368_n 0.0265302f $X=0.475 $Y=0.945 $X2=0.65
+ $Y2=3.305
cc_235 N_A_M1010_g N_A_27_115#_c_368_n 0.0149699f $X=0.475 $Y=3.825 $X2=0.65
+ $Y2=3.305
cc_236 N_A_c_227_n N_A_27_115#_c_368_n 0.00766302f $X=0.475 $Y=2.505 $X2=0.65
+ $Y2=3.305
cc_237 N_A_c_228_n N_A_27_115#_c_368_n 0.0456533f $X=0.27 $Y=2.505 $X2=0.65
+ $Y2=3.305
cc_238 A N_A_27_115#_c_368_n 0.00758489f $X=0.275 $Y=3.07 $X2=0.65 $Y2=3.305
cc_239 N_A_M1010_g N_A_27_115#_c_435_n 0.00884152f $X=0.475 $Y=3.825 $X2=0.65
+ $Y2=3.475
cc_240 N_B_M1003_g N_A_27_115#_M1002_g 0.0276217f $X=0.835 $Y=0.945 $X2=1.335
+ $Y2=0.945
cc_241 N_B_M1005_g N_A_27_115#_c_301_n 0.00773101f $X=0.905 $Y=3.825 $X2=1.37
+ $Y2=2.55
cc_242 N_B_c_261_n N_A_27_115#_c_301_n 0.0206104f $X=0.95 $Y=2.165 $X2=1.37
+ $Y2=2.55
cc_243 N_B_c_262_n N_A_27_115#_c_301_n 0.0033451f $X=0.95 $Y=2.165 $X2=1.37
+ $Y2=2.55
cc_244 N_B_M1003_g N_A_27_115#_c_309_n 0.0104742f $X=0.835 $Y=0.945 $X2=1.84
+ $Y2=1.585
cc_245 N_B_M1005_g N_A_27_115#_c_348_n 0.0410292f $X=0.905 $Y=3.825 $X2=1.352
+ $Y2=2.625
cc_246 N_B_c_262_n N_A_27_115#_c_348_n 0.00173699f $X=0.95 $Y=2.165 $X2=1.352
+ $Y2=2.625
cc_247 B N_A_27_115#_c_348_n 0.00389258f $X=0.955 $Y=2.7 $X2=1.352 $Y2=2.625
cc_248 N_B_M1003_g N_A_27_115#_c_365_n 0.0182215f $X=0.835 $Y=0.945 $X2=1.43
+ $Y2=1.675
cc_249 N_B_c_261_n N_A_27_115#_c_365_n 0.00258465f $X=0.95 $Y=2.165 $X2=1.43
+ $Y2=1.675
cc_250 N_B_c_262_n N_A_27_115#_c_365_n 0.0101796f $X=0.95 $Y=2.165 $X2=1.43
+ $Y2=1.675
cc_251 N_B_M1003_g N_A_27_115#_c_368_n 0.00755919f $X=0.835 $Y=0.945 $X2=0.65
+ $Y2=3.305
cc_252 N_B_M1005_g N_A_27_115#_c_368_n 0.0137515f $X=0.905 $Y=3.825 $X2=0.65
+ $Y2=3.305
cc_253 N_B_c_262_n N_A_27_115#_c_368_n 0.0541375f $X=0.95 $Y=2.165 $X2=0.65
+ $Y2=3.305
cc_254 B N_A_27_115#_c_368_n 0.00866797f $X=0.955 $Y=2.7 $X2=0.65 $Y2=3.305
cc_255 B N_A_27_115#_c_435_n 0.00281588f $X=0.955 $Y=2.7 $X2=0.65 $Y2=3.475
cc_256 N_B_c_262_n N_Y_c_543_n 0.0149875f $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.33
cc_257 B N_Y_c_543_n 0.00649253f $X=0.955 $Y=2.7 $X2=1.55 $Y2=2.33
cc_258 N_B_M1003_g N_Y_c_561_n 3.57178e-19 $X=0.835 $Y=0.945 $X2=1.55 $Y2=1.335
cc_259 N_B_c_261_n N_Y_c_564_n 5.85867e-19 $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.215
cc_260 N_B_c_262_n N_Y_c_564_n 0.00592261f $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.215
cc_261 N_B_M1003_g Y 6.71108e-19 $X=0.835 $Y=0.945 $X2=1.555 $Y2=1.96
cc_262 N_B_c_262_n Y 0.00695761f $X=0.95 $Y=2.165 $X2=1.555 $Y2=1.96
cc_263 N_A_27_115#_M1002_g N_Y_c_538_n 9.07985e-19 $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=0.74
cc_264 N_A_27_115#_M1008_g N_Y_c_538_n 8.52215e-19 $X=1.765 $Y=0.945 $X2=1.55
+ $Y2=0.74
cc_265 N_A_27_115#_c_309_n N_Y_c_538_n 0.00171364f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=0.74
cc_266 N_A_27_115#_c_365_n N_Y_c_538_n 0.00500271f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.74
cc_267 N_A_27_115#_c_369_n N_Y_c_543_n 0.00287202f $X=1.335 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_268 N_A_27_115#_c_301_n N_Y_c_543_n 0.00744772f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_269 N_A_27_115#_c_302_n N_Y_c_543_n 0.0156184f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_270 N_A_27_115#_c_374_n N_Y_c_543_n 0.00401146f $X=1.765 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_271 N_A_27_115#_c_309_n N_Y_c_543_n 0.00182797f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.33
cc_272 N_A_27_115#_c_365_n N_Y_c_543_n 0.00273485f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_273 N_A_27_115#_M1009_g N_Y_c_544_n 8.52215e-19 $X=2.195 $Y=0.945 $X2=2.41
+ $Y2=0.74
cc_274 N_A_27_115#_c_315_n N_Y_c_544_n 0.00280419f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=0.74
cc_275 N_A_27_115#_M1012_g N_Y_c_544_n 8.52215e-19 $X=2.625 $Y=0.945 $X2=2.41
+ $Y2=0.74
cc_276 N_A_27_115#_c_381_n N_Y_c_549_n 0.00401146f $X=2.195 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_277 N_A_27_115#_c_315_n N_Y_c_549_n 0.00250559f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.33
cc_278 N_A_27_115#_c_316_n N_Y_c_549_n 0.021445f $X=2.55 $Y=2.625 $X2=2.41
+ $Y2=2.33
cc_279 N_A_27_115#_c_386_n N_Y_c_549_n 0.00401146f $X=2.625 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_280 N_A_27_115#_c_328_n N_Y_c_549_n 0.00361281f $X=3.055 $Y=2.55 $X2=2.41
+ $Y2=2.33
cc_281 N_A_27_115#_M1014_g N_Y_c_550_n 8.52215e-19 $X=3.055 $Y=0.945 $X2=3.27
+ $Y2=0.74
cc_282 N_A_27_115#_c_329_n N_Y_c_550_n 0.00280419f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=0.74
cc_283 N_A_27_115#_M1015_g N_Y_c_550_n 8.52215e-19 $X=3.485 $Y=0.945 $X2=3.27
+ $Y2=0.74
cc_284 N_A_27_115#_c_328_n N_Y_c_555_n 0.00721971f $X=3.055 $Y=2.55 $X2=3.27
+ $Y2=2.33
cc_285 N_A_27_115#_c_392_n N_Y_c_555_n 0.00401146f $X=3.055 $Y=2.7 $X2=3.27
+ $Y2=2.33
cc_286 N_A_27_115#_c_329_n N_Y_c_555_n 0.00250559f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=2.33
cc_287 N_A_27_115#_c_330_n N_Y_c_555_n 0.021445f $X=3.41 $Y=2.625 $X2=3.27
+ $Y2=2.33
cc_288 N_A_27_115#_c_397_n N_Y_c_555_n 0.00401146f $X=3.485 $Y=2.7 $X2=3.27
+ $Y2=2.33
cc_289 N_A_27_115#_M1016_g N_Y_c_556_n 8.52215e-19 $X=3.915 $Y=0.945 $X2=4.13
+ $Y2=0.74
cc_290 N_A_27_115#_c_342_n N_Y_c_556_n 0.00280419f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=0.74
cc_291 N_A_27_115#_M1017_g N_Y_c_556_n 8.52215e-19 $X=4.345 $Y=0.945 $X2=4.13
+ $Y2=0.74
cc_292 N_A_27_115#_c_403_n N_Y_c_560_n 0.00401146f $X=3.915 $Y=2.7 $X2=4.13
+ $Y2=2.33
cc_293 N_A_27_115#_c_342_n N_Y_c_560_n 0.00250559f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=2.33
cc_294 N_A_27_115#_c_343_n N_Y_c_560_n 0.0206674f $X=4.27 $Y=2.625 $X2=4.13
+ $Y2=2.33
cc_295 N_A_27_115#_c_408_n N_Y_c_560_n 0.00401146f $X=4.345 $Y=2.7 $X2=4.13
+ $Y2=2.33
cc_296 N_A_27_115#_M1002_g N_Y_c_561_n 0.00345902f $X=1.335 $Y=0.945 $X2=1.55
+ $Y2=1.335
cc_297 N_A_27_115#_M1008_g N_Y_c_561_n 0.00134358f $X=1.765 $Y=0.945 $X2=1.55
+ $Y2=1.335
cc_298 N_A_27_115#_c_365_n N_Y_c_561_n 0.00238892f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=1.335
cc_299 N_A_27_115#_c_301_n N_Y_c_564_n 0.00821104f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.215
cc_300 N_A_27_115#_c_302_n N_Y_c_564_n 0.00186325f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.215
cc_301 N_A_27_115#_c_309_n N_Y_c_564_n 0.00194187f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.215
cc_302 N_A_27_115#_c_365_n N_Y_c_564_n 0.00181779f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.215
cc_303 N_A_27_115#_M1002_g Y 0.00251111f $X=1.335 $Y=0.945 $X2=1.555 $Y2=1.96
cc_304 N_A_27_115#_c_301_n Y 0.00892438f $X=1.37 $Y=2.55 $X2=1.555 $Y2=1.96
cc_305 N_A_27_115#_M1008_g Y 0.00251111f $X=1.765 $Y=0.945 $X2=1.555 $Y2=1.96
cc_306 N_A_27_115#_c_309_n Y 0.0131748f $X=1.84 $Y=1.585 $X2=1.555 $Y2=1.96
cc_307 N_A_27_115#_c_365_n Y 0.0148238f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_308 N_A_27_115#_M1008_g N_Y_c_566_n 0.0120124f $X=1.765 $Y=0.945 $X2=2.265
+ $Y2=1.22
cc_309 N_A_27_115#_c_307_n N_Y_c_566_n 0.00213861f $X=2.12 $Y=1.585 $X2=2.265
+ $Y2=1.22
cc_310 N_A_27_115#_M1009_g N_Y_c_566_n 0.0120124f $X=2.195 $Y=0.945 $X2=2.265
+ $Y2=1.22
cc_311 N_A_27_115#_c_309_n N_Y_c_568_n 0.0121767f $X=1.84 $Y=1.585 $X2=2.265
+ $Y2=2.33
cc_312 N_A_27_115#_c_349_n N_Y_c_568_n 0.0158479f $X=1.765 $Y=2.625 $X2=2.265
+ $Y2=2.33
cc_313 N_A_27_115#_M1009_g N_Y_c_569_n 0.00251111f $X=2.195 $Y=0.945 $X2=2.41
+ $Y2=2.215
cc_314 N_A_27_115#_c_315_n N_Y_c_569_n 0.0177725f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_315 N_A_27_115#_M1012_g N_Y_c_569_n 0.00251111f $X=2.625 $Y=0.945 $X2=2.41
+ $Y2=2.215
cc_316 N_A_27_115#_c_328_n N_Y_c_569_n 0.00843025f $X=3.055 $Y=2.55 $X2=2.41
+ $Y2=2.215
cc_317 N_A_27_115#_M1012_g N_Y_c_570_n 0.0120124f $X=2.625 $Y=0.945 $X2=3.125
+ $Y2=1.22
cc_318 N_A_27_115#_c_321_n N_Y_c_570_n 0.00213861f $X=2.98 $Y=1.585 $X2=3.125
+ $Y2=1.22
cc_319 N_A_27_115#_M1014_g N_Y_c_570_n 0.0126623f $X=3.055 $Y=0.945 $X2=3.125
+ $Y2=1.22
cc_320 N_A_27_115#_M1009_g N_Y_c_572_n 0.00134358f $X=2.195 $Y=0.945 $X2=2.555
+ $Y2=1.22
cc_321 N_A_27_115#_M1012_g N_Y_c_572_n 0.00134358f $X=2.625 $Y=0.945 $X2=2.555
+ $Y2=1.22
cc_322 N_A_27_115#_c_328_n N_Y_c_575_n 0.0155956f $X=3.055 $Y=2.55 $X2=3.125
+ $Y2=2.33
cc_323 N_A_27_115#_c_352_n N_Y_c_575_n 0.00894336f $X=2.625 $Y=1.585 $X2=3.125
+ $Y2=2.33
cc_324 N_A_27_115#_c_353_n N_Y_c_575_n 0.00903839f $X=2.625 $Y=2.625 $X2=3.125
+ $Y2=2.33
cc_325 N_A_27_115#_c_315_n N_Y_c_576_n 0.00140336f $X=2.55 $Y=1.585 $X2=2.555
+ $Y2=2.33
cc_326 N_A_27_115#_c_328_n N_Y_c_576_n 0.0012308f $X=3.055 $Y=2.55 $X2=2.555
+ $Y2=2.33
cc_327 N_A_27_115#_c_350_n N_Y_c_576_n 0.00140336f $X=2.195 $Y=1.585 $X2=2.555
+ $Y2=2.33
cc_328 N_A_27_115#_c_351_n N_Y_c_576_n 0.00372651f $X=2.195 $Y=2.625 $X2=2.555
+ $Y2=2.33
cc_329 N_A_27_115#_M1014_g N_Y_c_577_n 0.00136818f $X=3.055 $Y=0.945 $X2=3.27
+ $Y2=1.335
cc_330 N_A_27_115#_M1015_g N_Y_c_577_n 0.00245758f $X=3.485 $Y=0.945 $X2=3.27
+ $Y2=1.335
cc_331 N_A_27_115#_M1014_g N_Y_c_580_n 0.00251111f $X=3.055 $Y=0.945 $X2=3.27
+ $Y2=2.215
cc_332 N_A_27_115#_c_328_n N_Y_c_580_n 0.0108556f $X=3.055 $Y=2.55 $X2=3.27
+ $Y2=2.215
cc_333 N_A_27_115#_c_329_n N_Y_c_580_n 0.0177725f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=2.215
cc_334 N_A_27_115#_M1015_g N_Y_c_580_n 0.00251111f $X=3.485 $Y=0.945 $X2=3.27
+ $Y2=2.215
cc_335 N_A_27_115#_c_356_n N_Y_c_581_n 0.0121767f $X=3.485 $Y=1.585 $X2=3.985
+ $Y2=2.33
cc_336 N_A_27_115#_c_357_n N_Y_c_581_n 0.0158479f $X=3.485 $Y=2.625 $X2=3.985
+ $Y2=2.33
cc_337 N_A_27_115#_c_328_n N_Y_c_582_n 0.00618817f $X=3.055 $Y=2.55 $X2=3.415
+ $Y2=2.33
cc_338 N_A_27_115#_c_329_n N_Y_c_582_n 0.00268861f $X=3.41 $Y=1.585 $X2=3.415
+ $Y2=2.33
cc_339 N_A_27_115#_c_330_n N_Y_c_582_n 0.00357274f $X=3.41 $Y=2.625 $X2=3.415
+ $Y2=2.33
cc_340 N_A_27_115#_M1016_g N_Y_c_583_n 0.00134358f $X=3.915 $Y=0.945 $X2=4.13
+ $Y2=1.335
cc_341 N_A_27_115#_M1017_g N_Y_c_583_n 0.00541892f $X=4.345 $Y=0.945 $X2=4.13
+ $Y2=1.335
cc_342 N_A_27_115#_M1016_g N_Y_c_586_n 0.00251111f $X=3.915 $Y=0.945 $X2=4.13
+ $Y2=2.215
cc_343 N_A_27_115#_c_342_n N_Y_c_586_n 0.0184054f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=2.215
cc_344 N_A_27_115#_M1017_g N_Y_c_586_n 0.00251111f $X=4.345 $Y=0.945 $X2=4.13
+ $Y2=2.215
cc_345 N_A_27_115#_c_358_n N_Y_c_586_n 0.00140336f $X=3.915 $Y=1.585 $X2=4.13
+ $Y2=2.215
cc_346 N_A_27_115#_c_359_n N_Y_c_586_n 0.00372651f $X=3.915 $Y=2.625 $X2=4.13
+ $Y2=2.215
cc_347 N_A_27_115#_c_335_n N_Y_c_587_n 0.00213861f $X=3.84 $Y=1.585 $X2=4.13
+ $Y2=1.22
cc_348 N_A_27_115#_M1016_g N_Y_c_587_n 0.0120182f $X=3.915 $Y=0.945 $X2=4.13
+ $Y2=1.22
