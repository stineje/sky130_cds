* File: sky130_osu_sc_18T_hs__dffr_l.spice
* Created: Thu Oct 29 17:07:33 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_hs__dffr_l.pex.spice"
.subckt sky130_osu_sc_18T_hs__dffr_l  GND VDD RN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* RN	RN
* VDD	VDD
* GND	GND
MM1015 N_A_110_115#_M1015_d N_RN_M1015_g N_GND_M1015_s N_GND_M1015_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1012 N_A_217_817#_M1012_d N_A_110_115#_M1012_g N_GND_M1012_s N_GND_M1015_b
+ NLOWVT L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1001 N_GND_M1001_d N_A_342_518#_M1001_g N_A_217_817#_M1012_d N_GND_M1015_b
+ NLOWVT L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 A_576_115# N_D_M1003_g N_GND_M1003_s N_GND_M1015_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1031 N_A_342_518#_M1031_d N_A_618_89#_M1031_g A_576_115# N_GND_M1015_b NLOWVT
+ L=0.15 W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1
+ R=6.66667 SA=75000.5 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1025 A_768_115# N_CK_M1025_g N_A_342_518#_M1031_d N_GND_M1015_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.1 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1028 N_GND_M1028_d N_A_217_817#_M1028_g A_768_115# N_GND_M1015_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.5
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1022 A_926_115# N_A_217_817#_M1022_g N_GND_M1028_d N_GND_M1015_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1013 N_A_998_115#_M1013_d N_CK_M1013_g A_926_115# N_GND_M1015_b NLOWVT L=0.15
+ W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1 R=6.66667
+ SA=75002.3 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1014 A_1118_115# N_A_618_89#_M1014_g N_A_998_115#_M1013_d N_GND_M1015_b NLOWVT
+ L=0.15 W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1
+ R=6.66667 SA=75002.9 SB=75001 A=0.15 P=2.3 MULT=1
MM1018 N_GND_M1018_d N_A_1160_89#_M1018_g A_1118_115# N_GND_M1015_b NLOWVT
+ L=0.15 W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667
+ SA=75003.3 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_618_89#_M1005_d N_CK_M1005_g N_GND_M1018_d N_GND_M1015_b NLOWVT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_1160_89#_M1006_d N_A_998_115#_M1006_g N_GND_M1006_s N_GND_M1015_b
+ NLOWVT L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_GND_M1007_d N_A_110_115#_M1007_g N_A_1160_89#_M1006_d N_GND_M1015_b
+ NLOWVT L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_GND_M1008_d N_A_1160_89#_M1008_g N_QN_M1008_s N_GND_M1015_b NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_Q_M1004_d N_QN_M1004_g N_GND_M1008_d N_GND_M1015_b NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_110_115#_M1011_d N_RN_M1011_g N_VDD_M1011_s N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1029 A_300_817# N_A_110_115#_M1029_g N_A_217_817#_M1029_s N_VDD_M1011_b PSHORT
+ L=0.15 W=2 AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.5 A=0.3 P=4.3 MULT=1
MM1021 N_VDD_M1021_d N_A_342_518#_M1021_g A_300_817# N_VDD_M1011_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.21 PD=4.53 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75000.5
+ SB=75000.2 A=0.3 P=4.3 MULT=1
MM1000 A_576_617# N_D_M1000_g N_VDD_M1000_s N_VDD_M1011_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.2
+ SB=75003.7 A=0.45 P=6.3 MULT=1
MM1030 N_A_342_518#_M1030_d N_CK_M1030_g A_576_617# N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75000.5 SB=75003.3 A=0.45 P=6.3 MULT=1
MM1023 A_768_617# N_A_618_89#_M1023_g N_A_342_518#_M1030_d N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75001.1 SB=75002.7 A=0.45 P=6.3 MULT=1
MM1026 N_VDD_M1026_d N_A_217_817#_M1026_g A_768_617# N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.5
+ SB=75002.4 A=0.45 P=6.3 MULT=1
MM1019 A_926_617# N_A_217_817#_M1019_g N_VDD_M1026_d N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75001.9
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1009 N_A_998_115#_M1009_d N_A_618_89#_M1009_g A_926_617# N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75002.3 SB=75001.6 A=0.45 P=6.3 MULT=1
MM1010 A_1118_617# N_CK_M1010_g N_A_998_115#_M1009_d N_VDD_M1011_b PSHORT L=0.15
+ W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75002.9 SB=75001 A=0.45 P=6.3 MULT=1
MM1016 N_VDD_M1016_d N_A_1160_89#_M1016_g A_1118_617# N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20
+ SA=75003.3 SB=75000.6 A=0.45 P=6.3 MULT=1
MM1002 N_A_618_89#_M1002_d N_CK_M1002_g N_VDD_M1016_d N_VDD_M1011_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.7
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1024 A_1466_817# N_A_998_115#_M1024_g N_A_1160_89#_M1024_s N_VDD_M1011_b
+ PSHORT L=0.15 W=2 AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1
+ R=13.3333 SA=75000.2 SB=75000.5 A=0.3 P=4.3 MULT=1
MM1017 N_VDD_M1017_d N_A_110_115#_M1017_g A_1466_817# N_VDD_M1011_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.21 PD=4.53 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333
+ SA=75000.5 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1027 N_VDD_M1027_d N_A_1160_89#_M1027_g N_QN_M1027_s N_VDD_M1011_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1020 N_Q_M1020_d N_QN_M1020_g N_VDD_M1027_d N_VDD_M1011_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX32_noxref N_GND_M1015_b N_VDD_M1011_b NWDIODE A=36.613 P=26.87
pX33_noxref noxref_24 RN RN PROBETYPE=1
pX34_noxref noxref_25 D D PROBETYPE=1
pX35_noxref noxref_26 CK CK PROBETYPE=1
pX36_noxref noxref_27 QN QN PROBETYPE=1
pX37_noxref noxref_28 Q Q PROBETYPE=1
c_1602 A_926_617# 0 1.57671e-19 $X=4.63 $Y=3.085
*
.include "sky130_osu_sc_18T_hs__dffr_l.pxi.spice"
*
.ends
*
*
