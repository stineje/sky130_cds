* File: sky130_osu_sc_18T_ms__inv_6.pxi.spice
* Created: Thu Oct 29 17:30:07 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__INV_6%GND N_GND_M1000_d N_GND_M1002_d N_GND_M1006_d
+ N_GND_M1010_d N_GND_M1000_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p N_GND_c_17_p
+ N_GND_c_23_p N_GND_c_36_p N_GND_c_30_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_MS__INV_6%GND
x_PM_SKY130_OSU_SC_18T_MS__INV_6%VDD N_VDD_M1001_d N_VDD_M1003_d N_VDD_M1007_d
+ N_VDD_M1011_d N_VDD_M1001_b N_VDD_c_84_p N_VDD_c_85_p N_VDD_c_90_p
+ N_VDD_c_96_p N_VDD_c_101_p N_VDD_c_111_p N_VDD_c_107_p VDD N_VDD_c_86_p
+ PM_SKY130_OSU_SC_18T_MS__INV_6%VDD
x_PM_SKY130_OSU_SC_18T_MS__INV_6%A N_A_c_141_n N_A_M1000_g N_A_c_145_n
+ N_A_c_194_n N_A_M1001_g N_A_c_146_n N_A_c_147_n N_A_c_148_n N_A_M1002_g
+ N_A_c_199_n N_A_M1003_g N_A_c_152_n N_A_c_154_n N_A_c_155_n N_A_M1004_g
+ N_A_c_205_n N_A_M1005_g N_A_c_159_n N_A_c_160_n N_A_c_161_n N_A_M1006_g
+ N_A_c_210_n N_A_M1007_g N_A_c_165_n N_A_c_167_n N_A_c_168_n N_A_M1008_g
+ N_A_c_172_n N_A_c_216_n N_A_M1009_g N_A_c_173_n N_A_c_174_n N_A_c_175_n
+ N_A_M1010_g N_A_c_221_n N_A_M1011_g N_A_c_179_n N_A_c_180_n N_A_c_181_n
+ N_A_c_182_n N_A_c_183_n N_A_c_184_n N_A_c_185_n N_A_c_186_n N_A_c_187_n
+ N_A_c_188_n N_A_c_189_n N_A_c_190_n N_A_c_191_n A N_A_c_192_n N_A_c_193_n
+ PM_SKY130_OSU_SC_18T_MS__INV_6%A
x_PM_SKY130_OSU_SC_18T_MS__INV_6%Y N_Y_M1000_s N_Y_M1004_s N_Y_M1008_s
+ N_Y_M1001_s N_Y_M1005_s N_Y_M1009_s N_Y_c_320_n N_Y_c_349_n Y N_Y_c_324_n
+ N_Y_c_350_n N_Y_c_326_n N_Y_c_327_n N_Y_c_329_n N_Y_c_352_n N_Y_c_354_n
+ N_Y_c_332_n N_Y_c_335_n N_Y_c_356_n N_Y_c_359_n N_Y_c_362_n N_Y_c_336_n
+ N_Y_c_340_n N_Y_c_345_n PM_SKY130_OSU_SC_18T_MS__INV_6%Y
cc_1 N_GND_M1000_b N_A_c_141_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.7
cc_2 N_GND_c_2_p N_A_c_141_n 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.7
cc_3 N_GND_c_3_p N_A_c_141_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.7
cc_4 N_GND_c_4_p N_A_c_141_n 0.00468827f $X=2.38 $Y=0.17 $X2=0.475 $Y2=1.7
cc_5 N_GND_M1000_b N_A_c_145_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.81
cc_6 N_GND_M1000_b N_A_c_146_n 0.01476f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.775
cc_7 N_GND_M1000_b N_A_c_147_n 0.00981662f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.885
cc_8 N_GND_M1000_b N_A_c_148_n 0.0166526f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.7
cc_9 N_GND_c_3_p N_A_c_148_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.7
cc_10 N_GND_c_10_p N_A_c_148_n 0.00356864f $X=1.12 $Y=0.825 $X2=0.905 $Y2=1.7
cc_11 N_GND_c_4_p N_A_c_148_n 0.00468827f $X=2.38 $Y=0.17 $X2=0.905 $Y2=1.7
cc_12 N_GND_M1000_b N_A_c_152_n 0.0213783f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.775
cc_13 N_GND_c_10_p N_A_c_152_n 0.00283047f $X=1.12 $Y=0.825 $X2=1.26 $Y2=1.775
cc_14 N_GND_M1000_b N_A_c_154_n 0.0173499f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.885
cc_15 N_GND_M1000_b N_A_c_155_n 0.0166526f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.7
cc_16 N_GND_c_10_p N_A_c_155_n 0.00356864f $X=1.12 $Y=0.825 $X2=1.335 $Y2=1.7
cc_17 N_GND_c_17_p N_A_c_155_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.335 $Y2=1.7
cc_18 N_GND_c_4_p N_A_c_155_n 0.00468827f $X=2.38 $Y=0.17 $X2=1.335 $Y2=1.7
cc_19 N_GND_M1000_b N_A_c_159_n 0.0195339f $X=-0.045 $Y=0 $X2=1.69 $Y2=1.775
cc_20 N_GND_M1000_b N_A_c_160_n 0.0145324f $X=-0.045 $Y=0 $X2=1.69 $Y2=2.885
cc_21 N_GND_M1000_b N_A_c_161_n 0.0166526f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.7
cc_22 N_GND_c_17_p N_A_c_161_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.765 $Y2=1.7
cc_23 N_GND_c_23_p N_A_c_161_n 0.00356864f $X=1.98 $Y=0.825 $X2=1.765 $Y2=1.7
cc_24 N_GND_c_4_p N_A_c_161_n 0.00468827f $X=2.38 $Y=0.17 $X2=1.765 $Y2=1.7
cc_25 N_GND_M1000_b N_A_c_165_n 0.0164591f $X=-0.045 $Y=0 $X2=2.12 $Y2=1.775
cc_26 N_GND_c_23_p N_A_c_165_n 0.00283047f $X=1.98 $Y=0.825 $X2=2.12 $Y2=1.775
cc_27 N_GND_M1000_b N_A_c_167_n 0.0124307f $X=-0.045 $Y=0 $X2=2.12 $Y2=2.885
cc_28 N_GND_M1000_b N_A_c_168_n 0.0166526f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.7
cc_29 N_GND_c_23_p N_A_c_168_n 0.00356864f $X=1.98 $Y=0.825 $X2=2.195 $Y2=1.7
cc_30 N_GND_c_30_p N_A_c_168_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.195 $Y2=1.7
cc_31 N_GND_c_4_p N_A_c_168_n 0.00468827f $X=2.38 $Y=0.17 $X2=2.195 $Y2=1.7
cc_32 N_GND_M1000_b N_A_c_172_n 0.0685082f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.81
cc_33 N_GND_M1000_b N_A_c_173_n 0.0385034f $X=-0.045 $Y=0 $X2=2.55 $Y2=1.775
cc_34 N_GND_M1000_b N_A_c_174_n 0.0295863f $X=-0.045 $Y=0 $X2=2.55 $Y2=2.885
cc_35 N_GND_M1000_b N_A_c_175_n 0.0208613f $X=-0.045 $Y=0 $X2=2.625 $Y2=1.7
cc_36 N_GND_c_36_p N_A_c_175_n 0.00713292f $X=2.84 $Y=0.825 $X2=2.625 $Y2=1.7
cc_37 N_GND_c_30_p N_A_c_175_n 0.00606474f $X=2.755 $Y=0.152 $X2=2.625 $Y2=1.7
cc_38 N_GND_c_4_p N_A_c_175_n 0.00468827f $X=2.38 $Y=0.17 $X2=2.625 $Y2=1.7
cc_39 N_GND_M1000_b N_A_c_179_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.775
cc_40 N_GND_M1000_b N_A_c_180_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.885
cc_41 N_GND_M1000_b N_A_c_181_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.775
cc_42 N_GND_M1000_b N_A_c_182_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.885
cc_43 N_GND_M1000_b N_A_c_183_n 0.0106787f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.775
cc_44 N_GND_M1000_b N_A_c_184_n 0.00980309f $X=-0.045 $Y=0 $X2=1.335 $Y2=2.885
cc_45 N_GND_M1000_b N_A_c_185_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.775
cc_46 N_GND_M1000_b N_A_c_186_n 0.00980309f $X=-0.045 $Y=0 $X2=1.765 $Y2=2.885
cc_47 N_GND_M1000_b N_A_c_187_n 0.0023879f $X=-0.045 $Y=0 $X2=2.195 $Y2=1.775
cc_48 N_GND_M1000_b N_A_c_188_n 0.00151234f $X=-0.045 $Y=0 $X2=2.195 $Y2=2.885
cc_49 N_GND_M1000_b N_A_c_189_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.305
cc_50 N_GND_M1000_b N_A_c_190_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_51 N_GND_M1000_b N_A_c_191_n 0.0382476f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_52 N_GND_M1000_b N_A_c_192_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.33
cc_53 N_GND_M1000_b N_A_c_193_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.14
cc_54 N_GND_M1000_b N_Y_c_320_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.595
cc_55 N_GND_c_2_p N_Y_c_320_n 0.00134236f $X=0.26 $Y=0.825 $X2=0.69 $Y2=1.595
cc_56 N_GND_c_10_p N_Y_c_320_n 7.53951e-19 $X=1.12 $Y=0.825 $X2=0.69 $Y2=1.595
cc_57 N_GND_M1000_b Y 0.0456345f $X=-0.045 $Y=0 $X2=0.76 $Y2=2.2
cc_58 N_GND_M1002_d N_Y_c_324_n 0.0127699f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1.48
cc_59 N_GND_c_10_p N_Y_c_324_n 0.0142303f $X=1.12 $Y=0.825 $X2=1.405 $Y2=1.48
cc_60 N_GND_M1000_b N_Y_c_326_n 0.0591815f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.845
cc_61 N_GND_M1006_d N_Y_c_327_n 0.0127699f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.48
cc_62 N_GND_c_23_p N_Y_c_327_n 0.0142303f $X=1.98 $Y=0.825 $X2=2.265 $Y2=1.48
cc_63 N_GND_M1000_b N_Y_c_329_n 0.00409378f $X=-0.045 $Y=0 $X2=1.695 $Y2=1.48
cc_64 N_GND_c_10_p N_Y_c_329_n 7.53951e-19 $X=1.12 $Y=0.825 $X2=1.695 $Y2=1.48
cc_65 N_GND_c_23_p N_Y_c_329_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=1.695 $Y2=1.48
cc_66 N_GND_M1000_b N_Y_c_332_n 0.00409378f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.595
cc_67 N_GND_c_23_p N_Y_c_332_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=1.595
cc_68 N_GND_c_36_p N_Y_c_332_n 0.00134236f $X=2.84 $Y=0.825 $X2=2.41 $Y2=1.595
cc_69 N_GND_M1000_b N_Y_c_335_n 0.0581802f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.845
cc_70 N_GND_M1000_b N_Y_c_336_n 0.00155118f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_71 N_GND_c_3_p N_Y_c_336_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.825
cc_72 N_GND_c_10_p N_Y_c_336_n 8.14297e-19 $X=1.12 $Y=0.825 $X2=0.69 $Y2=0.825
cc_73 N_GND_c_4_p N_Y_c_336_n 0.00475776f $X=2.38 $Y=0.17 $X2=0.69 $Y2=0.825
cc_74 N_GND_M1000_b N_Y_c_340_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_75 N_GND_c_10_p N_Y_c_340_n 8.14297e-19 $X=1.12 $Y=0.825 $X2=1.55 $Y2=0.825
cc_76 N_GND_c_17_p N_Y_c_340_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.825
cc_77 N_GND_c_23_p N_Y_c_340_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=0.825
cc_78 N_GND_c_4_p N_Y_c_340_n 0.00475776f $X=2.38 $Y=0.17 $X2=1.55 $Y2=0.825
cc_79 N_GND_M1000_b N_Y_c_345_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.825
cc_80 N_GND_c_23_p N_Y_c_345_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=0.825
cc_81 N_GND_c_30_p N_Y_c_345_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.825
cc_82 N_GND_c_4_p N_Y_c_345_n 0.00475776f $X=2.38 $Y=0.17 $X2=2.41 $Y2=0.825
cc_83 N_VDD_M1001_b N_A_c_194_n 0.0181616f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=2.96
cc_84 N_VDD_c_84_p N_A_c_194_n 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=2.96
cc_85 N_VDD_c_85_p N_A_c_194_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=2.96
cc_86 N_VDD_c_86_p N_A_c_194_n 0.00468827f $X=2.38 $Y=6.49 $X2=0.475 $Y2=2.96
cc_87 N_VDD_M1001_b N_A_c_147_n 0.00448664f $X=-0.045 $Y=2.905 $X2=0.83
+ $Y2=2.885
cc_88 N_VDD_M1001_b N_A_c_199_n 0.0159283f $X=-0.045 $Y=2.905 $X2=0.905 $Y2=2.96
cc_89 N_VDD_c_85_p N_A_c_199_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=2.96
cc_90 N_VDD_c_90_p N_A_c_199_n 0.00354579f $X=1.12 $Y=3.455 $X2=0.905 $Y2=2.96
cc_91 N_VDD_c_86_p N_A_c_199_n 0.00468827f $X=2.38 $Y=6.49 $X2=0.905 $Y2=2.96
cc_92 N_VDD_M1001_b N_A_c_154_n 0.00500158f $X=-0.045 $Y=2.905 $X2=1.26
+ $Y2=2.885
cc_93 N_VDD_c_90_p N_A_c_154_n 0.00341318f $X=1.12 $Y=3.455 $X2=1.26 $Y2=2.885
cc_94 N_VDD_M1001_b N_A_c_205_n 0.0159283f $X=-0.045 $Y=2.905 $X2=1.335 $Y2=2.96
cc_95 N_VDD_c_90_p N_A_c_205_n 0.00354579f $X=1.12 $Y=3.455 $X2=1.335 $Y2=2.96
cc_96 N_VDD_c_96_p N_A_c_205_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.335 $Y2=2.96
cc_97 N_VDD_c_86_p N_A_c_205_n 0.00468827f $X=2.38 $Y=6.49 $X2=1.335 $Y2=2.96
cc_98 N_VDD_M1001_b N_A_c_160_n 0.00448664f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.885
cc_99 N_VDD_M1001_b N_A_c_210_n 0.0159283f $X=-0.045 $Y=2.905 $X2=1.765 $Y2=2.96
cc_100 N_VDD_c_96_p N_A_c_210_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.765 $Y2=2.96
cc_101 N_VDD_c_101_p N_A_c_210_n 0.00354579f $X=1.98 $Y=3.455 $X2=1.765 $Y2=2.96
cc_102 N_VDD_c_86_p N_A_c_210_n 0.00468827f $X=2.38 $Y=6.49 $X2=1.765 $Y2=2.96
cc_103 N_VDD_M1001_b N_A_c_167_n 0.00500158f $X=-0.045 $Y=2.905 $X2=2.12
+ $Y2=2.885
cc_104 N_VDD_c_101_p N_A_c_167_n 0.00341318f $X=1.98 $Y=3.455 $X2=2.12 $Y2=2.885
cc_105 N_VDD_M1001_b N_A_c_216_n 0.0159283f $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.96
cc_106 N_VDD_c_101_p N_A_c_216_n 0.00354579f $X=1.98 $Y=3.455 $X2=2.195 $Y2=2.96
cc_107 N_VDD_c_107_p N_A_c_216_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.195
+ $Y2=2.96
cc_108 N_VDD_c_86_p N_A_c_216_n 0.00468827f $X=2.38 $Y=6.49 $X2=2.195 $Y2=2.96
cc_109 N_VDD_M1001_b N_A_c_174_n 0.00840215f $X=-0.045 $Y=2.905 $X2=2.55
+ $Y2=2.885
cc_110 N_VDD_M1001_b N_A_c_221_n 0.0204783f $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=2.96
cc_111 N_VDD_c_111_p N_A_c_221_n 0.00713292f $X=2.84 $Y=3.455 $X2=2.625 $Y2=2.96
cc_112 N_VDD_c_107_p N_A_c_221_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.625
+ $Y2=2.96
cc_113 N_VDD_c_86_p N_A_c_221_n 0.00468827f $X=2.38 $Y=6.49 $X2=2.625 $Y2=2.96
cc_114 N_VDD_M1001_b N_A_c_180_n 0.00244521f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.885
cc_115 N_VDD_M1001_b N_A_c_182_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=2.885
cc_116 N_VDD_M1001_b N_A_c_184_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.885
cc_117 N_VDD_M1001_b N_A_c_186_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.885
cc_118 N_VDD_M1001_b N_A_c_188_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.885
cc_119 N_VDD_M1001_d A 0.0162774f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.325
cc_120 N_VDD_c_84_p A 0.00522047f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.325
cc_121 N_VDD_c_90_p A 9.09141e-19 $X=1.12 $Y=3.455 $X2=0.32 $Y2=3.325
cc_122 N_VDD_M1001_d N_A_c_192_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_123 N_VDD_M1001_b N_A_c_192_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.32
+ $Y2=3.33
cc_124 N_VDD_c_84_p N_A_c_192_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_125 N_VDD_M1001_b N_Y_c_349_n 0.00248543f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.845
cc_126 N_VDD_M1001_b N_Y_c_350_n 0.00520877f $X=-0.045 $Y=2.905 $X2=1.405
+ $Y2=2.96
cc_127 N_VDD_c_90_p N_Y_c_350_n 0.0090257f $X=1.12 $Y=3.455 $X2=1.405 $Y2=2.96
cc_128 N_VDD_M1001_b N_Y_c_352_n 0.00520877f $X=-0.045 $Y=2.905 $X2=2.265
+ $Y2=2.96
cc_129 N_VDD_c_101_p N_Y_c_352_n 0.0090257f $X=1.98 $Y=3.455 $X2=2.265 $Y2=2.96
cc_130 N_VDD_M1001_b N_Y_c_354_n 0.00409378f $X=-0.045 $Y=2.905 $X2=1.695
+ $Y2=2.96
cc_131 N_VDD_M1001_b N_Y_c_335_n 0.00409378f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.845
cc_132 N_VDD_M1001_b N_Y_c_356_n 0.00361433f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.96
cc_133 N_VDD_c_85_p N_Y_c_356_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69 $Y2=2.96
cc_134 N_VDD_c_86_p N_Y_c_356_n 0.00475776f $X=2.38 $Y=6.49 $X2=0.69 $Y2=2.96
cc_135 N_VDD_M1001_b N_Y_c_359_n 0.00465961f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=2.96
cc_136 N_VDD_c_96_p N_Y_c_359_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55 $Y2=2.96
cc_137 N_VDD_c_86_p N_Y_c_359_n 0.00475776f $X=2.38 $Y=6.49 $X2=1.55 $Y2=2.96
cc_138 N_VDD_M1001_b N_Y_c_362_n 0.00465961f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.96
cc_139 N_VDD_c_107_p N_Y_c_362_n 0.00734006f $X=2.755 $Y=6.507 $X2=2.41 $Y2=2.96
cc_140 N_VDD_c_86_p N_Y_c_362_n 0.00475776f $X=2.38 $Y=6.49 $X2=2.41 $Y2=2.96
cc_141 A N_Y_M1001_s 0.00251573f $X=0.32 $Y=3.325 $X2=0.55 $Y2=3.085
cc_142 N_A_c_141_n N_Y_c_320_n 0.00942005f $X=0.475 $Y=1.7 $X2=0.69 $Y2=1.595
cc_143 N_A_c_148_n N_Y_c_320_n 0.00259753f $X=0.905 $Y=1.7 $X2=0.69 $Y2=1.595
cc_144 N_A_c_191_n N_Y_c_320_n 0.0011424f $X=0.535 $Y=2.305 $X2=0.69 $Y2=1.595
cc_145 N_A_c_194_n N_Y_c_349_n 0.00169643f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.845
cc_146 N_A_c_147_n N_Y_c_349_n 0.00270155f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.845
cc_147 N_A_c_199_n N_Y_c_349_n 0.00144225f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.845
cc_148 N_A_c_180_n N_Y_c_349_n 0.00102602f $X=0.475 $Y=2.885 $X2=0.69 $Y2=2.845
cc_149 N_A_c_182_n N_Y_c_349_n 0.00150284f $X=0.905 $Y=2.885 $X2=0.69 $Y2=2.845
cc_150 N_A_c_190_n N_Y_c_349_n 0.00173027f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.845
cc_151 N_A_c_191_n N_Y_c_349_n 8.31386e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.845
cc_152 A N_Y_c_349_n 0.00815006f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.845
cc_153 N_A_c_192_n N_Y_c_349_n 0.0071561f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.845
cc_154 N_A_c_141_n Y 0.00150089f $X=0.475 $Y=1.7 $X2=0.76 $Y2=2.2
cc_155 N_A_c_145_n Y 0.00792324f $X=0.475 $Y=2.81 $X2=0.76 $Y2=2.2
cc_156 N_A_c_146_n Y 0.0161013f $X=0.83 $Y=1.775 $X2=0.76 $Y2=2.2
cc_157 N_A_c_147_n Y 0.00363305f $X=0.83 $Y=2.885 $X2=0.76 $Y2=2.2
cc_158 N_A_c_148_n Y 0.00150089f $X=0.905 $Y=1.7 $X2=0.76 $Y2=2.2
cc_159 N_A_c_190_n Y 0.0178517f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_160 N_A_c_191_n Y 0.00668675f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_161 N_A_c_192_n Y 0.0182346f $X=0.32 $Y=3.33 $X2=0.76 $Y2=2.2
cc_162 N_A_c_193_n Y 0.00675469f $X=0.535 $Y=2.14 $X2=0.76 $Y2=2.2
cc_163 N_A_c_148_n N_Y_c_324_n 0.0129682f $X=0.905 $Y=1.7 $X2=1.405 $Y2=1.48
cc_164 N_A_c_152_n N_Y_c_324_n 0.0022289f $X=1.26 $Y=1.775 $X2=1.405 $Y2=1.48
cc_165 N_A_c_155_n N_Y_c_324_n 0.0129682f $X=1.335 $Y=1.7 $X2=1.405 $Y2=1.48
cc_166 N_A_c_199_n N_Y_c_350_n 0.00693713f $X=0.905 $Y=2.96 $X2=1.405 $Y2=2.96
cc_167 N_A_c_154_n N_Y_c_350_n 0.0120397f $X=1.26 $Y=2.885 $X2=1.405 $Y2=2.96
cc_168 N_A_c_205_n N_Y_c_350_n 0.00693713f $X=1.335 $Y=2.96 $X2=1.405 $Y2=2.96
cc_169 N_A_c_182_n N_Y_c_350_n 0.00560085f $X=0.905 $Y=2.885 $X2=1.405 $Y2=2.96
cc_170 N_A_c_184_n N_Y_c_350_n 0.00560085f $X=1.335 $Y=2.885 $X2=1.405 $Y2=2.96
cc_171 N_A_c_155_n N_Y_c_326_n 0.00150089f $X=1.335 $Y=1.7 $X2=1.55 $Y2=2.845
cc_172 N_A_c_159_n N_Y_c_326_n 0.0177499f $X=1.69 $Y=1.775 $X2=1.55 $Y2=2.845
cc_173 N_A_c_160_n N_Y_c_326_n 0.00562481f $X=1.69 $Y=2.885 $X2=1.55 $Y2=2.845
cc_174 N_A_c_161_n N_Y_c_326_n 0.00150089f $X=1.765 $Y=1.7 $X2=1.55 $Y2=2.845
cc_175 N_A_c_172_n N_Y_c_326_n 0.0141566f $X=2.195 $Y=2.81 $X2=1.55 $Y2=2.845
cc_176 N_A_c_161_n N_Y_c_327_n 0.0129682f $X=1.765 $Y=1.7 $X2=2.265 $Y2=1.48
cc_177 N_A_c_165_n N_Y_c_327_n 0.0022289f $X=2.12 $Y=1.775 $X2=2.265 $Y2=1.48
cc_178 N_A_c_168_n N_Y_c_327_n 0.0136594f $X=2.195 $Y=1.7 $X2=2.265 $Y2=1.48
cc_179 N_A_c_155_n N_Y_c_329_n 0.00259753f $X=1.335 $Y=1.7 $X2=1.695 $Y2=1.48
cc_180 N_A_c_161_n N_Y_c_329_n 0.00259753f $X=1.765 $Y=1.7 $X2=1.695 $Y2=1.48
cc_181 N_A_c_210_n N_Y_c_352_n 0.00693713f $X=1.765 $Y=2.96 $X2=2.265 $Y2=2.96
cc_182 N_A_c_167_n N_Y_c_352_n 0.0125508f $X=2.12 $Y=2.885 $X2=2.265 $Y2=2.96
cc_183 N_A_c_216_n N_Y_c_352_n 0.00693713f $X=2.195 $Y=2.96 $X2=2.265 $Y2=2.96
cc_184 N_A_c_186_n N_Y_c_352_n 0.00560085f $X=1.765 $Y=2.885 $X2=2.265 $Y2=2.96
cc_185 N_A_c_188_n N_Y_c_352_n 0.00642784f $X=2.195 $Y=2.885 $X2=2.265 $Y2=2.96
cc_186 N_A_c_205_n N_Y_c_354_n 0.00144225f $X=1.335 $Y=2.96 $X2=1.695 $Y2=2.96
cc_187 N_A_c_160_n N_Y_c_354_n 0.00397642f $X=1.69 $Y=2.885 $X2=1.695 $Y2=2.96
cc_188 N_A_c_210_n N_Y_c_354_n 0.00144225f $X=1.765 $Y=2.96 $X2=1.695 $Y2=2.96
cc_189 N_A_c_184_n N_Y_c_354_n 0.00150284f $X=1.335 $Y=2.885 $X2=1.695 $Y2=2.96
cc_190 N_A_c_186_n N_Y_c_354_n 0.00150284f $X=1.765 $Y=2.885 $X2=1.695 $Y2=2.96
cc_191 N_A_c_168_n N_Y_c_332_n 0.00262362f $X=2.195 $Y=1.7 $X2=2.41 $Y2=1.595
cc_192 N_A_c_175_n N_Y_c_332_n 0.00939395f $X=2.625 $Y=1.7 $X2=2.41 $Y2=1.595
cc_193 N_A_c_168_n N_Y_c_335_n 0.00150089f $X=2.195 $Y=1.7 $X2=2.41 $Y2=2.845
cc_194 N_A_c_172_n N_Y_c_335_n 0.0182294f $X=2.195 $Y=2.81 $X2=2.41 $Y2=2.845
cc_195 N_A_c_216_n N_Y_c_335_n 0.00144225f $X=2.195 $Y=2.96 $X2=2.41 $Y2=2.845
cc_196 N_A_c_173_n N_Y_c_335_n 0.0169795f $X=2.55 $Y=1.775 $X2=2.41 $Y2=2.845
cc_197 N_A_c_174_n N_Y_c_335_n 0.0141541f $X=2.55 $Y=2.885 $X2=2.41 $Y2=2.845
cc_198 N_A_c_175_n N_Y_c_335_n 0.00150089f $X=2.625 $Y=1.7 $X2=2.41 $Y2=2.845
cc_199 N_A_c_221_n N_Y_c_335_n 0.00541616f $X=2.625 $Y=2.96 $X2=2.41 $Y2=2.845
cc_200 N_A_c_188_n N_Y_c_335_n 0.00153387f $X=2.195 $Y=2.885 $X2=2.41 $Y2=2.845
cc_201 N_A_c_194_n N_Y_c_356_n 0.00199065f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.96
cc_202 N_A_c_147_n N_Y_c_356_n 0.00899372f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.96
cc_203 N_A_c_199_n N_Y_c_356_n 0.0035213f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.96
cc_204 N_A_c_190_n N_Y_c_356_n 0.00165526f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_205 N_A_c_191_n N_Y_c_356_n 5.06602e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_206 A N_Y_c_356_n 0.00938699f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.96
cc_207 N_A_c_192_n N_Y_c_356_n 0.0226156f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_208 N_A_c_205_n N_Y_c_359_n 0.0035213f $X=1.335 $Y=2.96 $X2=1.55 $Y2=2.96
cc_209 N_A_c_160_n N_Y_c_359_n 0.0108863f $X=1.69 $Y=2.885 $X2=1.55 $Y2=2.96
cc_210 N_A_c_210_n N_Y_c_359_n 0.0035213f $X=1.765 $Y=2.96 $X2=1.55 $Y2=2.96
cc_211 N_A_c_216_n N_Y_c_362_n 0.0035213f $X=2.195 $Y=2.96 $X2=2.41 $Y2=2.96
cc_212 N_A_c_174_n N_Y_c_362_n 0.0105836f $X=2.55 $Y=2.885 $X2=2.41 $Y2=2.96
cc_213 N_A_c_221_n N_Y_c_362_n 0.0035213f $X=2.625 $Y=2.96 $X2=2.41 $Y2=2.96
cc_214 N_A_c_141_n N_Y_c_336_n 0.00231637f $X=0.475 $Y=1.7 $X2=0.69 $Y2=0.825
cc_215 N_A_c_146_n N_Y_c_336_n 0.00256118f $X=0.83 $Y=1.775 $X2=0.69 $Y2=0.825
cc_216 N_A_c_148_n N_Y_c_336_n 0.00231637f $X=0.905 $Y=1.7 $X2=0.69 $Y2=0.825
cc_217 N_A_c_190_n N_Y_c_336_n 0.00110256f $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_218 N_A_c_191_n N_Y_c_336_n 3.64468e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_219 N_A_c_155_n N_Y_c_340_n 0.00231637f $X=1.335 $Y=1.7 $X2=1.55 $Y2=0.825
cc_220 N_A_c_159_n N_Y_c_340_n 0.00317228f $X=1.69 $Y=1.775 $X2=1.55 $Y2=0.825
cc_221 N_A_c_161_n N_Y_c_340_n 0.00231637f $X=1.765 $Y=1.7 $X2=1.55 $Y2=0.825
cc_222 N_A_c_168_n N_Y_c_345_n 0.00231637f $X=2.195 $Y=1.7 $X2=2.41 $Y2=0.825
cc_223 N_A_c_173_n N_Y_c_345_n 0.00317228f $X=2.55 $Y=1.775 $X2=2.41 $Y2=0.825
cc_224 N_A_c_175_n N_Y_c_345_n 0.00231637f $X=2.625 $Y=1.7 $X2=2.41 $Y2=0.825
