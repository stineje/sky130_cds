* File: sky130_osu_sc_12T_ms__dffsr_l.pex.spice
* Created: Fri Nov 12 15:23:21 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%GND 1 2 3 4 5 6 7 8 9 127 131 133 140
+ 142 152 154 158 160 170 172 182 184 191 193 203 205 212 238 240
c265 191 0 1.63226e-19 $X=7.47 $Y=0.755
c266 182 0 3.34232e-19 $X=6.52 $Y=0.755
c267 158 0 3.07651e-19 $X=3.02 $Y=0.755
c268 152 0 2.98797e-19 $X=2.5 $Y=0.755
c269 127 0 1.91032e-19 $X=-0.05 $Y=0
r270 238 240 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.855 $Y2=0.152
r271 214 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=0.152
+ $X2=9.71 $Y2=0.152
r272 210 234 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.152
r273 210 212 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.755
r274 206 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.152
+ $X2=8.75 $Y2=0.152
r275 205 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=0.152
+ $X2=9.71 $Y2=0.152
r276 201 233 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.152
r277 201 203 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.74
r278 194 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.152
+ $X2=7.47 $Y2=0.152
r279 193 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.152
+ $X2=8.75 $Y2=0.152
r280 189 232 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.152
r281 189 191 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.755
r282 184 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=0.152
+ $X2=7.47 $Y2=0.152
r283 180 182 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.52 $Y=0.305
+ $X2=6.52 $Y2=0.755
r284 173 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.152
+ $X2=4.77 $Y2=0.152
r285 168 228 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.152
r286 168 170 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.74
r287 160 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.152
+ $X2=4.77 $Y2=0.152
r288 156 158 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.02 $Y=0.305
+ $X2=3.02 $Y2=0.755
r289 155 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.152
+ $X2=2.5 $Y2=0.152
r290 154 155 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=2.935 $Y=0.152
+ $X2=2.585 $Y2=0.152
r291 150 224 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.152
r292 150 152 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.755
r293 143 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0.152
+ $X2=1.22 $Y2=0.152
r294 142 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.152
+ $X2=2.5 $Y2=0.152
r295 138 223 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.152
r296 138 140 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.74
r297 133 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.152
+ $X2=1.22 $Y2=0.152
r298 129 131 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r299 127 240 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=0.19
+ $X2=9.855 $Y2=0.19
r300 127 238 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r301 127 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.52 $Y2=0.305
r302 127 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.435 $Y2=0.152
r303 127 185 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.605 $Y2=0.152
r304 127 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.02 $Y2=0.305
r305 127 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=2.935 $Y2=0.152
r306 127 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.105 $Y2=0.152
r307 127 129 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r308 127 134 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r309 127 214 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.855 $Y=0.152
+ $X2=9.795 $Y2=0.152
r310 127 205 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=9.625 $Y2=0.152
r311 127 206 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.835 $Y2=0.152
r312 127 193 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.665 $Y2=0.152
r313 127 194 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=7.815 $Y=0.152
+ $X2=7.555 $Y2=0.152
r314 127 184 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.385 $Y2=0.152
r315 127 185 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.605 $Y2=0.152
r316 127 172 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.435 $Y2=0.152
r317 127 173 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.855 $Y2=0.152
r318 127 160 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=4.685 $Y2=0.152
r319 127 161 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.105 $Y2=0.152
r320 127 142 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.415 $Y2=0.152
r321 127 143 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.305 $Y2=0.152
r322 127 133 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.135 $Y2=0.152
r323 127 134 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r324 9 212 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.57
+ $Y=0.575 $X2=9.71 $Y2=0.755
r325 8 203 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.61
+ $Y=0.575 $X2=8.75 $Y2=0.74
r326 7 191 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.755
r327 6 182 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.755
r328 5 170 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.575 $X2=4.77 $Y2=0.74
r329 4 158 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.575 $X2=3.02 $Y2=0.755
r330 3 152 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.575 $X2=2.5 $Y2=0.755
r331 2 140 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.575 $X2=1.22 $Y2=0.74
r332 1 131 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%VDD 1 2 3 4 5 6 7 89 93 95 103 105 111
+ 113 121 123 131 133 139 141 149 153 168 172
r166 168 172 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=4.287
+ $X2=9.855 $Y2=4.287
r167 156 168 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=4.25
+ $X2=0.335 $Y2=4.25
r168 153 172 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=4.25
+ $X2=9.855 $Y2=4.25
r169 151 166 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=4.287
+ $X2=9.71 $Y2=4.287
r170 151 153 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.795 $Y=4.287
+ $X2=9.855 $Y2=4.287
r171 147 166 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.71 $Y=4.135
+ $X2=9.71 $Y2=4.287
r172 147 149 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=9.71 $Y=4.135
+ $X2=9.71 $Y2=3.265
r173 144 146 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=8.495 $Y=4.287
+ $X2=9.175 $Y2=4.287
r174 142 165 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=4.287
+ $X2=7.9 $Y2=4.287
r175 142 144 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=7.985 $Y=4.287
+ $X2=8.495 $Y2=4.287
r176 141 166 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=4.287
+ $X2=9.71 $Y2=4.287
r177 141 146 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.625 $Y=4.287
+ $X2=9.175 $Y2=4.287
r178 137 165 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=4.287
r179 137 139 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=3.7
r180 134 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=4.287
+ $X2=6.52 $Y2=4.287
r181 134 136 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=6.605 $Y=4.287
+ $X2=7.135 $Y2=4.287
r182 133 165 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=4.287
+ $X2=7.9 $Y2=4.287
r183 133 136 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=4.287
+ $X2=7.135 $Y2=4.287
r184 129 163 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.52 $Y=4.135
+ $X2=6.52 $Y2=4.287
r185 129 131 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.52 $Y=4.135
+ $X2=6.52 $Y2=3.21
r186 126 128 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=4.287
+ $X2=5.775 $Y2=4.287
r187 124 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=4.287
+ $X2=4.77 $Y2=4.287
r188 124 126 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=4.855 $Y=4.287
+ $X2=5.095 $Y2=4.287
r189 123 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=4.287
+ $X2=6.52 $Y2=4.287
r190 123 128 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=6.435 $Y=4.287
+ $X2=5.775 $Y2=4.287
r191 119 161 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.77 $Y=4.135
+ $X2=4.77 $Y2=4.287
r192 119 121 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.77 $Y=4.135
+ $X2=4.77 $Y2=3.295
r193 116 118 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=4.287
+ $X2=4.415 $Y2=4.287
r194 114 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=4.287
+ $X2=3.02 $Y2=4.287
r195 114 116 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.105 $Y=4.287
+ $X2=3.735 $Y2=4.287
r196 113 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=4.287
+ $X2=4.77 $Y2=4.287
r197 113 118 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.685 $Y=4.287
+ $X2=4.415 $Y2=4.287
r198 109 160 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.02 $Y=4.135
+ $X2=3.02 $Y2=4.287
r199 109 111 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.02 $Y=4.135
+ $X2=3.02 $Y2=3.295
r200 106 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=4.287
+ $X2=2.07 $Y2=4.287
r201 106 108 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.155 $Y=4.287
+ $X2=2.375 $Y2=4.287
r202 105 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=4.287
+ $X2=3.02 $Y2=4.287
r203 105 108 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=2.935 $Y=4.287
+ $X2=2.375 $Y2=4.287
r204 101 158 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.07 $Y=4.135
+ $X2=2.07 $Y2=4.287
r205 101 103 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=4.135
+ $X2=2.07 $Y2=3.7
r206 98 100 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=4.287
+ $X2=1.695 $Y2=4.287
r207 96 156 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r208 96 98 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.015 $Y2=4.287
r209 95 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=4.287
+ $X2=2.07 $Y2=4.287
r210 95 100 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.985 $Y=4.287
+ $X2=1.695 $Y2=4.287
r211 91 156 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r212 91 93 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r213 89 153 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=9.65 $Y=4.135 $X2=9.855 $Y2=4.22
r214 89 146 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=4.135 $X2=9.175 $Y2=4.22
r215 89 144 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=4.135 $X2=8.495 $Y2=4.22
r216 89 165 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=4.135 $X2=7.815 $Y2=4.22
r217 89 136 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=4.135 $X2=7.135 $Y2=4.22
r218 89 163 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=4.135 $X2=6.455 $Y2=4.22
r219 89 128 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=4.135 $X2=5.775 $Y2=4.22
r220 89 126 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=4.135 $X2=5.095 $Y2=4.22
r221 89 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=4.135 $X2=4.415 $Y2=4.22
r222 89 116 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=4.135 $X2=3.735 $Y2=4.22
r223 89 160 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=4.135 $X2=3.055 $Y2=4.22
r224 89 108 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=4.135 $X2=2.375 $Y2=4.22
r225 89 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=4.135 $X2=1.695 $Y2=4.22
r226 89 98 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=4.135 $X2=1.015 $Y2=4.22
r227 89 156 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=4.135 $X2=0.335 $Y2=4.22
r228 7 149 300 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=2 $X=9.57
+ $Y=3.025 $X2=9.71 $Y2=3.265
r229 6 139 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.605 $X2=7.9 $Y2=3.7
r230 5 131 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=3.21
r231 4 121 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=4.63
+ $Y=2.605 $X2=4.77 $Y2=3.295
r232 3 111 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.605 $X2=3.02 $Y2=3.295
r233 2 103 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.605 $X2=2.07 $Y2=3.7
r234 1 93 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%RN 3 5 7 13 15 21
c42 21 0 7.48684e-20 $X=0.325 $Y=2.85
c43 3 0 1.41286e-20 $X=0.475 $Y=0.835
r44 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=2.85
+ $X2=0.325 $Y2=2.85
r45 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.53 $Y2=1.825
r46 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r47 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=1.99
+ $X2=0.32 $Y2=1.825
r48 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=1.99 $X2=0.32
+ $Y2=2.85
r49 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.825 $X2=0.53 $Y2=1.825
r50 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.53 $Y2=1.825
r51 5 7 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=3.235
r52 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.53 $Y2=1.825
r53 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_110_115# 1 3 10 13 15 17 18 20 23 26
+ 29 33 36 39 43 47 54 57 62 65 68 72 73 74 78 81 82
c228 78 0 5.45583e-20 $X=0.87 $Y=1.37
c229 72 0 1.41286e-20 $X=0.87 $Y=1.255
c230 68 0 1.57074e-19 $X=8.86 $Y=1.21
c231 65 0 7.48684e-20 $X=0.87 $Y=2.26
c232 54 0 1.68724e-19 $X=0.87 $Y=1.37
c233 39 0 1.09867e-19 $X=8.545 $Y=2.27
r234 81 82 0.0806629 $w=2.95e-07 $l=1.15e-07 $layer=MET1_cond $X=8.862 $Y=1.37
+ $X2=8.862 $Y2=1.255
r235 75 82 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=8.86 $Y=1.085
+ $X2=8.86 $Y2=1.255
r236 73 75 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=8.775 $Y=1
+ $X2=8.86 $Y2=1.085
r237 73 74 7.52974 $w=1.7e-07 $l=7.82e-06 $layer=MET1_cond $X=8.775 $Y=1
+ $X2=0.955 $Y2=1
r238 72 78 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.87 $Y=1.255
+ $X2=0.87 $Y2=1.37
r239 71 74 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.87 $Y=1.085
+ $X2=0.955 $Y2=1
r240 71 72 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=0.87 $Y=1.085
+ $X2=0.87 $Y2=1.255
r241 70 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.86 $Y=1.37
+ $X2=8.86 $Y2=1.37
r242 68 70 7.74603 $w=2.52e-07 $l=1.6e-07 $layer=LI1_cond $X=8.86 $Y=1.21
+ $X2=8.86 $Y2=1.37
r243 63 65 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.26
+ $X2=0.87 $Y2=2.26
r244 61 62 14.2597 $w=1.73e-07 $l=2.25e-07 $layer=LI1_cond $X=0.87 $Y=1.207
+ $X2=1.095 $Y2=1.207
r245 59 61 11.4078 $w=1.73e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.207
+ $X2=0.87 $Y2=1.207
r246 57 62 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.23 $Y=1.21
+ $X2=1.095 $Y2=1.21
r247 54 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.87 $Y=1.37
+ $X2=0.87 $Y2=1.37
r248 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=2.26
r249 52 54 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=1.37
r250 51 61 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.207
r251 51 54 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.37
r252 47 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r253 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.26
r254 45 47 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.955
r255 41 59 0.89264 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=0.69 $Y=1.12
+ $X2=0.69 $Y2=1.207
r256 41 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=1.12
+ $X2=0.69 $Y2=0.755
r257 39 40 60.25 $w=2.04e-07 $l=2.55e-07 $layer=POLY_cond $X=8.545 $Y=2.27
+ $X2=8.8 $Y2=2.27
r258 38 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.86
+ $Y=1.21 $X2=8.86 $Y2=1.21
r259 36 38 12.05 $w=2.4e-07 $l=6e-08 $layer=POLY_cond $X=8.8 $Y=1.21 $X2=8.86
+ $Y2=1.21
r260 32 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.21 $X2=1.23 $Y2=1.21
r261 32 33 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.23 $Y=1.21 $X2=1.29
+ $Y2=1.21
r262 27 29 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.29 $Y=2.34
+ $X2=1.425 $Y2=2.34
r263 26 40 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.8 $Y=2.125
+ $X2=8.8 $Y2=2.27
r264 25 36 13.7767 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=1.375
+ $X2=8.8 $Y2=1.21
r265 25 26 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=8.8 $Y=1.375
+ $X2=8.8 $Y2=2.125
r266 21 39 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.545 $Y=2.415
+ $X2=8.545 $Y2=2.27
r267 21 23 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.545 $Y=2.415
+ $X2=8.545 $Y2=3.235
r268 18 36 53.2208 $w=2.4e-07 $l=3.37565e-07 $layer=POLY_cond $X=8.535 $Y=1.045
+ $X2=8.8 $Y2=1.21
r269 18 20 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.535 $Y=1.045
+ $X2=8.535 $Y2=0.755
r270 15 33 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.435 $Y=1.045
+ $X2=1.29 $Y2=1.21
r271 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.435 $Y=1.045
+ $X2=1.435 $Y2=0.755
r272 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=2.415
+ $X2=1.425 $Y2=2.34
r273 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.425 $Y=2.415
+ $X2=1.425 $Y2=3.235
r274 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=2.265
+ $X2=1.29 $Y2=2.34
r275 9 33 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.375
+ $X2=1.29 $Y2=1.21
r276 9 10 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.29 $Y=1.375
+ $X2=1.29 $Y2=2.265
r277 3 49 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r278 3 47 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r279 1 43 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%SN 1 2 5 9 13 17 22 25 29 32 34 37 39
+ 45 47 48 49 56
c192 48 0 1.36413e-19 $X=7.79 $Y=2.85
c193 29 0 1.5152e-19 $X=1.71 $Y=2.62
r194 54 56 0.00223214 $w=2.8e-07 $l=5e-09 $layer=MET1_cond $X=7.935 $Y=2.802
+ $X2=7.94 $Y2=2.802
r195 49 51 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=2.195 $Y=2.85
+ $X2=2.055 $Y2=2.85
r196 48 54 0.0838839 $w=2.8e-07 $l=1.67287e-07 $layer=MET1_cond $X=7.79 $Y=2.85
+ $X2=7.935 $Y2=2.802
r197 48 49 5.38733 $w=1.7e-07 $l=5.595e-06 $layer=MET1_cond $X=7.79 $Y=2.85
+ $X2=2.195 $Y2=2.85
r198 42 45 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.935 $Y=1.815
+ $X2=8.025 $Y2=1.815
r199 41 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.055 $Y=2.85
+ $X2=2.055 $Y2=2.85
r200 39 41 17.9872 $w=2.34e-07 $l=3.45e-07 $layer=LI1_cond $X=1.71 $Y=2.777
+ $X2=2.055 $Y2=2.777
r201 34 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.935 $Y=2.845
+ $X2=7.935 $Y2=2.845
r202 32 47 5.51377 $w=1.73e-07 $l=8.7e-08 $layer=LI1_cond $X=7.937 $Y=2.482
+ $X2=7.937 $Y2=2.395
r203 32 34 23.0057 $w=1.73e-07 $l=3.63e-07 $layer=LI1_cond $X=7.937 $Y=2.482
+ $X2=7.937 $Y2=2.845
r204 30 42 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=1.94
+ $X2=7.935 $Y2=1.815
r205 30 47 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=7.935 $Y=1.94
+ $X2=7.935 $Y2=2.395
r206 29 39 2.60974 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.71 $Y=2.62
+ $X2=1.71 $Y2=2.777
r207 28 37 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.975
+ $X2=1.71 $Y2=1.89
r208 28 29 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.71 $Y=1.975
+ $X2=1.71 $Y2=2.62
r209 25 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.025
+ $Y=1.775 $X2=8.025 $Y2=1.775
r210 25 27 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=1.775
+ $X2=8.035 $Y2=1.94
r211 25 26 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=1.775
+ $X2=8.035 $Y2=1.61
r212 22 23 5.53115 $w=3.05e-07 $l=3.5e-08 $layer=POLY_cond $X=1.855 $Y=1.89
+ $X2=1.89 $Y2=1.89
r213 21 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.89 $X2=1.71 $Y2=1.89
r214 21 22 22.9148 $w=3.05e-07 $l=1.45e-07 $layer=POLY_cond $X=1.71 $Y=1.89
+ $X2=1.855 $Y2=1.89
r215 17 27 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=8.115 $Y=3.235
+ $X2=8.115 $Y2=1.94
r216 13 26 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=8.045 $Y=0.835
+ $X2=8.045 $Y2=1.61
r217 9 19 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.925 $Y=0.835
+ $X2=1.925 $Y2=1.295
r218 3 22 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=2.055
+ $X2=1.855 $Y2=1.89
r219 3 5 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.855 $Y=2.055
+ $X2=1.855 $Y2=3.235
r220 2 23 10.4756 $w=2.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.725
+ $X2=1.89 $Y2=1.89
r221 1 19 38.6248 $w=2.2e-07 $l=1.1e-07 $layer=POLY_cond $X=1.89 $Y=1.405
+ $X2=1.89 $Y2=1.295
r222 1 2 93.3405 $w=2.2e-07 $l=3.2e-07 $layer=POLY_cond $X=1.89 $Y=1.405
+ $X2=1.89 $Y2=1.725
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_432_424# 1 3 11 15 18 22 23 24 25 28
+ 29 30 32 35 41
c109 41 0 1.72079e-19 $X=3.795 $Y=0.755
c110 30 0 1.07085e-19 $X=2.855 $Y=2.705
c111 23 0 1.29912e-19 $X=3.71 $Y=1.285
c112 11 0 1.32807e-19 $X=2.285 $Y=0.835
r113 41 43 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=3.795 $Y=0.755
+ $X2=3.895 $Y2=0.755
r114 35 37 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=3.895 $Y=2.955
+ $X2=3.895 $Y2=3.635
r115 33 35 2.03372 $w=3.38e-07 $l=6e-08 $layer=LI1_cond $X=3.895 $Y=2.895
+ $X2=3.895 $Y2=2.955
r116 31 41 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.795 $Y=0.935
+ $X2=3.795 $Y2=0.755
r117 31 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.795 $Y=0.935
+ $X2=3.795 $Y2=1.2
r118 29 33 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=3.725 $Y=2.705
+ $X2=3.895 $Y2=2.895
r119 29 30 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.725 $Y=2.705
+ $X2=2.855 $Y2=2.705
r120 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=2.62
+ $X2=2.855 $Y2=2.705
r121 27 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.77 $Y=2.37
+ $X2=2.77 $Y2=2.62
r122 26 40 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.38 $Y=2.285
+ $X2=2.295 $Y2=2.325
r123 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.685 $Y=2.285
+ $X2=2.77 $Y2=2.37
r124 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.685 $Y=2.285
+ $X2=2.38 $Y2=2.285
r125 23 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=1.285
+ $X2=3.795 $Y2=1.2
r126 23 24 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.71 $Y=1.285
+ $X2=2.38 $Y2=1.285
r127 22 40 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=2.2
+ $X2=2.295 $Y2=2.325
r128 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=1.37
+ $X2=2.38 $Y2=1.285
r129 21 22 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.295 $Y=1.37
+ $X2=2.295 $Y2=2.2
r130 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=2.285 $X2=2.295 $Y2=2.285
r131 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.285
+ $X2=2.295 $Y2=2.45
r132 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.285
+ $X2=2.295 $Y2=2.12
r133 15 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.285 $Y=3.235
+ $X2=2.285 $Y2=2.45
r134 11 19 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=2.285 $Y=0.835
+ $X2=2.285 $Y2=2.12
r135 3 37 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.605 $X2=3.895 $Y2=3.635
r136 3 35 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.605 $X2=3.895 $Y2=2.955
r137 1 43 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.575 $X2=3.895 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%D 3 7 10 14 19
c38 19 0 1.41836e-19 $X=3.295 $Y=1.74
c39 10 0 1.12321e-19 $X=3.295 $Y=1.74
c40 7 0 1.07085e-19 $X=3.235 $Y=3.235
r41 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.295 $Y=1.74
+ $X2=3.295 $Y2=1.74
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.74 $X2=3.295 $Y2=1.74
r43 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.74
+ $X2=3.295 $Y2=1.905
r44 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.74
+ $X2=3.295 $Y2=1.575
r45 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.235 $Y=3.235
+ $X2=3.235 $Y2=1.905
r46 3 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.235 $Y=0.835
+ $X2=3.235 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c254 76 0 1.37846e-19 $X=6.735 $Y=2.11
c255 74 0 8.87231e-20 $X=5.74 $Y=2.11
c256 55 0 6.79641e-20 $X=5.49 $Y=2.11
c257 48 0 1.98654e-19 $X=4.135 $Y=1.37
c258 44 0 1.86602e-19 $X=4.05 $Y=2.11
c259 37 0 4.76307e-20 $X=5.885 $Y=2.285
c260 30 0 1.29912e-19 $X=4.135 $Y=1.205
c261 25 0 1.41836e-19 $X=3.655 $Y=2.285
r262 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.03 $Y=2.11
+ $X2=5.885 $Y2=2.11
r263 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.735 $Y=2.11
+ $X2=6.88 $Y2=2.11
r264 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.735 $Y=2.11
+ $X2=6.03 $Y2=2.11
r265 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.8 $Y=2.11
+ $X2=3.655 $Y2=2.11
r266 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.74 $Y=2.11
+ $X2=5.885 $Y2=2.11
r267 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.74 $Y=2.11
+ $X2=3.8 $Y2=2.11
r268 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=2.11
+ $X2=5.885 $Y2=2.11
r269 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.885 $Y=2.11
+ $X2=5.885 $Y2=2.285
r270 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.655 $Y=2.11
+ $X2=3.655 $Y2=2.11
r271 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.655 $Y=2.11
+ $X2=3.655 $Y2=2.285
r272 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.88 $Y=2.11
+ $X2=6.88 $Y2=2.11
r273 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.88 $Y=2.11
+ $X2=6.88 $Y2=2.285
r274 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.11
+ $X2=5.885 $Y2=2.11
r275 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.8 $Y=2.11
+ $X2=5.49 $Y2=2.11
r276 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.405 $Y=2.025
+ $X2=5.49 $Y2=2.11
r277 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.405 $Y=2.025
+ $X2=5.405 $Y2=1.37
r278 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.135 $Y=2.025
+ $X2=4.135 $Y2=1.37
r279 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=2.11
+ $X2=3.655 $Y2=2.11
r280 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.05 $Y=2.11
+ $X2=4.135 $Y2=2.025
r281 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.05 $Y=2.11
+ $X2=3.74 $Y2=2.11
r282 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=2.285 $X2=6.88 $Y2=2.285
r283 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.762 $Y=1.205
+ $X2=6.762 $Y2=1.355
r284 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=2.285 $X2=5.885 $Y2=2.285
r285 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=2.285
+ $X2=5.885 $Y2=2.45
r286 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.37 $X2=5.405 $Y2=1.37
r287 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.37
+ $X2=5.405 $Y2=1.205
r288 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.37 $X2=4.135 $Y2=1.37
r289 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.37
+ $X2=4.135 $Y2=1.205
r290 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=2.285 $X2=3.655 $Y2=2.285
r291 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=2.285
+ $X2=3.655 $Y2=2.45
r292 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.79 $Y=2.12
+ $X2=6.837 $Y2=2.285
r293 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.79 $Y=2.12
+ $X2=6.79 $Y2=1.355
r294 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.735 $Y=2.45
+ $X2=6.837 $Y2=2.285
r295 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.735 $Y=2.45
+ $X2=6.735 $Y2=3.235
r296 17 40 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.735 $Y=0.835
+ $X2=6.735 $Y2=1.205
r297 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.945 $Y=3.235
+ $X2=5.945 $Y2=2.45
r298 10 34 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.345 $Y=0.835
+ $X2=5.345 $Y2=1.205
r299 7 30 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.195 $Y=0.835
+ $X2=4.195 $Y2=1.205
r300 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.595 $Y=3.235
+ $X2=3.595 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_217_521# 1 3 11 15 17 18 21 22 27 31
+ 35 37 38 41 47 52 53 54 59
c161 54 0 1.32807e-19 $X=1.855 $Y=1.37
c162 53 0 2.71143e-19 $X=4.49 $Y=1.37
c163 47 0 1.5821e-19 $X=4.725 $Y=2.285
c164 41 0 1.63226e-19 $X=1.71 $Y=0.755
c165 37 0 2.23283e-19 $X=1.565 $Y=1.55
c166 31 0 6.36774e-20 $X=4.985 $Y=3.235
c167 22 0 1.86602e-19 $X=4.63 $Y=2.285
c168 21 0 6.79641e-20 $X=4.91 $Y=2.285
c169 15 0 6.36774e-20 $X=4.555 $Y=3.235
r170 54 56 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.37
+ $X2=1.71 $Y2=1.37
r171 53 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.49 $Y=1.37
+ $X2=4.635 $Y2=1.37
r172 53 54 2.53719 $w=1.7e-07 $l=2.635e-06 $layer=MET1_cond $X=4.49 $Y=1.37
+ $X2=1.855 $Y2=1.37
r173 50 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.37
+ $X2=4.635 $Y2=1.37
r174 50 52 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=4.635 $Y=1.33
+ $X2=4.725 $Y2=1.33
r175 45 52 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.725 $Y=1.455
+ $X2=4.725 $Y2=1.33
r176 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.725 $Y=1.455
+ $X2=4.725 $Y2=2.285
r177 44 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.37
+ $X2=1.71 $Y2=1.37
r178 41 44 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.71 $Y=0.755
+ $X2=1.71 $Y2=1.37
r179 39 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.455
+ $X2=1.71 $Y2=1.37
r180 37 39 6.81649 $w=1.7e-07 $l=1.86548e-07 $layer=LI1_cond $X=1.565 $Y=1.55
+ $X2=1.71 $Y2=1.455
r181 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.565 $Y=1.55
+ $X2=1.295 $Y2=1.55
r182 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.635
+ $X2=1.295 $Y2=1.55
r183 33 35 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=1.21 $Y=1.635
+ $X2=1.21 $Y2=3.295
r184 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.985 $Y=2.42
+ $X2=4.985 $Y2=3.235
r185 25 27 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.985 $Y=1.235
+ $X2=4.985 $Y2=0.835
r186 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=2.285 $X2=4.725 $Y2=2.285
r187 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=2.285
+ $X2=4.725 $Y2=2.285
r188 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=2.285
+ $X2=4.985 $Y2=2.42
r189 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=2.285
+ $X2=4.725 $Y2=2.285
r190 20 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=1.37 $X2=4.725 $Y2=1.37
r191 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=1.37
+ $X2=4.725 $Y2=1.37
r192 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=1.37
+ $X2=4.985 $Y2=1.235
r193 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=1.37
+ $X2=4.725 $Y2=1.37
r194 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.63 $Y2=2.285
r195 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.555 $Y2=3.235
r196 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.235
+ $X2=4.63 $Y2=1.37
r197 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.555 $Y=1.235
+ $X2=4.555 $Y2=0.835
r198 3 35 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.605 $X2=1.21 $Y2=3.295
r199 1 41 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.575 $X2=1.71 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_704_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 50 54 59 63 67 69 70 75
c209 70 0 4.76307e-20 $X=6.05 $Y=1.725
c210 59 0 1.36413e-19 $X=7.22 $Y=2.62
c211 44 0 2.26569e-19 $X=5.885 $Y=1.725
c212 34 0 1.98654e-19 $X=3.715 $Y=1.28
c213 18 0 1.12321e-19 $X=4.195 $Y=3.235
r214 70 72 0.116207 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=6.05 $Y=1.725
+ $X2=5.885 $Y2=1.725
r215 69 75 0.0841272 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=6.835 $Y=1.725
+ $X2=6.95 $Y2=1.725
r216 69 70 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=6.835 $Y=1.725
+ $X2=6.05 $Y2=1.725
r217 65 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=2.705
+ $X2=7.22 $Y2=2.705
r218 62 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.95 $Y=1.725
+ $X2=6.95 $Y2=1.725
r219 62 63 16.1867 $w=1.83e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=1.717
+ $X2=7.22 $Y2=1.717
r220 59 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.62
+ $X2=7.22 $Y2=2.705
r221 58 63 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=7.22 $Y=1.81
+ $X2=7.22 $Y2=1.717
r222 58 59 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=7.22 $Y=1.81
+ $X2=7.22 $Y2=2.62
r223 54 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.95 $Y=2.955
+ $X2=6.95 $Y2=3.635
r224 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=2.79
+ $X2=6.95 $Y2=2.705
r225 52 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=2.79
+ $X2=6.95 $Y2=2.955
r226 48 62 1.22693 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=6.95 $Y=1.625
+ $X2=6.95 $Y2=1.717
r227 48 50 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.95 $Y=1.625
+ $X2=6.95 $Y2=0.755
r228 44 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=1.725
+ $X2=5.885 $Y2=1.725
r229 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=1.725 $X2=5.885 $Y2=1.725
r230 39 41 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=5.885 $Y=1.725
+ $X2=5.885 $Y2=1.82
r231 39 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.725
+ $X2=5.885 $Y2=1.56
r232 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.595 $Y=1.28
+ $X2=3.715 $Y2=1.28
r233 30 40 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=5.945 $Y=0.835
+ $X2=5.945 $Y2=1.56
r234 27 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=1.82
+ $X2=5.345 $Y2=1.82
r235 26 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.75 $Y=1.82
+ $X2=5.885 $Y2=1.82
r236 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.75 $Y=1.82
+ $X2=5.42 $Y2=1.82
r237 22 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.345 $Y=1.895
+ $X2=5.345 $Y2=1.82
r238 22 24 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=5.345 $Y=1.895
+ $X2=5.345 $Y2=3.235
r239 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=1.82
+ $X2=4.195 $Y2=1.82
r240 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=1.82
+ $X2=5.345 $Y2=1.82
r241 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.27 $Y=1.82 $X2=4.27
+ $Y2=1.82
r242 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=1.895
+ $X2=4.195 $Y2=1.82
r243 16 18 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=4.195 $Y=1.895
+ $X2=4.195 $Y2=3.235
r244 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=1.82
+ $X2=4.195 $Y2=1.82
r245 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.12 $Y=1.82
+ $X2=3.79 $Y2=1.82
r246 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=1.745
+ $X2=3.79 $Y2=1.82
r247 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.715 $Y=1.355
+ $X2=3.715 $Y2=1.28
r248 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.715 $Y=1.355
+ $X2=3.715 $Y2=1.745
r249 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.205
+ $X2=3.595 $Y2=1.28
r250 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.595 $Y=1.205
+ $X2=3.595 $Y2=0.835
r251 3 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=2.605 $X2=6.95 $Y2=3.635
r252 3 54 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=2.605 $X2=6.95 $Y2=2.955
r253 1 50 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.575 $X2=6.95 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_1246_89# 1 3 11 15 23 27 30 34 35 38
+ 39 40 42 49 53 55 57 62 65 66 67 71 73
c213 49 0 1.63226e-19 $X=8.26 $Y=0.755
c214 42 0 1.6261e-19 $X=6.365 $Y=1.71
c215 39 0 8.77106e-20 $X=9.47 $Y=2.375
c216 35 0 1.57074e-19 $X=9.382 $Y=1.545
c217 34 0 2.20654e-19 $X=9.38 $Y=1.71
c218 11 0 1.35097e-19 $X=6.305 $Y=0.835
r219 69 71 0.105038 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=6.365 $Y=2.48
+ $X2=6.515 $Y2=2.48
r220 66 73 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.235 $Y=1.71
+ $X2=9.38 $Y2=1.71
r221 66 67 1.79096 $w=1.7e-07 $l=1.86e-06 $layer=MET1_cond $X=9.235 $Y=1.71
+ $X2=7.375 $Y2=1.71
r222 64 67 0.0706952 $w=1.7e-07 $l=1.14782e-07 $layer=MET1_cond $X=7.305
+ $Y=1.795 $X2=7.375 $Y2=1.71
r223 64 65 0.736385 $w=1.4e-07 $l=5.95e-07 $layer=MET1_cond $X=7.305 $Y=1.795
+ $X2=7.305 $Y2=2.39
r224 62 65 0.0709685 $w=1.75e-07 $l=1.80222e-07 $layer=MET1_cond $X=7.165
+ $Y=2.482 $X2=7.305 $Y2=2.39
r225 62 71 0.588306 $w=1.75e-07 $l=6.5e-07 $layer=MET1_cond $X=7.165 $Y=2.482
+ $X2=6.515 $Y2=2.482
r226 57 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.38 $Y=1.71
+ $X2=9.38 $Y2=1.71
r227 55 57 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.845 $Y=1.71
+ $X2=9.38 $Y2=1.71
r228 51 55 5.37722 $w=2.41e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=1.795
+ $X2=8.845 $Y2=1.71
r229 51 53 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=8.76 $Y=1.795
+ $X2=8.76 $Y2=3.295
r230 47 51 25.3112 $w=2.41e-07 $l=6.89202e-07 $layer=LI1_cond $X=8.26 $Y=1.345
+ $X2=8.76 $Y2=1.795
r231 47 49 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.26 $Y=1.345
+ $X2=8.26 $Y2=0.755
r232 45 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.365 $Y=2.48
+ $X2=6.365 $Y2=2.48
r233 42 45 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.365 $Y=1.71
+ $X2=6.365 $Y2=2.48
r234 39 40 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=2.375
+ $X2=9.47 $Y2=2.525
r235 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=1.17 $X2=9.47
+ $Y2=1.32
r236 36 39 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.445 $Y=1.875
+ $X2=9.445 $Y2=2.375
r237 35 38 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.445 $Y=1.545
+ $X2=9.445 $Y2=1.32
r238 34 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.38
+ $Y=1.71 $X2=9.38 $Y2=1.71
r239 34 36 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=1.71
+ $X2=9.382 $Y2=1.875
r240 34 35 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=1.71
+ $X2=9.382 $Y2=1.545
r241 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=1.71 $X2=6.365 $Y2=1.71
r242 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.71
+ $X2=6.365 $Y2=1.875
r243 30 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.71
+ $X2=6.365 $Y2=1.545
r244 27 40 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=9.495 $Y=3.445
+ $X2=9.495 $Y2=2.525
r245 23 37 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=9.495 $Y=0.755
+ $X2=9.495 $Y2=1.17
r246 15 32 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=6.305 $Y=3.235
+ $X2=6.305 $Y2=1.875
r247 11 31 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.305 $Y=0.835
+ $X2=6.305 $Y2=1.545
r248 3 53 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=8.62
+ $Y=2.605 $X2=8.76 $Y2=3.295
r249 1 49 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=8.12
+ $Y=0.575 $X2=8.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_1084_115# 1 3 10 11 13 16 20 26 30 32
+ 33 36 40 43 49 52 53 54 55 62
c174 55 0 1.35097e-19 $X=5.89 $Y=1.37
c175 53 0 1.5821e-19 $X=5.21 $Y=1.37
c176 49 0 1.71621e-19 $X=5.645 $Y=0.755
c177 30 0 1.57671e-19 $X=5.065 $Y=1.37
c178 16 0 6.36774e-20 $X=7.685 $Y=3.235
r179 55 60 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=5.89 $Y=1.37
+ $X2=5.745 $Y2=1.34
r180 54 62 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=1.37
+ $X2=7.595 $Y2=1.37
r181 54 55 1.5021 $w=1.7e-07 $l=1.56e-06 $layer=MET1_cond $X=7.45 $Y=1.37
+ $X2=5.89 $Y2=1.37
r182 53 57 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.21 $Y=1.37
+ $X2=5.065 $Y2=1.37
r183 52 60 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=5.6 $Y=1.37
+ $X2=5.745 $Y2=1.34
r184 52 53 0.375524 $w=1.7e-07 $l=3.9e-07 $layer=MET1_cond $X=5.6 $Y=1.37
+ $X2=5.21 $Y2=1.37
r185 49 51 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=5.652 $Y=0.755
+ $X2=5.652 $Y2=1.035
r186 43 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=1.37
+ $X2=7.595 $Y2=1.37
r187 43 46 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.595 $Y=1.37
+ $X2=7.595 $Y2=2.285
r188 40 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=1.34
r189 40 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=1.035
r190 34 36 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=5.645 $Y=2.79
+ $X2=5.645 $Y2=3.295
r191 32 34 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=2.705
+ $X2=5.645 $Y2=2.79
r192 32 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=2.705
+ $X2=5.15 $Y2=2.705
r193 30 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.065 $Y=1.37
+ $X2=5.065 $Y2=1.37
r194 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=2.62
+ $X2=5.15 $Y2=2.705
r195 28 30 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.065 $Y=2.62
+ $X2=5.065 $Y2=1.37
r196 25 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=2.285 $X2=7.595 $Y2=2.285
r197 25 26 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=2.285
+ $X2=7.685 $Y2=2.285
r198 22 25 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=2.285
+ $X2=7.595 $Y2=2.285
r199 18 20 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=7.505 $Y=1.29
+ $X2=7.685 $Y2=1.29
r200 14 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.685 $Y=2.42
+ $X2=7.685 $Y2=2.285
r201 14 16 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=7.685 $Y=2.42
+ $X2=7.685 $Y2=3.235
r202 11 20 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.685 $Y=1.21
+ $X2=7.685 $Y2=1.29
r203 11 13 120.5 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=7.685 $Y=1.21
+ $X2=7.685 $Y2=0.835
r204 10 22 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.505 $Y=2.15
+ $X2=7.505 $Y2=2.285
r205 9 18 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.505 $Y=1.37
+ $X2=7.505 $Y2=1.29
r206 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.505 $Y=1.37
+ $X2=7.505 $Y2=2.15
r207 3 36 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=5.42
+ $Y=2.605 $X2=5.645 $Y2=3.295
r208 1 49 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=5.42
+ $Y=0.575 $X2=5.645 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c90 42 0 8.77106e-20 $X=9.285 $Y=2.48
c91 33 0 9.99996e-20 $X=9.78 $Y=2.285
c92 31 0 1.20654e-19 $X=9.78 $Y=1.37
c93 27 0 1.09867e-19 $X=9.28 $Y=2.48
r94 40 42 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=9.28 $Y=2.48
+ $X2=9.285 $Y2=2.48
r95 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.865 $Y=2.2
+ $X2=9.865 $Y2=1.915
r96 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.865 $Y=1.455
+ $X2=9.865 $Y2=1.915
r97 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=2.285
+ $X2=9.865 $Y2=2.2
r98 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=2.285
+ $X2=9.365 $Y2=2.285
r99 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.37
+ $X2=9.865 $Y2=1.455
r100 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=1.37
+ $X2=9.365 $Y2=1.37
r101 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=2.48
+ $X2=9.28 $Y2=2.48
r102 27 29 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=9.28 $Y=2.48
+ $X2=9.28 $Y2=3.265
r103 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=2.37
+ $X2=9.365 $Y2=2.285
r104 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.28 $Y=2.37
+ $X2=9.28 $Y2=2.48
r105 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=1.285
+ $X2=9.365 $Y2=1.37
r106 21 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.28 $Y=1.285
+ $X2=9.28 $Y2=0.755
r107 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.865
+ $Y=1.915 $X2=9.865 $Y2=1.915
r108 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=1.915
+ $X2=9.865 $Y2=2.08
r109 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=1.915
+ $X2=9.865 $Y2=1.75
r110 15 20 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=9.925 $Y=3.445
+ $X2=9.925 $Y2=2.08
r111 11 19 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=9.925 $Y=0.755
+ $X2=9.925 $Y2=1.75
r112 3 29 300 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=2 $X=9.155
+ $Y=3.025 $X2=9.28 $Y2=3.265
r113 1 23 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.575 $X2=9.28 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_300_521# 1 2 11 13 14 17
c20 1 0 1.5152e-19 $X=1.5 $Y=2.605
r21 15 17 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.5 $Y=3.275 $X2=2.5
+ $Y2=3.295
r22 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=3.19
+ $X2=2.5 $Y2=3.275
r23 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.415 $Y=3.19
+ $X2=1.725 $Y2=3.19
r24 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.275
+ $X2=1.725 $Y2=3.19
r25 9 11 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.64 $Y=3.275 $X2=1.64
+ $Y2=3.295
r26 2 17 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=2.605 $X2=2.5 $Y2=3.295
r27 1 11 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.605 $X2=1.64 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%A_1469_521# 1 2 11 13 14 17
r20 15 17 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.33 $Y=3.27
+ $X2=8.33 $Y2=3.295
r21 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.245 $Y=3.185
+ $X2=8.33 $Y2=3.27
r22 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.245 $Y=3.185
+ $X2=7.555 $Y2=3.185
r23 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=3.27
+ $X2=7.555 $Y2=3.185
r24 9 11 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.47 $Y=3.27 $X2=7.47
+ $Y2=3.295
r25 2 17 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=2.605 $X2=8.33 $Y2=3.295
r26 1 11 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=2.605 $X2=7.47 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFFSR_L%Q 1 3 10 13 20 22 26 28 31
r24 28 29 8.56905 $w=1.68e-07 $l=1.18e-07 $layer=LI1_cond $X=10.137 $Y=2.61
+ $X2=10.255 $Y2=2.61
r25 24 26 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=1.035
+ $X2=10.255 $Y2=1.035
r26 20 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.255 $Y=2.11
+ $X2=10.255 $Y2=2.11
r27 18 29 0.644183 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=2.525
+ $X2=10.255 $Y2=2.61
r28 18 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=10.255 $Y=2.525
+ $X2=10.255 $Y2=2.11
r29 17 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=1.12
+ $X2=10.255 $Y2=1.035
r30 17 20 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=10.255 $Y=1.12
+ $X2=10.255 $Y2=2.11
r31 11 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=0.95
+ $X2=10.14 $Y2=1.035
r32 11 13 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.14 $Y=0.95
+ $X2=10.14 $Y2=0.755
r33 10 22 1.39429 $w=1.73e-07 $l=2.2e-08 $layer=LI1_cond $X=10.137 $Y=3.243
+ $X2=10.137 $Y2=3.265
r34 9 28 0.502328 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.137 $Y=2.695
+ $X2=10.137 $Y2=2.61
r35 9 10 34.7304 $w=1.73e-07 $l=5.48e-07 $layer=LI1_cond $X=10.137 $Y=2.695
+ $X2=10.137 $Y2=3.243
r36 3 22 300 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=2 $X=10
+ $Y=3.025 $X2=10.14 $Y2=3.265
r37 1 13 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=10 $Y=0.575
+ $X2=10.14 $Y2=0.755
.ends

