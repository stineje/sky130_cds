* File: sky130_osu_sc_12T_ms__addh_l.pex.spice
* Created: Fri Nov 12 15:20:01 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%GND 1 2 45 47 55 57 70 86 88
r104 86 88 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r105 72 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r106 68 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r107 68 70 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.755
r108 58 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r109 57 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r110 53 81 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r111 53 55 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.755
r112 47 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r113 45 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r114 45 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r115 45 72 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r116 45 57 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r117 45 58 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r118 45 47 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r119 2 70 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.755
r120 1 55 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%VDD 1 2 3 37 39 46 50 56 58 66 72 80 84
r57 80 84 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=3.74 $Y2=4.287
r58 72 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=4.25
+ $X2=3.74 $Y2=4.25
r59 70 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=4.287
+ $X2=3.05 $Y2=4.287
r60 70 72 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=4.287
+ $X2=3.74 $Y2=4.287
r61 66 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.05 $Y=2.955
+ $X2=3.05 $Y2=3.635
r62 64 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=4.135
+ $X2=3.05 $Y2=4.287
r63 64 69 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.05 $Y=4.135 $X2=3.05
+ $Y2=3.635
r64 61 63 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=4.287
+ $X2=2.38 $Y2=4.287
r65 59 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=4.287
+ $X2=1.61 $Y2=4.287
r66 59 61 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=4.287
+ $X2=1.7 $Y2=4.287
r67 58 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=4.287
+ $X2=3.05 $Y2=4.287
r68 58 63 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=4.287
+ $X2=2.38 $Y2=4.287
r69 54 76 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=4.135
+ $X2=1.61 $Y2=4.287
r70 54 56 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.61 $Y=4.135
+ $X2=1.61 $Y2=3.295
r71 51 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=4.287
+ $X2=0.75 $Y2=4.287
r72 51 53 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=4.287
+ $X2=1.02 $Y2=4.287
r73 50 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=4.287
+ $X2=1.61 $Y2=4.287
r74 50 53 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=4.287
+ $X2=1.02 $Y2=4.287
r75 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.75 $Y=2.955
+ $X2=0.75 $Y2=3.635
r76 44 75 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=4.135
+ $X2=0.75 $Y2=4.287
r77 44 49 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.75 $Y=4.135 $X2=0.75
+ $Y2=3.635
r78 41 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r79 39 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=4.287
+ $X2=0.75 $Y2=4.287
r80 39 41 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=4.287
+ $X2=0.34 $Y2=4.287
r81 37 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r82 37 78 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r83 37 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r84 37 61 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r85 37 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r86 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r87 3 56 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.605 $X2=1.61 $Y2=3.295
r88 2 49 400 $w=1.7e-07 $l=6.97872e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.03 $X2=0.75 $Y2=3.635
r89 2 46 400 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.03 $X2=0.75 $Y2=2.955
r90 1 69 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=2.605 $X2=3.05 $Y2=3.635
r91 1 66 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=2.605 $X2=3.05 $Y2=2.955
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%CON 1 7 8 23 27 30 37 39 40 43 47 49 51
+ 54 56 57 61 67 68 73 76 81 82 87 90
c140 90 0 2.7119e-19 $X=3.42 $Y=1.37
c141 82 0 1.57622e-19 $X=0.78 $Y=1.37
c142 68 0 4.75316e-20 $X=2.99 $Y=0.635
c143 54 0 1.92558e-19 $X=3.42 $Y=1.285
r144 82 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.37
+ $X2=0.635 $Y2=1.37
r145 81 87 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.37
+ $X2=2.62 $Y2=1.37
r146 81 82 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.37
+ $X2=0.78 $Y2=1.37
r147 76 79 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.85 $Y=0.635
+ $X2=3.85 $Y2=0.755
r148 75 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.37
+ $X2=3.42 $Y2=1.37
r149 68 71 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.99 $Y=0.635
+ $X2=2.99 $Y2=0.755
r150 66 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.37
+ $X2=2.62 $Y2=1.37
r151 61 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.84 $Y=2.955
+ $X2=3.84 $Y2=3.635
r152 59 61 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.84 $Y=2.555
+ $X2=3.84 $Y2=2.955
r153 58 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=0.635
+ $X2=3.42 $Y2=0.635
r154 57 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.85 $Y2=0.635
r155 57 58 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.505 $Y2=0.635
r156 54 75 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.285
+ $X2=3.42 $Y2=1.37
r157 54 56 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.42 $Y=1.285
+ $X2=3.42 $Y2=0.755
r158 53 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.72
+ $X2=3.42 $Y2=0.635
r159 53 56 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.42 $Y=0.72
+ $X2=3.42 $Y2=0.755
r160 52 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.635
+ $X2=2.99 $Y2=0.635
r161 51 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.635
+ $X2=3.42 $Y2=0.635
r162 51 52 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.335 $Y=0.635
+ $X2=3.075 $Y2=0.635
r163 50 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.47
+ $X2=2.62 $Y2=2.47
r164 49 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.47
+ $X2=3.84 $Y2=2.555
r165 49 50 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.47
+ $X2=2.705 $Y2=2.47
r166 48 66 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.37
+ $X2=2.62 $Y2=1.37
r167 47 75 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.37
+ $X2=3.42 $Y2=1.37
r168 47 48 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.37
+ $X2=2.705 $Y2=1.37
r169 43 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.62 $Y=2.955
+ $X2=2.62 $Y2=3.635
r170 41 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.555
+ $X2=2.62 $Y2=2.47
r171 41 43 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.62 $Y=2.555
+ $X2=2.62 $Y2=2.955
r172 40 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.385
+ $X2=2.62 $Y2=2.47
r173 39 66 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.455
+ $X2=2.62 $Y2=1.37
r174 39 40 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.455
+ $X2=2.62 $Y2=2.385
r175 37 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.37
+ $X2=0.635 $Y2=1.37
r176 34 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.35 $Y=1.37
+ $X2=0.635 $Y2=1.37
r177 30 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.37 $X2=0.35 $Y2=1.37
r178 30 32 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.37
+ $X2=0.382 $Y2=1.535
r179 30 31 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.37
+ $X2=0.382 $Y2=1.205
r180 27 32 980.409 $w=1.5e-07 $l=1.912e-06 $layer=POLY_cond $X=0.475 $Y=3.447
+ $X2=0.475 $Y2=1.535
r181 23 31 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.475 $Y=0.755
+ $X2=0.475 $Y2=1.205
r182 8 63 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=2.605 $X2=3.84 $Y2=3.635
r183 8 61 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=2.605 $X2=3.84 $Y2=2.955
r184 7 45 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.605 $X2=2.62 $Y2=3.635
r185 7 43 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.605 $X2=2.62 $Y2=2.955
r186 1 79 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.755
r187 1 56 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=0.755
r188 1 71 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%B 3 7 11 15 18 22 25 30 39 42 44
c101 44 0 4.99902e-20 $X=3.21 $Y=1.74
c102 22 0 1.42567e-19 $X=3.205 $Y=1.74
c103 18 0 1.57622e-19 $X=0.905 $Y=1.74
c104 11 0 4.75316e-20 $X=3.205 $Y=0.835
r105 41 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=3.205 $Y=1.74
+ $X2=3.21 $Y2=1.74
r106 41 42 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.205 $Y=1.74
+ $X2=3.06 $Y2=1.74
r107 39 42 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=1.742
+ $X2=3.06 $Y2=1.742
r108 37 39 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=1.74
+ $X2=1.05 $Y2=1.74
r109 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=1.74
+ $X2=3.205 $Y2=1.74
r110 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=1.74
+ $X2=0.905 $Y2=1.74
r111 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.74 $X2=3.205 $Y2=1.74
r112 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.74
+ $X2=3.205 $Y2=1.905
r113 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.74 $X2=0.905 $Y2=1.74
r114 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.74
+ $X2=0.905 $Y2=1.905
r115 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.74
+ $X2=0.905 $Y2=1.575
r116 15 23 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.265 $Y=3.235
+ $X2=3.265 $Y2=1.905
r117 9 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.575
+ $X2=3.205 $Y2=1.74
r118 9 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.205 $Y=1.575
+ $X2=3.205 $Y2=0.835
r119 7 20 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.965 $Y=3.235
+ $X2=0.965 $Y2=1.905
r120 3 19 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.965 $Y=0.835
+ $X2=0.965 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%A 3 7 11 15 18 22 26 31 40 42 43
c88 22 0 1.74252e-19 $X=3.685 $Y=2.11
r89 42 43 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.11
+ $X2=3.54 $Y2=2.11
r90 40 43 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.107
+ $X2=3.54 $Y2=2.107
r91 38 40 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.11
+ $X2=1.53 $Y2=2.11
r92 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.11
+ $X2=3.685 $Y2=2.11
r93 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.11
+ $X2=1.385 $Y2=2.11
r94 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.11 $X2=3.685 $Y2=2.11
r95 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.11
+ $X2=3.685 $Y2=2.275
r96 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.11
+ $X2=3.685 $Y2=1.945
r97 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.11 $X2=1.385 $Y2=2.11
r98 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.11
+ $X2=1.385 $Y2=2.275
r99 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.11
+ $X2=1.385 $Y2=1.945
r100 15 23 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=3.635 $Y=0.835
+ $X2=3.635 $Y2=1.945
r101 11 24 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.625 $Y=3.235
+ $X2=3.625 $Y2=2.275
r102 7 20 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.395 $Y=3.235
+ $X2=1.395 $Y2=2.275
r103 3 19 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.325 $Y=0.835
+ $X2=1.325 $Y2=1.945
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%A_208_521# 1 3 10 13 15 17 21 23 27 31
+ 33 38 39 42 44 45 48 51 53
c113 31 0 2.52869e-20 $X=2.835 $Y=3.235
c114 23 0 9.69384e-20 $X=2.7 $Y=1.32
r115 53 55 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.475
+ $X2=1.825 $Y2=1.475
r116 52 53 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.475
+ $X2=1.725 $Y2=1.475
r117 50 53 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.64
+ $X2=1.725 $Y2=1.475
r118 50 51 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=1.64
+ $X2=1.725 $Y2=2.445
r119 46 52 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.31
+ $X2=1.54 $Y2=1.475
r120 46 48 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.54 $Y=1.31
+ $X2=1.54 $Y2=0.755
r121 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=2.53
+ $X2=1.725 $Y2=2.445
r122 44 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=2.53
+ $X2=1.265 $Y2=2.53
r123 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=2.615
+ $X2=1.265 $Y2=2.53
r124 40 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.18 $Y=2.615
+ $X2=1.18 $Y2=3.295
r125 36 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.475 $X2=1.825 $Y2=1.475
r126 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.475
+ $X2=1.825 $Y2=1.64
r127 33 36 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.32
+ $X2=1.825 $Y2=1.475
r128 29 31 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.835 $Y=2.265
+ $X2=2.835 $Y2=3.235
r129 25 27 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.775 $Y=1.245
+ $X2=2.775 $Y2=0.835
r130 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.32
+ $X2=2.285 $Y2=1.32
r131 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.32
+ $X2=2.775 $Y2=1.245
r132 23 24 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.32 $X2=2.36
+ $Y2=1.32
r133 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.245
+ $X2=2.285 $Y2=1.32
r134 19 21 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.285 $Y=1.245
+ $X2=2.285 $Y2=0.755
r135 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.19
+ $X2=1.885 $Y2=2.19
r136 17 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.19
+ $X2=2.835 $Y2=2.265
r137 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.19 $X2=1.96
+ $Y2=2.19
r138 16 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.32
+ $X2=1.825 $Y2=1.32
r139 15 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.32
+ $X2=2.285 $Y2=1.32
r140 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.32
+ $X2=1.96 $Y2=1.32
r141 11 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.265
+ $X2=1.885 $Y2=2.19
r142 11 13 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.885 $Y=2.265
+ $X2=1.885 $Y2=3.445
r143 10 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.115
+ $X2=1.885 $Y2=2.19
r144 10 37 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.115
+ $X2=1.885 $Y2=1.64
r145 3 42 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.605 $X2=1.18 $Y2=3.295
r146 1 48 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.4 $Y=0.575
+ $X2=1.54 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%S 1 3 10 16 24 27 30
r33 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=2.735
+ $X2=0.26 $Y2=2.85
r34 22 24 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=2.735
+ $X2=0.26 $Y2=1.905
r35 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.11
+ $X2=0.26 $Y2=0.995
r36 21 24 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.11
+ $X2=0.26 $Y2=1.905
r37 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.85
+ $X2=0.26 $Y2=2.85
r38 16 19 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.26 $Y=2.85
+ $X2=0.26 $Y2=3.275
r39 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=0.995
+ $X2=0.26 $Y2=0.995
r40 10 13 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=0.74
+ $X2=0.26 $Y2=0.995
r41 3 19 300 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.03 $X2=0.26 $Y2=3.275
r42 1 10 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__ADDH_L%CO 1 3 11 15 21 24 25 28
c54 24 0 2.52869e-20 $X=2.175 $Y=2.48
r55 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.48
+ $X2=2.175 $Y2=2.48
r56 24 26 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.48
+ $X2=2.137 $Y2=2.565
r57 24 25 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.48
+ $X2=2.137 $Y2=2.395
r58 19 21 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=0.992
+ $X2=2.175 $Y2=0.992
r59 17 21 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.175 $Y=1.08
+ $X2=2.175 $Y2=0.992
r60 17 25 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.08
+ $X2=2.175 $Y2=2.395
r61 15 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.1 $Y=3.275 $X2=2.1
+ $Y2=2.565
r62 9 19 0.89264 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.07 $Y=0.905 $X2=2.07
+ $Y2=0.992
r63 9 11 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0.905
+ $X2=2.07 $Y2=0.74
r64 3 15 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=3.025 $X2=2.1 $Y2=3.275
r65 1 11 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.74
.ends

