* File: sky130_osu_sc_12T_ms__nor2_1.pex.spice
* Created: Fri Nov 12 15:25:29 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_1%GND 1 2 21 25 27 35 41 44
r28 41 44 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r29 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r30 27 33 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.305
r31 23 25 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r32 21 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r33 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r34 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r35 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r36 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r37 2 35 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
r38 1 25 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_1%VDD 1 13 15 21 27 30
r18 27 30 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r19 24 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r20 19 24 4.25596 $w=1.7e-07 $l=2.13185e-07 $layer=LI1_cond $X=1.05 $Y=4.135
+ $X2=1.197 $Y2=4.287
r21 19 21 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.05 $Y=4.135 $X2=1.05
+ $Y2=3.635
r22 15 24 3.30228 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=0.965 $Y=4.287
+ $X2=1.197 $Y2=4.287
r23 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=4.287
+ $X2=0.34 $Y2=4.287
r24 13 24 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r25 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r26 1 21 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.605 $X2=1.05 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_1%B 3 7 10 13 19 22
r49 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.65 $Y=2.48
+ $X2=0.65 $Y2=2.48
r50 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.65 $Y=1.695
+ $X2=0.65 $Y2=2.48
r51 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=1.61
+ $X2=0.65 $Y2=1.695
r52 13 15 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.565 $Y=1.61
+ $X2=0.415 $Y2=1.61
r53 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.61 $X2=0.415 $Y2=1.61
r54 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.61
+ $X2=0.415 $Y2=1.775
r55 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.61
+ $X2=0.415 $Y2=1.445
r56 7 12 748.638 $w=1.5e-07 $l=1.46e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=1.775
r57 3 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.445
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_1%A 3 7 10 14 20
r36 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=2.85
+ $X2=0.99 $Y2=2.85
r37 14 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.99 $Y=2.275
+ $X2=0.99 $Y2=2.85
r38 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.275 $X2=0.99 $Y2=2.275
r39 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.275
+ $X2=0.942 $Y2=2.44
r40 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.275
+ $X2=0.942 $Y2=2.11
r41 7 11 653.777 $w=1.5e-07 $l=1.275e-06 $layer=POLY_cond $X=0.905 $Y=0.835
+ $X2=0.905 $Y2=2.11
r42 3 12 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.835 $Y=3.235
+ $X2=0.835 $Y2=2.44
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_1%Y 1 3 10 18 23 24 28 34
r42 26 28 0.519956 $w=1.7e-07 $l=5.4e-07 $layer=MET1_cond $X=0.69 $Y=2.025
+ $X2=0.69 $Y2=1.485
r43 25 34 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1
r44 25 28 0.356266 $w=1.7e-07 $l=3.7e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1.485
r45 24 31 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=2.11
+ $X2=0.26 $Y2=2.11
r46 23 26 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=2.11
+ $X2=0.69 $Y2=2.025
r47 23 24 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=2.11
+ $X2=0.405 $Y2=2.11
r48 21 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1 $X2=0.69
+ $Y2=1
r49 18 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0.755
+ $X2=0.69 $Y2=1
r50 13 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r51 10 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.11
+ $X2=0.26 $Y2=2.11
r52 10 13 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.26 $Y=2.11
+ $X2=0.26 $Y2=2.955
r53 3 15 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r54 3 13 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r55 1 18 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

