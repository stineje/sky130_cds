magic
tech sky130A
magscale 1 2
timestamp 1612373520
<< nwell >>
rect -9 529 286 1119
<< nmoslvt >>
rect 80 115 110 243
rect 152 115 182 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 115 152 243
rect 182 215 235 243
rect 182 131 193 215
rect 227 131 235 215
rect 182 115 235 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 949 166 965
rect 110 605 121 949
rect 155 605 166 949
rect 110 565 166 605
rect 196 949 249 965
rect 196 673 207 949
rect 241 673 249 949
rect 196 565 249 673
<< ndiffc >>
rect 35 131 69 215
rect 193 131 227 215
<< pdiffc >>
rect 35 741 69 949
rect 121 605 155 949
rect 207 673 241 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 80 518 110 565
rect 37 502 110 518
rect 37 468 47 502
rect 81 468 110 502
rect 37 452 110 468
rect 80 243 110 452
rect 166 425 196 565
rect 152 409 210 425
rect 152 375 166 409
rect 200 375 210 409
rect 152 359 210 375
rect 152 243 182 359
rect 80 89 110 115
rect 152 89 182 115
<< polycont >>
rect 47 468 81 502
rect 166 375 200 409
<< locali >>
rect 0 1089 286 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 286 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 121 949 155 965
rect 47 502 81 597
rect 47 452 81 468
rect 207 949 241 1049
rect 207 657 241 673
rect 121 483 155 605
rect 195 409 229 523
rect 150 375 166 409
rect 200 375 229 409
rect 35 215 69 227
rect 35 115 69 131
rect 193 215 227 231
rect 193 61 227 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 47 597 81 631
rect 121 449 155 483
rect 195 523 229 557
rect 35 227 69 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 286 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 286 1089
rect 0 1049 286 1055
rect 35 631 93 637
rect 35 597 47 631
rect 81 597 115 631
rect 35 591 93 597
rect 183 557 241 563
rect 161 523 195 557
rect 229 523 241 557
rect 183 517 241 523
rect 109 483 167 489
rect 109 449 121 483
rect 155 449 167 483
rect 109 443 167 449
rect 23 261 81 267
rect 121 261 155 443
rect 23 227 35 261
rect 69 227 155 261
rect 23 221 81 227
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 136 418 136 418 1 Y
port 1 n
rlabel viali 64 614 64 614 1 A
port 2 n
rlabel viali 212 540 212 540 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
