* File: sky130_osu_sc_15T_ls__oai21_l.pex.spice
* Created: Fri Nov 12 14:58:55 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%GND 1 17 19 26 35 38
r37 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r38 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r39 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r40 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r41 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r42 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r43 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r44 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r45 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%VDD 1 13 15 21 26 29 32
r26 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r27 26 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r28 19 26 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.05 $Y=5.245
+ $X2=1.05 $Y2=5.397
r29 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.05 $Y=5.245
+ $X2=1.05 $Y2=4.225
r30 15 26 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=5.397
+ $X2=1.05 $Y2=5.397
r31 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=5.397
+ $X2=0.34 $Y2=5.397
r32 13 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r33 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r34 1 21 300 $w=1.7e-07 $l=1.46833e-06 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.825 $X2=1.05 $Y2=4.225
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%A0 3 5 8 12 15 16 19 25
r37 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.415 $Y=3.07
+ $X2=0.415 $Y2=3.07
r38 19 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.415 $Y=2.5
+ $X2=0.415 $Y2=3.07
r39 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=2.5 $X2=0.415 $Y2=2.5
r40 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.5
+ $X2=0.415 $Y2=2.665
r41 15 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.5
+ $X2=0.415 $Y2=2.335
r42 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=0.355 $Y=1.515
+ $X2=0.475 $Y2=1.515
r43 8 17 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.665
r44 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=1.515
r45 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=0.945
r46 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.355 $Y=1.59
+ $X2=0.355 $Y2=1.515
r47 1 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.355 $Y=1.59
+ $X2=0.355 $Y2=2.335
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%A1 3 7 10 15 18 22
r55 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.895 $Y=2.7
+ $X2=0.895 $Y2=2.7
r56 18 19 5.0779 $w=2.18e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.7 $X2=0.87
+ $Y2=2.615
r57 15 19 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.845 $Y=1.96
+ $X2=0.845 $Y2=2.615
r58 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.96 $X2=0.845 $Y2=1.96
r59 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.845 $Y=1.96
+ $X2=0.845 $Y2=2.095
r60 10 11 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.845 $Y=1.96
+ $X2=0.845 $Y2=1.825
r61 7 11 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=1.825
r62 3 12 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=0.835 $Y=3.825
+ $X2=0.835 $Y2=2.095
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%B0 1 3 7 13 15 17 20
r52 15 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.285 $Y=1.62
+ $X2=1.395 $Y2=1.62
r53 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.33 $X2=1.2
+ $Y2=2.33
r54 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=1.705
+ $X2=1.285 $Y2=1.62
r55 11 13 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.2 $Y=1.705
+ $X2=1.2 $Y2=2.33
r56 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.62 $X2=1.395 $Y2=1.62
r57 5 10 38.8629 $w=2.72e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.335 $Y=1.455
+ $X2=1.39 $Y2=1.62
r58 5 7 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.335 $Y=1.455
+ $X2=1.335 $Y2=0.945
r59 1 10 38.8629 $w=2.72e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.325 $Y=1.785
+ $X2=1.39 $Y2=1.62
r60 1 3 1235.77 $w=1.5e-07 $l=2.41e-06 $layer=POLY_cond $X=1.325 $Y=1.785
+ $X2=1.325 $Y2=4.195
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%Y 1 3 4 15 19 20 23 27 30 35 39 40 45
r57 39 40 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.54 $Y=1.96
+ $X2=1.54 $Y2=1.845
r58 36 45 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r59 36 40 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.845
r60 33 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r61 30 33 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.55 $Y=0.86
+ $X2=1.55 $Y2=1.22
r62 25 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.495
+ $X2=1.54 $Y2=3.41
r63 25 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.54 $Y=3.495
+ $X2=1.54 $Y2=4.225
r64 23 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.54 $Y=1.96
+ $X2=1.54 $Y2=1.96
r65 21 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.325
+ $X2=1.54 $Y2=3.41
r66 21 23 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.54 $Y=3.325
+ $X2=1.54 $Y2=1.96
r67 19 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=3.41
+ $X2=1.54 $Y2=3.41
r68 19 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.455 $Y=3.41
+ $X2=0.345 $Y2=3.41
r69 15 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r70 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.495
+ $X2=0.345 $Y2=3.41
r71 13 15 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.26 $Y=3.495
+ $X2=0.26 $Y2=3.885
r72 4 27 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=3.565 $X2=1.54 $Y2=4.225
r73 3 17 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r74 3 15 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
r75 1 30 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.86
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__OAI21_L%A_27_115# 1 2 11 13 14 17
r14 15 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.12 $Y=1.075
+ $X2=1.12 $Y2=0.865
r15 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=1.12 $Y2=1.075
r16 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.345 $Y2=1.16
r17 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.345 $Y2=1.16
r18 9 11 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.26 $Y2=0.865
r19 2 17 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r20 1 11 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

