* File: sky130_osu_sc_15T_hs__inv_2.spice
* Created: Fri Nov 12 14:30:42 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__inv_2.pex.spice"
.subckt sky130_osu_sc_15T_hs__inv_2  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1000 N_GND_M1000_d N_A_M1000_g N_Y_M1000_s N_GND_M1000_b NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1000_s N_GND_M1000_b NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_Y_M1001_s N_VDD_M1001_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g N_Y_M1001_s N_VDD_M1001_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX4_noxref N_GND_M1000_b N_VDD_M1001_b NWDIODE A=4.366 P=8.86
pX5_noxref noxref_5 A A PROBETYPE=1
pX6_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__inv_2.pxi.spice"
*
.ends
*
*
