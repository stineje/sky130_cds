* File: sky130_osu_sc_18T_hs__and2_1.pex.spice
* Created: Thu Oct 29 17:05:45 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__AND2_1%GND 1 12 14 21 26 29
r36 26 29 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r37 19 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r38 12 19 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r39 12 14 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r40 12 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r41 12 14 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r42 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__AND2_1%VDD 1 2 13 17 23 32 33 35 38
r29 38 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r30 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r31 32 42 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r32 32 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r33 29 42 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r34 29 31 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r35 23 26 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r36 21 33 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r37 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r38 17 20 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r39 15 31 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r40 15 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r41 13 42 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r42 13 31 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r43 2 26 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r44 2 23 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r45 1 20 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r46 1 17 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__AND2_1%A 3 7 12 15 18
r32 16 18 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.765
+ $X2=0.475 $Y2=2.765
r33 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.765 $X2=0.27 $Y2=2.765
r34 11 15 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=2.765
r35 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r36 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=2.765
r37 5 7 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=4.585
r38 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=2.765
r39 1 3 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__AND2_1%B 3 7 12 15 16
r41 16 18 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.59
r42 16 17 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.26
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.425 $X2=0.95 $Y2=2.425
r44 11 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.425
r45 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.96
r46 7 18 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.59
r47 3 17 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__AND2_1%A_27_115# 1 2 9 13 14 16 17 20 22 23 28
+ 34 37 38 39
r69 38 39 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.545
+ $X2=0.65 $Y2=3.715
r70 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r71 32 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=0.61 $Y2=1.935
r72 32 34 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=1.43 $Y2=1.935
r73 28 30 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.69 $Y=3.795
+ $X2=0.69 $Y2=5.835
r74 28 39 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.795 $X2=0.69
+ $Y2=3.715
r75 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=2.02 $X2=0.61
+ $Y2=1.935
r76 24 38 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r77 22 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.61 $Y2=1.935
r78 22 23 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.345 $Y2=1.935
r79 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.345 $Y2=1.935
r80 18 20 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r81 16 17 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.81
+ $X2=1.352 $Y2=2.96
r82 14 35 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.412 $Y2=1.935
r83 14 16 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1 $X2=1.37
+ $Y2=2.81
r84 13 17 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.96
r85 7 35 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.412 $Y2=1.935
r86 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r87 2 30 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r88 2 28 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.795
r89 1 20 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__AND2_1%Y 1 2 10 13 17 18 21
r35 28 30 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r36 18 28 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r37 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r38 14 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r39 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r40 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r41 8 10 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r42 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r43 7 10 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r44 2 30 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r45 2 28 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r46 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

