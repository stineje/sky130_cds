* File: sky130_osu_sc_18T_hs__xnor2_l.spice
* Created: Thu Oct 29 17:10:38 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_hs__xnor2_l.pex.spice"
.subckt sky130_osu_sc_18T_hs__xnor2_l  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1001 A_196_115# N_A_M1001_g N_GND_M1004_d N_GND_M1004_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1011 N_Y_M1011_d N_A_238_89#_M1011_g A_196_115# N_GND_M1004_b NLOWVT L=0.15
+ W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1 R=6.66667
+ SA=75001 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1007 A_388_115# N_A_27_115#_M1007_g N_Y_M1011_d N_GND_M1004_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.6 SB=75001 A=0.15 P=2.3 MULT=1
MM1009 N_GND_M1009_d N_B_M1009_g A_388_115# N_GND_M1004_b NLOWVT L=0.15 W=1
+ AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_238_89#_M1005_d N_B_M1005_g N_GND_M1009_d N_GND_M1004_b NLOWVT L=0.15
+ W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_VDD_M1002_d N_A_M1002_g N_A_27_115#_M1002_s N_VDD_M1002_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75002.4 A=0.45 P=6.3 MULT=1
MM1000 A_196_617# N_A_27_115#_M1000_g N_VDD_M1002_d N_VDD_M1002_b PSHORT L=0.15
+ W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.6
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1010 N_Y_M1010_d N_A_238_89#_M1010_g A_196_617# N_VDD_M1002_b PSHORT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20 SA=75001
+ SB=75001.6 A=0.45 P=6.3 MULT=1
MM1006 A_388_617# N_A_M1006_g N_Y_M1010_d N_VDD_M1002_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20 SA=75001.6
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1008 N_VDD_M1008_d N_B_M1008_g A_388_617# N_VDD_M1002_b PSHORT L=0.15 W=3
+ AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.9
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1003 N_A_238_89#_M1003_d N_B_M1003_g N_VDD_M1008_d N_VDD_M1002_b PSHORT L=0.15
+ W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.4
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX12_noxref N_GND_M1004_b N_VDD_M1002_b NWDIODE A=12.293 P=14.07
pX13_noxref noxref_12 A A PROBETYPE=1
pX14_noxref noxref_13 Y Y PROBETYPE=1
pX15_noxref noxref_14 B B PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__xnor2_l.pxi.spice"
*
.ends
*
*
