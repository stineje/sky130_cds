* File: sky130_osu_sc_18T_ms__nand2_1.pxi.spice
* Created: Thu Oct 29 17:30:30 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__NAND2_1%GND N_GND_M1001_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_9_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_MS__NAND2_1%GND
x_PM_SKY130_OSU_SC_18T_MS__NAND2_1%VDD N_VDD_M1003_s N_VDD_M1000_d N_VDD_M1003_b
+ N_VDD_c_27_p N_VDD_c_36_p N_VDD_c_28_p VDD N_VDD_c_29_p
+ PM_SKY130_OSU_SC_18T_MS__NAND2_1%VDD
x_PM_SKY130_OSU_SC_18T_MS__NAND2_1%A N_A_M1002_g N_A_M1003_g A N_A_c_50_n
+ N_A_c_51_n PM_SKY130_OSU_SC_18T_MS__NAND2_1%A
x_PM_SKY130_OSU_SC_18T_MS__NAND2_1%B N_B_M1001_g N_B_M1000_g N_B_c_82_n
+ N_B_c_84_n B N_B_c_86_n PM_SKY130_OSU_SC_18T_MS__NAND2_1%B
x_PM_SKY130_OSU_SC_18T_MS__NAND2_1%Y N_Y_M1002_s N_Y_M1003_d N_Y_c_115_n
+ N_Y_c_116_n Y N_Y_c_119_n N_Y_c_120_n N_Y_c_121_n
+ PM_SKY130_OSU_SC_18T_MS__NAND2_1%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.0889283f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=1.075
cc_4 N_GND_M1002_b N_A_M1003_g 0.00342256f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_5 N_GND_M1002_b N_A_c_50_n 0.00856875f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.685
cc_6 N_GND_M1002_b N_A_c_51_n 0.0490341f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.685
cc_7 N_GND_M1002_b N_B_M1001_g 0.0461967f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_8 N_GND_c_2_p N_B_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=1.075
cc_9 N_GND_c_9_p N_B_M1001_g 0.00713292f $X=1.05 $Y=0.825 $X2=0.835 $Y2=1.075
cc_10 N_GND_c_3_p N_B_M1001_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.835 $Y2=1.075
cc_11 N_GND_M1002_b N_B_M1000_g 0.0316271f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_12 N_GND_M1002_b N_B_c_82_n 0.0353546f $X=-0.045 $Y=0 $X2=0.915 $Y2=2.22
cc_13 N_GND_c_9_p N_B_c_82_n 0.00231535f $X=1.05 $Y=0.825 $X2=0.915 $Y2=2.22
cc_14 N_GND_M1002_b N_B_c_84_n 0.0122574f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.22
cc_15 N_GND_M1002_b B 0.00492682f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.96
cc_16 N_GND_M1002_b N_B_c_86_n 0.0195876f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.96
cc_17 N_GND_c_9_p N_Y_c_115_n 6.82281e-19 $X=1.05 $Y=0.825 $X2=0.605 $Y2=1.48
cc_18 N_GND_M1002_b N_Y_c_116_n 0.0206417f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.48
cc_19 N_GND_c_9_p N_Y_c_116_n 5.67165e-19 $X=1.05 $Y=0.825 $X2=0.405 $Y2=1.48
cc_20 N_GND_M1002_b Y 0.013296f $X=-0.045 $Y=0 $X2=0.68 $Y2=2.35
cc_21 N_GND_M1002_b N_Y_c_119_n 0.00518799f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.59
cc_22 N_GND_M1002_b N_Y_c_120_n 0.00851145f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.59
cc_23 N_GND_M1002_b N_Y_c_121_n 0.00156053f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.825
cc_24 N_GND_c_2_p N_Y_c_121_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26 $Y2=0.825
cc_25 N_GND_c_3_p N_Y_c_121_n 0.00476261f $X=1.02 $Y=0.17 $X2=0.26 $Y2=0.825
cc_26 N_VDD_M1003_b N_A_M1003_g 0.0225637f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_27 N_VDD_c_27_p N_A_M1003_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_28 N_VDD_c_28_p N_A_M1003_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=4.585
cc_29 N_VDD_c_29_p N_A_M1003_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=4.585
cc_30 N_VDD_M1003_s A 0.0150401f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_31 N_VDD_c_27_p A 0.00522047f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_32 N_VDD_M1003_s N_A_c_50_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32 $Y2=2.685
cc_33 N_VDD_M1003_b N_A_c_50_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=2.685
cc_34 N_VDD_c_27_p N_A_c_50_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=2.685
cc_35 N_VDD_M1003_b N_B_M1000_g 0.0222331f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_36 N_VDD_c_36_p N_B_M1000_g 0.00713292f $X=1.12 $Y=3.795 $X2=0.905 $Y2=4.585
cc_37 N_VDD_c_28_p N_B_M1000_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=4.585
cc_38 N_VDD_c_29_p N_B_M1000_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.905 $Y2=4.585
cc_39 N_VDD_M1003_b B 0.012337f $X=-0.045 $Y=2.905 $X2=1.06 $Y2=2.96
cc_40 N_VDD_c_36_p B 0.00509939f $X=1.12 $Y=3.795 $X2=1.06 $Y2=2.96
cc_41 N_VDD_M1003_b N_B_c_86_n 0.00337476f $X=-0.045 $Y=2.905 $X2=1.06 $Y2=2.96
cc_42 N_VDD_c_36_p N_B_c_86_n 0.00252359f $X=1.12 $Y=3.795 $X2=1.06 $Y2=2.96
cc_43 N_VDD_M1003_b N_Y_c_120_n 0.00458137f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.59
cc_44 N_VDD_c_28_p N_Y_c_120_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69 $Y2=2.59
cc_45 N_VDD_c_29_p N_Y_c_120_n 0.00475776f $X=1.02 $Y=6.49 $X2=0.69 $Y2=2.59
cc_46 N_A_M1002_g N_B_M1001_g 0.120558f $X=0.475 $Y=1.075 $X2=0.835 $Y2=1.075
cc_47 N_A_M1002_g N_B_M1000_g 0.0440961f $X=0.475 $Y=1.075 $X2=0.905 $Y2=4.585
cc_48 N_A_M1002_g N_B_c_84_n 0.00282768f $X=0.475 $Y=1.075 $X2=1.06 $Y2=2.22
cc_49 N_A_M1002_g N_B_c_86_n 0.00112963f $X=0.475 $Y=1.075 $X2=1.06 $Y2=2.96
cc_50 A N_Y_M1003_d 0.00263091f $X=0.32 $Y=3.33 $X2=0.55 $Y2=3.085
cc_51 N_A_M1002_g N_Y_c_115_n 0.0136921f $X=0.475 $Y=1.075 $X2=0.605 $Y2=1.48
cc_52 N_A_M1002_g N_Y_c_116_n 0.00380596f $X=0.475 $Y=1.075 $X2=0.405 $Y2=1.48
cc_53 N_A_M1002_g Y 0.0123501f $X=0.475 $Y=1.075 $X2=0.68 $Y2=2.35
cc_54 N_A_M1002_g N_Y_c_119_n 0.00216533f $X=0.475 $Y=1.075 $X2=0.69 $Y2=2.59
cc_55 A N_Y_c_119_n 0.00150969f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.59
cc_56 N_A_c_50_n N_Y_c_119_n 0.00474021f $X=0.32 $Y=2.685 $X2=0.69 $Y2=2.59
cc_57 N_A_c_51_n N_Y_c_119_n 0.00278592f $X=0.32 $Y=2.685 $X2=0.69 $Y2=2.59
cc_58 N_A_M1002_g N_Y_c_120_n 0.00546744f $X=0.475 $Y=1.075 $X2=0.69 $Y2=2.59
cc_59 A N_Y_c_120_n 0.00831114f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.59
cc_60 N_A_c_50_n N_Y_c_120_n 0.0420549f $X=0.32 $Y=2.685 $X2=0.69 $Y2=2.59
cc_61 N_A_M1002_g N_Y_c_121_n 0.00587516f $X=0.475 $Y=1.075 $X2=0.26 $Y2=0.825
cc_62 N_B_M1001_g N_Y_c_115_n 0.00790819f $X=0.835 $Y=1.075 $X2=0.605 $Y2=1.48
cc_63 N_B_M1001_g Y 0.0185298f $X=0.835 $Y=1.075 $X2=0.68 $Y2=2.35
cc_64 N_B_M1000_g Y 0.00128442f $X=0.905 $Y=4.585 $X2=0.68 $Y2=2.35
cc_65 N_B_c_82_n Y 0.00398874f $X=0.915 $Y=2.22 $X2=0.68 $Y2=2.35
cc_66 N_B_c_84_n Y 0.0139756f $X=1.06 $Y=2.22 $X2=0.68 $Y2=2.35
cc_67 N_B_c_86_n Y 0.0066619f $X=1.06 $Y=2.96 $X2=0.68 $Y2=2.35
cc_68 N_B_M1000_g N_Y_c_119_n 0.00339349f $X=0.905 $Y=4.585 $X2=0.69 $Y2=2.59
cc_69 N_B_c_82_n N_Y_c_119_n 0.00170653f $X=0.915 $Y=2.22 $X2=0.69 $Y2=2.59
cc_70 N_B_c_84_n N_Y_c_119_n 0.00261701f $X=1.06 $Y=2.22 $X2=0.69 $Y2=2.59
cc_71 B N_Y_c_119_n 0.0028041f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_72 N_B_c_86_n N_Y_c_119_n 0.00640429f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_73 N_B_M1000_g N_Y_c_120_n 0.00560092f $X=0.905 $Y=4.585 $X2=0.69 $Y2=2.59
cc_74 N_B_c_82_n N_Y_c_120_n 2.88224e-19 $X=0.915 $Y=2.22 $X2=0.69 $Y2=2.59
cc_75 N_B_c_84_n N_Y_c_120_n 0.00144012f $X=1.06 $Y=2.22 $X2=0.69 $Y2=2.59
cc_76 B N_Y_c_120_n 0.00831114f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_77 N_B_c_86_n N_Y_c_120_n 0.0295869f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_78 N_Y_c_115_n A_110_115# 0.0109071f $X=0.605 $Y=1.48 $X2=0.55 $Y2=0.575
