* File: sky130_osu_sc_18T_ms__inv_1.pxi.spice
* Created: Fri Nov 12 14:04:05 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__INV_1%GND N_GND_M1000_s N_GND_M1000_b N_GND_c_2_p
+ N_GND_c_3_p GND PM_SKY130_OSU_SC_18T_MS__INV_1%GND
x_PM_SKY130_OSU_SC_18T_MS__INV_1%VDD N_VDD_M1001_s N_VDD_M1001_b N_VDD_c_17_p
+ N_VDD_c_18_p VDD PM_SKY130_OSU_SC_18T_MS__INV_1%VDD
x_PM_SKY130_OSU_SC_18T_MS__INV_1%A N_A_M1000_g N_A_M1001_g N_A_c_33_n N_A_c_34_n
+ N_A_c_35_n N_A_c_36_n A PM_SKY130_OSU_SC_18T_MS__INV_1%A
x_PM_SKY130_OSU_SC_18T_MS__INV_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_67_n N_Y_c_69_n
+ Y N_Y_c_71_n N_Y_c_73_n PM_SKY130_OSU_SC_18T_MS__INV_1%Y
cc_1 N_GND_M1000_b N_A_M1000_g 0.0750619f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1000_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1000_g 0.00468827f $X=0.34 $Y=0.19 $X2=0.475 $Y2=1.075
cc_4 N_GND_M1000_b N_A_M1001_g 0.0337175f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_5 N_GND_M1000_b N_A_c_33_n 0.0393936f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_6 N_GND_M1000_b N_A_c_34_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.33
cc_7 N_GND_M1000_b N_A_c_35_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.305
cc_8 N_GND_M1000_b N_A_c_36_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_9 N_GND_M1000_b N_Y_c_67_n 0.00913846f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_10 N_GND_c_3_p N_Y_c_67_n 0.00476261f $X=0.34 $Y=0.19 $X2=0.69 $Y2=0.825
cc_11 N_GND_M1000_b N_Y_c_69_n 0.00237997f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_12 N_GND_M1000_b Y 0.0587019f $X=-0.045 $Y=0 $X2=0.755 $Y2=2.205
cc_13 N_GND_M1000_b N_Y_c_71_n 0.0126319f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.48
cc_14 N_GND_c_2_p N_Y_c_71_n 0.00125659f $X=0.26 $Y=0.825 $X2=0.69 $Y2=1.48
cc_15 N_GND_M1000_b N_Y_c_73_n 0.00507896f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_16 N_VDD_M1001_b N_A_M1001_g 0.028768f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=4.585
cc_17 N_VDD_c_17_p N_A_M1001_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_18 N_VDD_c_18_p N_A_M1001_g 0.00606474f $X=0.34 $Y=6.47 $X2=0.475 $Y2=4.585
cc_19 VDD N_A_M1001_g 0.00468827f $X=0.34 $Y=6.42 $X2=0.475 $Y2=4.585
cc_20 N_VDD_M1001_s N_A_c_34_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_21 N_VDD_M1001_b N_A_c_34_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=3.33
cc_22 N_VDD_c_17_p N_A_c_34_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_23 N_VDD_M1001_s A 0.0162774f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_24 N_VDD_c_17_p A 0.00522047f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_25 N_VDD_M1001_b N_Y_c_69_n 0.00592536f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_26 N_VDD_c_18_p N_Y_c_69_n 0.00757793f $X=0.34 $Y=6.47 $X2=0.69 $Y2=2.96
cc_27 VDD N_Y_c_69_n 0.00476261f $X=0.34 $Y=6.42 $X2=0.69 $Y2=2.96
cc_28 N_VDD_M1001_b N_Y_c_73_n 0.00914195f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_29 A N_Y_M1001_d 0.00251573f $X=0.32 $Y=3.33 $X2=0.55 $Y2=3.085
cc_30 N_A_M1000_g N_Y_c_67_n 0.0057847f $X=0.475 $Y=1.075 $X2=0.69 $Y2=0.825
cc_31 N_A_c_33_n N_Y_c_67_n 6.24081e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_32 N_A_c_36_n N_Y_c_67_n 0.00110256f $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_33 N_A_M1001_g N_Y_c_69_n 0.00866213f $X=0.475 $Y=4.585 $X2=0.69 $Y2=2.96
cc_34 N_A_c_33_n N_Y_c_69_n 8.13098e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_35 N_A_c_34_n N_Y_c_69_n 0.0228882f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_36 N_A_c_36_n N_Y_c_69_n 0.00202105f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_37 A N_Y_c_69_n 0.0149533f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_38 N_A_M1000_g Y 0.0127139f $X=0.475 $Y=1.075 $X2=0.755 $Y2=2.205
cc_39 N_A_M1001_g Y 0.00874077f $X=0.475 $Y=4.585 $X2=0.755 $Y2=2.205
cc_40 N_A_c_33_n Y 0.00719822f $X=0.535 $Y=2.305 $X2=0.755 $Y2=2.205
cc_41 N_A_c_34_n Y 0.0183799f $X=0.32 $Y=3.33 $X2=0.755 $Y2=2.205
cc_42 N_A_c_36_n Y 0.0178517f $X=0.535 $Y=2.305 $X2=0.755 $Y2=2.205
cc_43 N_A_M1000_g N_Y_c_71_n 0.0105261f $X=0.475 $Y=1.075 $X2=0.69 $Y2=1.48
cc_44 N_A_c_33_n N_Y_c_71_n 0.0011424f $X=0.535 $Y=2.305 $X2=0.69 $Y2=1.48
cc_45 N_A_M1001_g N_Y_c_73_n 0.00478745f $X=0.475 $Y=4.585 $X2=0.69 $Y2=2.96
cc_46 N_A_c_33_n N_Y_c_73_n 0.00126139f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_47 N_A_c_34_n N_Y_c_73_n 0.00640429f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_48 N_A_c_36_n N_Y_c_73_n 0.00194461f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_49 A N_Y_c_73_n 0.00815006f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
