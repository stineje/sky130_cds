* File: sky130_osu_sc_15T_hs__inv_10.pex.spice
* Created: Fri Nov 12 14:30:25 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__INV_10%GND 1 2 3 4 5 6 67 71 73 80 82 89 91 98
+ 100 107 109 117 132 134
r142 132 134 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r143 115 117 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.56 $Y2=0.865
r144 109 115 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.475
+ $Y=0.152 $X2=4.56 $Y2=0.305
r145 105 107 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.865
r146 101 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r147 96 125 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r148 96 98 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.865
r149 92 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r150 91 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r151 87 124 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r152 87 89 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.865
r153 83 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r154 82 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r155 78 123 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r156 78 80 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.865
r157 73 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r158 69 71 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r159 67 134 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r160 67 132 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r161 67 105 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.7 $Y2=0.305
r162 67 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.615 $Y2=0.152
r163 67 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.785 $Y2=0.152
r164 67 69 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r165 67 74 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r166 67 109 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.475 $Y2=0.152
r167 67 110 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=3.785 $Y2=0.152
r168 67 100 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r169 67 101 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r170 67 91 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r171 67 92 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r172 67 82 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r173 67 83 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r174 67 73 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r175 67 74 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r176 6 117 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.575 $X2=4.56 $Y2=0.865
r177 5 107 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.865
r178 4 98 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.865
r179 3 89 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.865
r180 2 80 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r181 1 71 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__INV_10%VDD 1 2 3 4 5 6 53 57 61 67 71 77 81 87
+ 91 97 101 108 121 125
r96 121 125 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=4.42 $Y2=5.397
r97 113 121 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r98 108 111 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.56 $Y=3.205
+ $X2=4.56 $Y2=4.565
r99 106 111 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.56 $Y=5.245
+ $X2=4.56 $Y2=4.565
r100 104 125 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=5.36
+ $X2=4.42 $Y2=5.36
r101 102 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=5.397
+ $X2=3.7 $Y2=5.397
r102 102 104 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=5.397
+ $X2=4.42 $Y2=5.397
r103 101 106 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.475 $Y=5.397
+ $X2=4.56 $Y2=5.245
r104 101 104 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.475 $Y=5.397
+ $X2=4.42 $Y2=5.397
r105 97 100 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.7 $Y=3.205
+ $X2=3.7 $Y2=4.565
r106 95 119 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.7 $Y=5.245
+ $X2=3.7 $Y2=5.397
r107 95 100 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=5.245
+ $X2=3.7 $Y2=4.565
r108 92 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=2.84 $Y2=5.397
r109 92 94 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=3.06 $Y2=5.397
r110 91 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.7 $Y2=5.397
r111 91 94 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.06 $Y2=5.397
r112 87 90 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.205
+ $X2=2.84 $Y2=4.565
r113 85 117 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=5.397
r114 85 90 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.565
r115 82 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r116 82 84 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r117 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.397
r118 81 84 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r119 77 80 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.205
+ $X2=1.98 $Y2=4.565
r120 75 116 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r121 75 80 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.565
r122 72 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r123 72 74 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r124 71 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r125 71 74 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r126 67 70 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=3.205
+ $X2=1.12 $Y2=4.565
r127 65 115 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r128 65 70 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r129 62 113 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r130 62 64 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r131 61 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r132 61 64 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r133 57 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r134 55 113 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r135 55 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r136 53 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=5.245 $X2=4.42 $Y2=5.33
r137 53 119 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r138 53 94 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r139 53 84 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r140 53 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r141 53 64 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r142 53 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r143 6 111 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.825 $X2=4.56 $Y2=4.565
r144 6 108 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.825 $X2=4.56 $Y2=3.205
r145 5 100 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=4.565
r146 5 97 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=3.205
r147 4 90 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.565
r148 4 87 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.205
r149 3 80 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.565
r150 3 77 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.205
r151 2 70 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r152 2 67 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.205
r153 1 60 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r154 1 57 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__INV_10%A 3 8 9 11 12 14 18 20 22 23 25 29 31 33
+ 34 36 40 42 44 45 47 51 54 55 57 58 60 64 66 68 69 71 75 77 79 80 82 86 88 90
+ 91 93 97 99 101 102 104 108 110 112 113 115 116 118 119 120 121 122 123 124
+ 125 126 127 128 129 130 131 132 133 134 137 139 141 144
c289 99 0 1.33323e-19 $X=3.915 $Y=2.7
c290 97 0 1.33323e-19 $X=3.915 $Y=0.895
c291 88 0 1.33323e-19 $X=3.485 $Y=2.7
c292 86 0 1.33323e-19 $X=3.485 $Y=0.895
c293 77 0 1.33323e-19 $X=3.055 $Y=2.7
c294 75 0 1.33323e-19 $X=3.055 $Y=0.895
c295 66 0 1.33323e-19 $X=2.625 $Y=2.7
c296 64 0 1.33323e-19 $X=2.625 $Y=0.895
c297 55 0 1.33323e-19 $X=2.195 $Y=2.7
c298 51 0 1.33323e-19 $X=2.195 $Y=0.895
c299 42 0 1.33323e-19 $X=1.765 $Y=2.7
c300 40 0 1.33323e-19 $X=1.765 $Y=0.895
c301 31 0 1.33323e-19 $X=1.335 $Y=2.7
c302 29 0 1.33323e-19 $X=1.335 $Y=0.895
c303 20 0 1.33323e-19 $X=0.905 $Y=2.7
c304 18 0 1.33323e-19 $X=0.905 $Y=0.895
r305 144 147 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=3.065
+ $X2=0.405 $Y2=3.07
r306 139 141 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.045
+ $X2=0.535 $Y2=2.045
r307 137 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r308 135 139 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.405 $Y2=2.045
r309 135 137 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.13
+ $X2=0.32 $Y2=3.07
r310 115 141 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.045 $X2=0.535 $Y2=2.045
r311 115 117 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=2.21
r312 115 116 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=1.88
r313 110 112 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=4.345 $Y=2.7
+ $X2=4.345 $Y2=3.825
r314 106 108 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.345 $Y=1.44
+ $X2=4.345 $Y2=0.895
r315 105 134 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=2.625
+ $X2=3.915 $Y2=2.625
r316 104 110 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=2.625
+ $X2=4.345 $Y2=2.7
r317 104 105 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=2.625
+ $X2=3.99 $Y2=2.625
r318 103 133 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.515
+ $X2=3.915 $Y2=1.515
r319 102 106 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=1.515
+ $X2=4.345 $Y2=1.44
r320 102 103 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.515
+ $X2=3.99 $Y2=1.515
r321 99 134 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=2.7
+ $X2=3.915 $Y2=2.625
r322 99 101 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.915 $Y=2.7
+ $X2=3.915 $Y2=3.825
r323 95 133 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=1.44
+ $X2=3.915 $Y2=1.515
r324 95 97 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.915 $Y=1.44
+ $X2=3.915 $Y2=0.895
r325 94 132 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.625
+ $X2=3.485 $Y2=2.625
r326 93 134 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.625
+ $X2=3.915 $Y2=2.625
r327 93 94 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.625
+ $X2=3.56 $Y2=2.625
r328 92 131 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.515
+ $X2=3.485 $Y2=1.515
r329 91 133 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.515
+ $X2=3.915 $Y2=1.515
r330 91 92 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.515
+ $X2=3.56 $Y2=1.515
r331 88 132 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=2.625
r332 88 90 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=3.825
r333 84 131 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.485 $Y2=1.515
r334 84 86 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.485 $Y2=0.895
r335 83 130 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.625
+ $X2=3.055 $Y2=2.625
r336 82 132 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.485 $Y2=2.625
r337 82 83 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.13 $Y2=2.625
r338 81 129 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.055 $Y2=1.515
r339 80 131 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.515
+ $X2=3.485 $Y2=1.515
r340 80 81 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.515
+ $X2=3.13 $Y2=1.515
r341 77 130 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=2.625
r342 77 79 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=3.825
r343 73 129 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=1.515
r344 73 75 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=0.895
r345 72 128 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.625
+ $X2=2.625 $Y2=2.625
r346 71 130 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=3.055 $Y2=2.625
r347 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=2.7 $Y2=2.625
r348 70 127 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.625 $Y2=1.515
r349 69 129 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=3.055 $Y2=1.515
r350 69 70 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=2.7 $Y2=1.515
r351 66 128 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=2.625
r352 66 68 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r353 62 127 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=1.515
r354 62 64 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.625 $Y=1.44
+ $X2=2.625 $Y2=0.895
r355 61 126 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r356 60 128 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.625
r357 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r358 59 125 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.515
+ $X2=2.195 $Y2=1.515
r359 58 127 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.625 $Y2=1.515
r360 58 59 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.27 $Y2=1.515
r361 55 126 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=2.625
r362 55 57 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r363 54 126 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.55
+ $X2=2.195 $Y2=2.625
r364 53 125 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.59
+ $X2=2.195 $Y2=1.515
r365 53 54 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.59
+ $X2=2.195 $Y2=2.55
r366 49 125 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.44
+ $X2=2.195 $Y2=1.515
r367 49 51 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.195 $Y=1.44
+ $X2=2.195 $Y2=0.895
r368 48 124 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r369 47 126 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r370 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r371 46 123 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.515
+ $X2=1.765 $Y2=1.515
r372 45 125 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.515
+ $X2=2.195 $Y2=1.515
r373 45 46 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.515
+ $X2=1.84 $Y2=1.515
r374 42 124 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r375 42 44 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r376 38 123 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.44
+ $X2=1.765 $Y2=1.515
r377 38 40 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.765 $Y=1.44
+ $X2=1.765 $Y2=0.895
r378 37 122 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.625
+ $X2=1.335 $Y2=2.625
r379 36 124 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r380 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.41 $Y2=2.625
r381 35 121 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.335 $Y2=1.515
r382 34 123 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.765 $Y2=1.515
r383 34 35 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.41 $Y2=1.515
r384 31 122 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=2.625
r385 31 33 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r386 27 121 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.44
+ $X2=1.335 $Y2=1.515
r387 27 29 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.335 $Y=1.44
+ $X2=1.335 $Y2=0.895
r388 26 120 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.625
+ $X2=0.905 $Y2=2.625
r389 25 122 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.625
+ $X2=1.335 $Y2=2.625
r390 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.625
+ $X2=0.98 $Y2=2.625
r391 24 119 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.515
+ $X2=0.905 $Y2=1.515
r392 23 121 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=1.335 $Y2=1.515
r393 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=0.98 $Y2=1.515
r394 20 120 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.7
+ $X2=0.905 $Y2=2.625
r395 20 22 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=2.7
+ $X2=0.905 $Y2=3.825
r396 16 119 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.44
+ $X2=0.905 $Y2=1.515
r397 16 18 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.905 $Y=1.44
+ $X2=0.905 $Y2=0.895
r398 15 118 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.625
+ $X2=0.475 $Y2=2.625
r399 14 120 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.625
+ $X2=0.905 $Y2=2.625
r400 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.625
+ $X2=0.55 $Y2=2.625
r401 13 113 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.515
+ $X2=0.475 $Y2=1.515
r402 12 119 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.515
+ $X2=0.905 $Y2=1.515
r403 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.515
+ $X2=0.55 $Y2=1.515
r404 9 118 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.7
+ $X2=0.475 $Y2=2.625
r405 9 11 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.475 $Y=2.7
+ $X2=0.475 $Y2=3.825
r406 8 118 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.55
+ $X2=0.475 $Y2=2.625
r407 8 117 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.55
+ $X2=0.475 $Y2=2.21
r408 5 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.59
+ $X2=0.475 $Y2=1.515
r409 5 116 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.59
+ $X2=0.475 $Y2=1.88
r410 1 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=1.515
r411 1 3 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.475 $Y=1.44
+ $X2=0.475 $Y2=0.895
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__INV_10%Y 1 2 3 4 5 11 12 13 14 15 42 48 56 62
+ 70 76 84 90 98 104 111 112 114 116 118 121 122 123 124 125 127 128 129 130 131
+ 133 134 135 136 137 138 139
c217 139 0 1.33323e-19 $X=4.13 $Y=2.585
c218 138 0 1.33323e-19 $X=4.13 $Y=1.335
c219 137 0 2.66647e-19 $X=3.415 $Y=2.7
c220 135 0 2.66647e-19 $X=3.415 $Y=1.22
c221 131 0 2.66647e-19 $X=2.555 $Y=2.7
c222 129 0 2.66647e-19 $X=2.555 $Y=1.22
c223 125 0 2.66647e-19 $X=1.695 $Y=2.7
c224 123 0 2.66647e-19 $X=1.695 $Y=1.22
c225 112 0 1.33323e-19 $X=0.69 $Y=2.585
c226 111 0 1.33323e-19 $X=0.69 $Y=1.335
r227 139 159 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=2.585
+ $X2=4.13 $Y2=2.7
r228 138 157 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.335
+ $X2=4.13 $Y2=1.22
r229 138 139 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=4.13 $Y=1.335
+ $X2=4.13 $Y2=2.585
r230 137 155 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=2.7
+ $X2=3.27 $Y2=2.7
r231 136 159 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=2.7
+ $X2=4.13 $Y2=2.7
r232 136 137 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=2.7
+ $X2=3.415 $Y2=2.7
r233 135 153 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=1.22
+ $X2=3.27 $Y2=1.22
r234 134 157 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=1.22
+ $X2=4.13 $Y2=1.22
r235 134 135 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=1.22
+ $X2=3.415 $Y2=1.22
r236 133 155 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.585
+ $X2=3.27 $Y2=2.7
r237 132 153 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=1.22
r238 132 133 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=2.585
r239 131 151 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.7
+ $X2=2.41 $Y2=2.7
r240 130 155 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.7
+ $X2=3.27 $Y2=2.7
r241 130 131 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.7
+ $X2=2.555 $Y2=2.7
r242 129 149 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.22
+ $X2=2.41 $Y2=1.22
r243 128 153 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=3.27 $Y2=1.22
r244 128 129 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=2.555 $Y2=1.22
r245 127 151 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.585
+ $X2=2.41 $Y2=2.7
r246 126 149 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r247 126 127 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.585
r248 125 147 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.7
+ $X2=1.55 $Y2=2.7
r249 124 151 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.7
+ $X2=2.41 $Y2=2.7
r250 124 125 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.7
+ $X2=1.695 $Y2=2.7
r251 123 145 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r252 122 149 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r253 122 123 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r254 121 147 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.585
+ $X2=1.55 $Y2=2.7
r255 120 145 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r256 120 121 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=2.585
r257 119 143 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.7
+ $X2=0.69 $Y2=2.7
r258 118 147 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.7
+ $X2=1.55 $Y2=2.7
r259 118 119 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.7
+ $X2=0.835 $Y2=2.7
r260 117 141 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.22
+ $X2=0.69 $Y2=1.22
r261 116 145 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.22
+ $X2=1.55 $Y2=1.22
r262 116 117 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.22
+ $X2=0.835 $Y2=1.22
r263 112 143 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=2.7
r264 112 114 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.585
+ $X2=0.69 $Y2=1.94
r265 111 141 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.22
r266 111 114 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.335
+ $X2=0.69 $Y2=1.94
r267 107 109 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.13 $Y=3.205
+ $X2=4.13 $Y2=4.565
r268 104 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=2.7
+ $X2=4.13 $Y2=2.7
r269 104 107 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.13 $Y=2.7
+ $X2=4.13 $Y2=3.205
r270 101 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=1.22
+ $X2=4.13 $Y2=1.22
r271 98 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.13 $Y=0.865
+ $X2=4.13 $Y2=1.22
r272 93 95 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.27 $Y=3.205
+ $X2=3.27 $Y2=4.565
r273 90 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.7
+ $X2=3.27 $Y2=2.7
r274 90 93 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.27 $Y=2.7
+ $X2=3.27 $Y2=3.205
r275 87 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.22
+ $X2=3.27 $Y2=1.22
r276 84 87 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.27 $Y=0.865
+ $X2=3.27 $Y2=1.22
r277 79 81 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.205
+ $X2=2.41 $Y2=4.565
r278 76 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.7
+ $X2=2.41 $Y2=2.7
r279 76 79 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.41 $Y=2.7
+ $X2=2.41 $Y2=3.205
r280 73 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r281 70 73 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.41 $Y=0.865
+ $X2=2.41 $Y2=1.22
r282 65 67 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.205
+ $X2=1.55 $Y2=4.565
r283 62 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.7
+ $X2=1.55 $Y2=2.7
r284 62 65 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.55 $Y=2.7
+ $X2=1.55 $Y2=3.205
r285 59 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r286 56 59 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.55 $Y=0.865
+ $X2=1.55 $Y2=1.22
r287 51 53 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r288 48 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=2.7
r289 48 51 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.69 $Y=2.7
+ $X2=0.69 $Y2=3.205
r290 45 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.22
+ $X2=0.69 $Y2=1.22
r291 42 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.69 $Y=0.865
+ $X2=0.69 $Y2=1.22
r292 15 109 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.825 $X2=4.13 $Y2=4.565
r293 15 107 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.825 $X2=4.13 $Y2=3.205
r294 14 95 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=4.565
r295 14 93 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=3.205
r296 13 81 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.565
r297 13 79 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.205
r298 12 67 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.565
r299 12 65 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.205
r300 11 53 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r301 11 51 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r302 5 98 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.865
r303 4 84 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.865
r304 3 70 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.865
r305 2 56 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.865
r306 1 42 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

