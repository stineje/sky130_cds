magic
tech sky130A
magscale 1 2
timestamp 1606864598
<< checkpaint >>
rect -1209 -1243 2569 2575
<< nwell >>
rect -9 581 1435 1341
<< nmos >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
rect 338 115 368 315
rect 410 115 440 315
rect 496 115 526 315
rect 582 115 612 315
rect 668 115 698 315
rect 754 115 784 315
rect 840 115 870 315
rect 922 115 952 315
rect 1004 115 1034 315
rect 1102 115 1132 315
rect 1292 115 1322 315
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
rect 338 617 368 1217
rect 410 617 440 1217
rect 496 617 526 1217
rect 582 617 612 1217
rect 668 617 698 1217
rect 754 617 784 1217
rect 840 617 870 1217
rect 922 617 952 1217
rect 1004 617 1034 1217
rect 1102 617 1132 1217
rect 1292 617 1322 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 199 166 315
rect 110 131 121 199
rect 155 131 166 199
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 267 338 315
rect 282 131 293 267
rect 327 131 338 267
rect 282 115 338 131
rect 368 115 410 315
rect 440 267 496 315
rect 440 131 451 267
rect 485 131 496 267
rect 440 115 496 131
rect 526 267 582 315
rect 526 131 537 267
rect 571 131 582 267
rect 526 115 582 131
rect 612 199 668 315
rect 612 131 623 199
rect 657 131 668 199
rect 612 115 668 131
rect 698 267 754 315
rect 698 131 709 267
rect 743 131 754 267
rect 698 115 754 131
rect 784 199 840 315
rect 784 131 795 199
rect 829 131 840 199
rect 784 115 840 131
rect 870 115 922 315
rect 952 115 1004 315
rect 1034 267 1102 315
rect 1034 131 1045 267
rect 1079 131 1102 267
rect 1034 115 1102 131
rect 1132 199 1185 315
rect 1132 131 1143 199
rect 1177 131 1185 199
rect 1132 115 1185 131
rect 1239 199 1292 315
rect 1239 131 1247 199
rect 1281 131 1292 199
rect 1239 115 1292 131
rect 1322 267 1375 315
rect 1322 131 1333 267
rect 1367 131 1375 267
rect 1322 115 1375 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 725 35 1201
rect 69 725 80 1201
rect 27 617 80 725
rect 110 1201 166 1217
rect 110 793 121 1201
rect 155 793 166 1201
rect 110 617 166 793
rect 196 1201 252 1217
rect 196 725 207 1201
rect 241 725 252 1201
rect 196 617 252 725
rect 282 1201 338 1217
rect 282 725 293 1201
rect 327 725 338 1201
rect 282 617 338 725
rect 368 617 410 1217
rect 440 1201 496 1217
rect 440 725 451 1201
rect 485 725 496 1201
rect 440 617 496 725
rect 526 1201 582 1217
rect 526 725 537 1201
rect 571 725 582 1201
rect 526 617 582 725
rect 612 1201 668 1217
rect 612 793 623 1201
rect 657 793 668 1201
rect 612 617 668 793
rect 698 1201 754 1217
rect 698 725 709 1201
rect 743 725 754 1201
rect 698 617 754 725
rect 784 1201 840 1217
rect 784 725 795 1201
rect 829 725 840 1201
rect 784 617 840 725
rect 870 617 922 1217
rect 952 617 1004 1217
rect 1034 1201 1102 1217
rect 1034 793 1045 1201
rect 1079 793 1102 1201
rect 1034 617 1102 793
rect 1132 1201 1185 1217
rect 1132 725 1143 1201
rect 1177 725 1185 1201
rect 1132 617 1185 725
rect 1239 1201 1292 1217
rect 1239 657 1247 1201
rect 1281 657 1292 1201
rect 1239 617 1292 657
rect 1322 1201 1375 1217
rect 1322 657 1333 1201
rect 1367 657 1375 1201
rect 1322 617 1375 657
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 199
rect 207 131 241 267
rect 293 131 327 267
rect 451 131 485 267
rect 537 131 571 267
rect 623 131 657 199
rect 709 131 743 267
rect 795 131 829 199
rect 1045 131 1079 267
rect 1143 131 1177 199
rect 1247 131 1281 199
rect 1333 131 1367 267
<< pdiffc >>
rect 35 725 69 1201
rect 121 793 155 1201
rect 207 725 241 1201
rect 293 725 327 1201
rect 451 725 485 1201
rect 537 725 571 1201
rect 623 793 657 1201
rect 709 725 743 1201
rect 795 725 829 1201
rect 1045 793 1079 1201
rect 1143 725 1177 1201
rect 1247 657 1281 1201
rect 1333 657 1367 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
rect 979 27 1003 61
rect 1037 27 1061 61
rect 1115 27 1139 61
rect 1173 27 1197 61
rect 1251 27 1275 61
rect 1309 27 1333 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
rect 707 1271 731 1305
rect 765 1271 789 1305
rect 843 1271 867 1305
rect 901 1271 925 1305
rect 979 1271 1003 1305
rect 1037 1271 1061 1305
rect 1115 1271 1139 1305
rect 1173 1271 1197 1305
rect 1251 1271 1275 1305
rect 1309 1271 1333 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
rect 1003 27 1037 61
rect 1139 27 1173 61
rect 1275 27 1309 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
rect 731 1271 765 1305
rect 867 1271 901 1305
rect 1003 1271 1037 1305
rect 1139 1271 1173 1305
rect 1275 1271 1309 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1245
rect 338 1217 368 1245
rect 410 1217 440 1243
rect 496 1217 526 1243
rect 582 1217 612 1245
rect 668 1217 698 1245
rect 754 1217 784 1245
rect 840 1217 870 1245
rect 922 1217 952 1245
rect 1004 1217 1034 1245
rect 1102 1217 1132 1245
rect 1292 1217 1322 1245
rect 80 403 110 617
rect 166 585 196 617
rect 152 569 206 585
rect 152 535 162 569
rect 196 535 206 569
rect 152 519 206 535
rect 70 387 124 403
rect 70 353 80 387
rect 114 353 124 387
rect 70 337 124 353
rect 80 315 110 337
rect 166 315 196 519
rect 252 477 282 617
rect 338 519 368 617
rect 410 592 440 617
rect 496 592 526 617
rect 410 562 526 592
rect 338 503 430 519
rect 238 461 292 477
rect 238 427 248 461
rect 282 427 292 461
rect 238 411 292 427
rect 338 469 386 503
rect 420 469 430 503
rect 338 453 430 469
rect 252 315 282 411
rect 338 315 368 453
rect 472 403 502 562
rect 582 403 612 617
rect 668 551 698 617
rect 656 535 710 551
rect 656 501 666 535
rect 700 501 710 535
rect 656 485 710 501
rect 472 387 526 403
rect 472 367 482 387
rect 410 353 482 367
rect 516 353 526 387
rect 410 337 526 353
rect 568 387 622 403
rect 568 353 578 387
rect 612 353 622 387
rect 568 337 622 353
rect 410 315 440 337
rect 496 315 526 337
rect 582 315 612 337
rect 668 315 698 485
rect 754 403 784 617
rect 840 551 870 617
rect 826 535 880 551
rect 826 501 836 535
rect 870 501 880 535
rect 826 485 880 501
rect 922 513 952 617
rect 1004 585 1034 617
rect 1004 555 1048 585
rect 1102 584 1132 617
rect 922 497 976 513
rect 742 387 796 403
rect 742 353 752 387
rect 786 353 796 387
rect 742 337 796 353
rect 754 315 784 337
rect 840 315 870 485
rect 922 463 932 497
rect 966 463 976 497
rect 922 447 976 463
rect 922 315 952 447
rect 1018 403 1048 555
rect 1090 568 1144 584
rect 1292 581 1322 617
rect 1090 534 1100 568
rect 1134 534 1144 568
rect 1090 518 1144 534
rect 1255 565 1322 581
rect 1255 531 1265 565
rect 1299 531 1322 565
rect 1004 387 1058 403
rect 1004 353 1014 387
rect 1048 353 1058 387
rect 1004 337 1058 353
rect 1004 315 1034 337
rect 1102 315 1132 518
rect 1255 515 1322 531
rect 1292 315 1322 515
rect 80 81 110 115
rect 166 82 196 115
rect 252 82 282 115
rect 338 82 368 115
rect 410 82 440 115
rect 496 82 526 115
rect 582 82 612 115
rect 668 82 698 115
rect 754 82 784 115
rect 840 82 870 115
rect 922 82 952 115
rect 1004 82 1034 115
rect 1102 80 1132 115
rect 1292 80 1322 115
<< polycont >>
rect 162 535 196 569
rect 80 353 114 387
rect 248 427 282 461
rect 386 469 420 503
rect 666 501 700 535
rect 482 353 516 387
rect 578 353 612 387
rect 836 501 870 535
rect 752 353 786 387
rect 932 463 966 497
rect 1100 534 1134 568
rect 1265 531 1299 565
rect 1014 353 1048 387
<< locali >>
rect 0 1311 1408 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 595 1311
rect 629 1271 731 1311
rect 765 1271 867 1311
rect 901 1271 1003 1311
rect 1037 1271 1139 1311
rect 1173 1271 1275 1311
rect 1309 1271 1408 1311
rect 35 1201 69 1217
rect 121 1201 155 1271
rect 121 777 155 793
rect 207 1201 241 1217
rect 35 709 69 725
rect 207 709 241 725
rect 35 675 241 709
rect 293 1201 327 1217
rect 293 642 327 725
rect 451 1201 485 1271
rect 451 709 485 725
rect 537 1201 571 1217
rect 623 1201 657 1271
rect 623 777 657 793
rect 709 1201 743 1217
rect 537 708 571 725
rect 709 708 743 725
rect 537 674 743 708
rect 795 1201 829 1217
rect 1045 1201 1079 1271
rect 1045 777 1079 793
rect 1143 1201 1177 1217
rect 795 684 829 725
rect 1143 684 1177 725
rect 795 650 1100 684
rect 293 605 350 642
rect 795 641 829 650
rect 80 535 162 569
rect 196 535 212 569
rect 248 461 282 477
rect 248 411 282 427
rect 64 353 80 387
rect 114 353 130 387
rect 316 370 350 605
rect 752 606 829 641
rect 578 535 612 541
rect 386 503 444 535
rect 420 501 444 503
rect 650 501 666 535
rect 700 501 716 535
rect 386 453 420 469
rect 578 387 612 501
rect 666 461 700 501
rect 752 461 786 606
rect 1066 584 1100 650
rect 1247 1201 1281 1271
rect 1177 650 1202 667
rect 1143 633 1202 650
rect 1247 641 1281 657
rect 1333 1201 1367 1217
rect 1066 568 1134 584
rect 1066 537 1100 568
rect 820 501 836 535
rect 870 501 886 535
rect 1089 534 1100 537
rect 1100 518 1134 534
rect 932 497 966 513
rect 932 461 966 463
rect 1168 461 1202 633
rect 1333 609 1367 657
rect 752 427 879 461
rect 1143 427 1202 461
rect 1265 565 1299 581
rect 293 336 350 370
rect 466 353 482 387
rect 516 353 532 387
rect 736 353 752 387
rect 786 353 811 387
rect 578 337 612 353
rect 293 313 327 336
rect 35 267 241 286
rect 69 252 207 267
rect 35 115 69 131
rect 121 199 155 215
rect 121 61 155 131
rect 207 114 241 131
rect 777 313 811 353
rect 293 267 327 279
rect 293 114 327 131
rect 451 267 485 283
rect 451 61 485 131
rect 537 267 743 286
rect 571 252 709 267
rect 537 114 571 131
rect 623 199 657 215
rect 623 61 657 131
rect 845 215 879 427
rect 998 353 1014 387
rect 1048 353 1064 387
rect 709 114 743 131
rect 795 199 879 215
rect 829 181 879 199
rect 1045 267 1079 283
rect 795 114 829 131
rect 1045 61 1079 131
rect 1143 199 1177 427
rect 1265 313 1299 531
rect 1245 279 1299 313
rect 1333 267 1367 575
rect 1143 115 1177 131
rect 1247 199 1281 215
rect 1247 61 1281 131
rect 1333 115 1367 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1003 61
rect 1037 21 1139 61
rect 1173 21 1275 61
rect 1309 21 1408 61
rect 0 0 1408 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 595 1305 629 1311
rect 595 1277 629 1305
rect 731 1305 765 1311
rect 731 1277 765 1305
rect 867 1305 901 1311
rect 867 1277 901 1305
rect 1003 1305 1037 1311
rect 1003 1277 1037 1305
rect 1139 1305 1173 1311
rect 1139 1277 1173 1305
rect 1275 1305 1309 1311
rect 1275 1277 1309 1305
rect 80 501 114 535
rect 248 427 282 461
rect 80 353 114 387
rect 444 501 478 535
rect 578 501 612 535
rect 666 427 700 461
rect 1143 650 1177 684
rect 836 501 870 535
rect 932 427 966 461
rect 482 353 516 387
rect 293 279 327 313
rect 777 279 811 313
rect 1014 353 1048 387
rect 1211 279 1245 313
rect 1333 575 1367 609
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
rect 1003 27 1037 55
rect 1003 21 1037 27
rect 1139 27 1173 55
rect 1139 21 1173 27
rect 1275 27 1309 55
rect 1275 21 1309 27
<< metal1 >>
rect 0 1311 1408 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 595 1311
rect 629 1277 731 1311
rect 765 1277 867 1311
rect 901 1277 1003 1311
rect 1037 1277 1139 1311
rect 1173 1277 1275 1311
rect 1309 1277 1408 1311
rect 0 1271 1408 1277
rect 1131 684 1189 690
rect 1109 650 1143 684
rect 1177 650 1189 684
rect 1131 644 1189 650
rect 1321 609 1379 615
rect 1299 575 1333 609
rect 1367 575 1379 609
rect 1321 569 1379 575
rect 68 535 126 541
rect 432 535 490 541
rect 566 535 624 541
rect 824 535 882 541
rect 68 501 80 535
rect 114 501 444 535
rect 478 501 578 535
rect 612 502 836 535
rect 612 501 734 502
rect 812 501 836 502
rect 870 501 882 535
rect 68 495 126 501
rect 432 495 490 501
rect 566 495 624 501
rect 824 495 882 501
rect 236 461 294 467
rect 654 461 712 467
rect 920 461 978 467
rect 80 427 248 461
rect 282 427 666 461
rect 700 427 932 461
rect 966 427 978 461
rect 236 421 294 427
rect 654 421 712 427
rect 920 421 978 427
rect 68 387 126 393
rect 470 387 528 393
rect 1002 387 1060 393
rect 68 353 80 387
rect 114 353 482 387
rect 516 353 1014 387
rect 1048 353 1060 387
rect 68 347 126 353
rect 470 347 528 353
rect 1002 347 1060 353
rect 281 313 339 319
rect 765 313 823 319
rect 1199 313 1257 319
rect 281 279 293 313
rect 327 279 777 313
rect 811 279 1211 313
rect 1245 279 1257 313
rect 281 273 339 279
rect 765 273 823 279
rect 1199 273 1257 279
rect 0 55 1408 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1003 55
rect 1037 21 1139 55
rect 1173 21 1275 55
rect 1309 21 1408 55
rect 0 0 1408 21
<< labels >>
rlabel metal1 97 370 97 370 1 A
port 1 n
rlabel metal1 265 444 265 444 1 CI
port 2 n
rlabel metal1 129 518 129 518 1 B
port 3 n
rlabel metal1 1228 296 1228 296 1 CON
port 4 n
rlabel metal1 1160 667 1160 667 1 S
port 5 n
rlabel metal1 1350 592 1350 592 1 CO
port 6 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
