* File: sky130_osu_sc_12T_hs__or2_8.pex.spice
* Created: Fri Nov 12 15:12:59 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__OR2_8%GND 1 2 3 4 5 6 67 71 73 80 82 89 91 98
+ 100 107 109 117 132 134
r141 132 134 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r142 115 117 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.56 $Y2=0.755
r143 109 115 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.475
+ $Y=0.152 $X2=4.56 $Y2=0.305
r144 105 107 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.755
r145 101 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r146 96 125 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r147 96 98 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.755
r148 92 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r149 91 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r150 87 124 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r151 87 89 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r152 83 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r153 82 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r154 78 123 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r155 78 80 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r156 73 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r157 69 71 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r158 67 134 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r159 67 132 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r160 67 105 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.7 $Y2=0.305
r161 67 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.615 $Y2=0.152
r162 67 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.785 $Y2=0.152
r163 67 69 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r164 67 74 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r165 67 109 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.475 $Y2=0.152
r166 67 110 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=3.785 $Y2=0.152
r167 67 100 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r168 67 101 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r169 67 91 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r170 67 92 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r171 67 82 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r172 67 83 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r173 67 73 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r174 67 74 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r175 6 117 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.575 $X2=4.56 $Y2=0.755
r176 5 107 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.755
r177 4 98 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.7 $Y=0.575
+ $X2=2.84 $Y2=0.755
r178 3 89 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.755
r179 2 80 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.755
r180 1 71 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__OR2_8%VDD 1 2 3 4 5 49 51 60 62 68 72 78 82 88
+ 92 99 109 113
r81 109 113 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=4.42 $Y2=4.287
r82 99 102 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.56 $Y=2.955
+ $X2=4.56 $Y2=3.635
r83 97 102 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.56 $Y=4.135
+ $X2=4.56 $Y2=3.635
r84 95 113 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=4.25
+ $X2=4.42 $Y2=4.25
r85 93 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=4.287
+ $X2=3.7 $Y2=4.287
r86 93 95 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=4.287
+ $X2=4.42 $Y2=4.287
r87 92 97 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.475 $Y=4.287
+ $X2=4.56 $Y2=4.135
r88 92 95 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.475 $Y=4.287
+ $X2=4.42 $Y2=4.287
r89 88 91 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.7 $Y=2.955 $X2=3.7
+ $Y2=3.635
r90 86 107 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.7 $Y=4.135
+ $X2=3.7 $Y2=4.287
r91 86 91 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.7 $Y=4.135 $X2=3.7
+ $Y2=3.635
r92 83 105 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=4.287
+ $X2=2.84 $Y2=4.287
r93 83 85 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=4.287
+ $X2=3.06 $Y2=4.287
r94 82 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=4.287
+ $X2=3.7 $Y2=4.287
r95 82 85 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=4.287
+ $X2=3.06 $Y2=4.287
r96 78 81 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=2.955
+ $X2=2.84 $Y2=3.635
r97 76 105 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=4.135
+ $X2=2.84 $Y2=4.287
r98 76 81 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.84 $Y=4.135 $X2=2.84
+ $Y2=3.635
r99 73 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=1.98 $Y2=4.287
r100 73 75 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=2.38 $Y2=4.287
r101 72 105 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.84 $Y2=4.287
r102 72 75 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.38 $Y2=4.287
r103 68 71 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r104 66 104 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=4.287
r105 66 71 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=3.635
r106 63 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r107 63 65 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r108 62 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.287
r109 62 65 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r110 58 103 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r111 58 60 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.635
r112 53 109 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r113 53 57 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r114 51 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r115 51 57 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r116 49 95 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=4.135 $X2=4.42 $Y2=4.22
r117 49 107 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r118 49 85 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r119 49 75 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r120 49 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r121 49 57 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r122 49 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r123 5 102 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=2.605 $X2=4.56 $Y2=3.635
r124 5 99 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=2.605 $X2=4.56 $Y2=2.955
r125 4 91 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=3.635
r126 4 88 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.605 $X2=3.7 $Y2=2.955
r127 3 81 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=3.635
r128 3 78 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=2.955
r129 2 71 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r130 2 68 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r131 1 60 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__OR2_8%B 3 7 12 15 21
r28 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.48
r29 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.195
+ $X2=0.27 $Y2=2.48
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.195 $X2=0.27 $Y2=2.195
r31 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.195
+ $X2=0.475 $Y2=2.195
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=2.195
r33 5 7 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=3.235
r34 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.03
+ $X2=0.475 $Y2=2.195
r35 1 3 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=0.475 $Y=2.03
+ $X2=0.475 $Y2=0.85
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__OR2_8%A 3 7 10 14 20
c44 7 0 1.37149e-19 $X=0.905 $Y=3.235
r45 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.85
+ $X2=0.95 $Y2=2.85
r46 14 17 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=2.85
r47 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.905 $X2=0.95 $Y2=1.905
r48 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=2.07
r49 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=1.74
r50 7 12 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.07
r51 3 11 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.905 $Y=0.85
+ $X2=0.905 $Y2=1.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__OR2_8%A_27_521# 1 3 11 13 15 17 18 22 24 26 27
+ 28 29 33 35 37 38 40 44 46 48 49 51 55 58 59 61 62 64 68 70 72 73 75 79 81 83
+ 84 86 90 92 94 95 101 102 103 104 105 106 107 108 109 110 111 114 116 117 119
+ 122 126 128
c243 68 0 1.33323e-19 $X=3.485 $Y=0.85
c244 55 0 1.33323e-19 $X=3.055 $Y=0.85
c245 44 0 1.33323e-19 $X=2.625 $Y=0.85
c246 33 0 1.33323e-19 $X=2.195 $Y=0.85
c247 22 0 1.33323e-19 $X=1.765 $Y=0.85
r248 124 128 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.455
+ $X2=0.65 $Y2=1.455
r249 124 126 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.455
+ $X2=1.43 $Y2=1.455
r250 120 128 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.65 $Y2=1.455
r251 120 122 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.69 $Y2=0.755
r252 118 128 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.65 $Y2=1.455
r253 118 119 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=3.065
r254 116 119 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.15
+ $X2=0.61 $Y2=3.065
r255 116 117 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.15
+ $X2=0.345 $Y2=3.15
r256 112 117 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.235
+ $X2=0.345 $Y2=3.15
r257 112 114 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.26 $Y=3.235
+ $X2=0.26 $Y2=3.295
r258 99 126 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.455 $X2=1.43 $Y2=1.455
r259 97 99 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.455
+ $X2=1.43 $Y2=1.455
r260 96 97 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.455
+ $X2=1.37 $Y2=1.455
r261 92 94 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=4.345 $Y=2.48
+ $X2=4.345 $Y2=3.235
r262 88 90 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.345 $Y=1.29
+ $X2=4.345 $Y2=0.85
r263 87 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=2.405
+ $X2=3.915 $Y2=2.405
r264 86 92 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=2.405
+ $X2=4.345 $Y2=2.48
r265 86 87 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=2.405
+ $X2=3.99 $Y2=2.405
r266 85 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.365
+ $X2=3.915 $Y2=1.365
r267 84 88 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=1.365
+ $X2=4.345 $Y2=1.29
r268 84 85 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.365
+ $X2=3.99 $Y2=1.365
r269 81 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=2.48
+ $X2=3.915 $Y2=2.405
r270 81 83 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.915 $Y=2.48
+ $X2=3.915 $Y2=3.235
r271 77 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=1.29
+ $X2=3.915 $Y2=1.365
r272 77 79 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.915 $Y=1.29
+ $X2=3.915 $Y2=0.85
r273 76 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.405
+ $X2=3.485 $Y2=2.405
r274 75 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.405
+ $X2=3.915 $Y2=2.405
r275 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.405
+ $X2=3.56 $Y2=2.405
r276 74 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.365
+ $X2=3.485 $Y2=1.365
r277 73 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.365
+ $X2=3.915 $Y2=1.365
r278 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.365
+ $X2=3.56 $Y2=1.365
r279 70 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.48
+ $X2=3.485 $Y2=2.405
r280 70 72 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.485 $Y=2.48
+ $X2=3.485 $Y2=3.235
r281 66 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.29
+ $X2=3.485 $Y2=1.365
r282 66 68 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.485 $Y=1.29
+ $X2=3.485 $Y2=0.85
r283 65 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.405
+ $X2=3.055 $Y2=2.405
r284 64 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.405
+ $X2=3.485 $Y2=2.405
r285 64 65 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.405
+ $X2=3.13 $Y2=2.405
r286 63 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.365
+ $X2=3.055 $Y2=1.365
r287 62 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.365
+ $X2=3.485 $Y2=1.365
r288 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.365
+ $X2=3.13 $Y2=1.365
r289 59 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.48
+ $X2=3.055 $Y2=2.405
r290 59 61 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.055 $Y=2.48
+ $X2=3.055 $Y2=3.235
r291 58 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.33
+ $X2=3.055 $Y2=2.405
r292 57 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=1.365
r293 57 58 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.055 $Y=1.44
+ $X2=3.055 $Y2=2.33
r294 53 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.29
+ $X2=3.055 $Y2=1.365
r295 53 55 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.055 $Y=1.29
+ $X2=3.055 $Y2=0.85
r296 52 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.405
+ $X2=2.625 $Y2=2.405
r297 51 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.405
+ $X2=3.055 $Y2=2.405
r298 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.405
+ $X2=2.7 $Y2=2.405
r299 50 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.365
+ $X2=2.625 $Y2=1.365
r300 49 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.365
+ $X2=3.055 $Y2=1.365
r301 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.365
+ $X2=2.7 $Y2=1.365
r302 46 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=2.405
r303 46 48 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=3.235
r304 42 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.29
+ $X2=2.625 $Y2=1.365
r305 42 44 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.625 $Y=1.29
+ $X2=2.625 $Y2=0.85
r306 41 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.405
+ $X2=2.195 $Y2=2.405
r307 40 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.625 $Y2=2.405
r308 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.27 $Y2=2.405
r309 39 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.365
+ $X2=2.195 $Y2=1.365
r310 38 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.365
+ $X2=2.625 $Y2=1.365
r311 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.365
+ $X2=2.27 $Y2=1.365
r312 35 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=2.405
r313 35 37 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=3.235
r314 31 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=1.365
r315 31 33 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=0.85
r316 30 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.405
+ $X2=1.765 $Y2=2.405
r317 29 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=2.195 $Y2=2.405
r318 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=1.84 $Y2=2.405
r319 27 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=2.195 $Y2=1.365
r320 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=1.84 $Y2=1.365
r321 24 101 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=2.405
r322 24 26 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r323 20 28 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.84 $Y2=1.365
r324 20 99 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.43 $Y2=1.455
r325 20 22 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=0.85
r326 19 95 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.405
+ $X2=1.352 $Y2=2.405
r327 18 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.405
r328 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.445 $Y2=2.405
r329 17 95 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.33
+ $X2=1.352 $Y2=2.405
r330 16 97 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=1.455
r331 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=2.33
r332 13 95 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.352 $Y2=2.405
r333 13 15 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r334 9 96 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=1.455
r335 9 11 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.85
r336 3 114 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.295
r337 1 122 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__OR2_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68 76
+ 82 89 90 92 94 96 99 100 101 102 103 104 105 106 107 110 111 125
c166 110 0 1.33323e-19 $X=4.13 $Y=1.115
c167 104 0 1.33323e-19 $X=3.27 $Y=1.115
c168 101 0 2.66647e-19 $X=2.555 $Y=1
c169 89 0 1.33323e-19 $X=1.55 $Y=1.115
c170 40 0 1.37149e-19 $X=1.55 $Y=2.11
r171 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.995
+ $X2=4.13 $Y2=2.11
r172 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.115
+ $X2=4.13 $Y2=1
r173 110 111 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=4.13 $Y=1.115
+ $X2=4.13 $Y2=1.995
r174 107 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=2.11
+ $X2=3.27 $Y2=2.11
r175 106 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=2.11
+ $X2=4.13 $Y2=2.11
r176 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=2.11
+ $X2=3.415 $Y2=2.11
r177 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.995
+ $X2=3.27 $Y2=2.11
r178 104 121 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.115
+ $X2=3.27 $Y2=1
r179 104 105 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=3.27 $Y=1.115
+ $X2=3.27 $Y2=1.995
r180 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.11
+ $X2=2.41 $Y2=2.11
r181 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.11
+ $X2=3.27 $Y2=2.11
r182 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.11
+ $X2=2.555 $Y2=2.11
r183 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1
+ $X2=2.41 $Y2=1
r184 100 121 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1
+ $X2=3.27 $Y2=1
r185 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1
+ $X2=2.555 $Y2=1
r186 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.995
+ $X2=2.41 $Y2=2.11
r187 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=1
r188 98 99 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=1.995
r189 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.11
+ $X2=1.55 $Y2=2.11
r190 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.11
+ $X2=2.41 $Y2=2.11
r191 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.11
+ $X2=1.695 $Y2=2.11
r192 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1
+ $X2=1.55 $Y2=1
r193 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=2.41 $Y2=1
r194 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=1.695 $Y2=1
r195 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=2.11
r196 90 92 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=1.74
r197 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r198 89 92 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.74
r199 85 87 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.13 $Y=2.955
+ $X2=4.13 $Y2=3.635
r200 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=2.11
+ $X2=4.13 $Y2=2.11
r201 82 85 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=4.13 $Y=2.11
+ $X2=4.13 $Y2=2.955
r202 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=1 $X2=4.13
+ $Y2=1
r203 76 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.13 $Y=0.755
+ $X2=4.13 $Y2=1
r204 71 73 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=2.955
+ $X2=3.27 $Y2=3.635
r205 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.11
+ $X2=3.27 $Y2=2.11
r206 68 71 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.27 $Y=2.11
+ $X2=3.27 $Y2=2.955
r207 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1 $X2=3.27
+ $Y2=1
r208 62 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.27 $Y=0.755
+ $X2=3.27 $Y2=1
r209 57 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=2.955
+ $X2=2.41 $Y2=3.635
r210 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.11
+ $X2=2.41 $Y2=2.11
r211 54 57 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.41 $Y=2.11
+ $X2=2.41 $Y2=2.955
r212 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1 $X2=2.41
+ $Y2=1
r213 48 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.41 $Y=0.755
+ $X2=2.41 $Y2=1
r214 43 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r215 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.11
r216 40 43 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.955
r217 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r218 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r219 12 87 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.605 $X2=4.13 $Y2=3.635
r220 12 85 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.605 $X2=4.13 $Y2=2.955
r221 11 73 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=3.635
r222 11 71 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.605 $X2=3.27 $Y2=2.955
r223 10 59 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=3.635
r224 10 57 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=2.955
r225 9 45 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r226 9 43 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r227 4 76 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.755
r228 3 62 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.755
r229 2 48 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.755
r230 1 34 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
.ends

