* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_12T_ms__pcgate_1
** N=23 EP=0 IP=0 FDC=31
M0 6 SE gnd gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=-900 $Y=575 $D=9
M1 gnd E 6 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=-470 $Y=575 $D=9
M2 gnd 5 9 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=480 $Y=575 $D=9
M3 17 6 gnd gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=910 $Y=575 $D=9
M4 5 8 17 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=1270 $Y=575 $D=9
M5 18 CK 5 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=1870 $Y=575 $D=9
M6 gnd 9 18 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=2230 $Y=575 $D=9
M7 8 CK gnd gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=2660 $Y=575 $D=9
M8 gnd 9 10 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=3700 $Y=575 $D=9
M9 15 10 gnd gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=4130 $Y=575 $D=9
M10 19 10 11 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=5080 $Y=575 $D=9
M11 gnd CK 19 gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=5440 $Y=575 $D=9
M12 ECK 11 gnd gnd nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=5940 $Y=575 $D=9
M13 12 SE 6 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=-900 $Y=2605 $D=79
M14 vdd E 12 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=-540 $Y=2605 $D=79
M15 vdd 5 9 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=480 $Y=2605 $D=79
M16 13 6 vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=910 $Y=2605 $D=79
M17 5 CK 13 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=1270 $Y=2605 $D=79
M18 14 8 5 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=1870 $Y=2605 $D=79
M19 vdd 9 14 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=2230 $Y=2605 $D=79
M20 8 CK vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=2660 $Y=2605 $D=79
M21 vdd 9 10 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=3700 $Y=2605 $D=79
M22 15 10 vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=4130 $Y=2605 $D=79
M23 11 10 vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=5080 $Y=2605 $D=79
M24 vdd CK 11 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=5510 $Y=2605 $D=79
M25 ECK 11 vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=5940 $Y=2605 $D=79
X26 gnd vdd Dpar a=16.3422 p=19.99 m=1 $[nwdiode] $X=-1345 $Y=2425 $D=185
X27 20 SE Probe probetype=1 $[SE] $X=-657 $Y=2478 $D=289
X28 21 E Probe probetype=1 $[E] $X=-312 $Y=2853 $D=289
X29 22 CK Probe probetype=1 $[CK] $X=2868 $Y=1368 $D=289
X30 23 ECK Probe probetype=1 $[ECK] $X=6223 $Y=1733 $D=289
.ENDS
***************************************
