* File: sky130_osu_sc_15T_ls__buf_1.spice
* Created: Fri Nov 12 14:54:42 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__buf_1.pex.spice"
.subckt sky130_osu_sc_15T_ls__buf_1  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1002_d N_GND_M1002_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_VDD_M1001_d N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.2 A=0.3 P=4.3 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=4.38075 P=8.87
pX5_noxref noxref_6 A A PROBETYPE=1
pX6_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__buf_1.pxi.spice"
*
.ends
*
*
