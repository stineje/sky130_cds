magic
tech sky130A
magscale 1 2
timestamp 1612373228
<< nwell >>
rect -10 529 2090 1119
<< nmoslvt >>
rect 80 115 110 243
rect 272 115 302 199
rect 370 115 400 243
rect 442 115 472 243
rect 632 115 662 243
rect 704 115 734 243
rect 824 115 854 243
rect 896 115 926 243
rect 982 115 1012 243
rect 1054 115 1084 243
rect 1174 115 1204 243
rect 1246 115 1276 243
rect 1332 115 1362 243
rect 1522 115 1552 243
rect 1594 115 1624 243
rect 1692 115 1722 199
rect 1884 115 1914 243
rect 1970 115 2000 243
<< pmos >>
rect 80 565 110 965
rect 270 565 300 965
rect 356 565 386 965
rect 442 565 472 965
rect 632 565 662 965
rect 704 565 734 965
rect 824 565 854 965
rect 896 565 926 965
rect 982 565 1012 965
rect 1054 565 1084 965
rect 1174 565 1204 965
rect 1246 565 1276 965
rect 1332 565 1362 965
rect 1522 565 1552 965
rect 1608 565 1638 965
rect 1694 565 1724 965
rect 1884 565 1914 965
rect 1970 565 2000 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 163 243
rect 110 131 121 215
rect 155 131 163 215
rect 317 215 370 243
rect 317 199 325 215
rect 110 115 163 131
rect 219 165 272 199
rect 219 131 227 165
rect 261 131 272 165
rect 219 115 272 131
rect 302 131 325 199
rect 359 131 370 215
rect 302 115 370 131
rect 400 115 442 243
rect 472 215 525 243
rect 472 131 483 215
rect 517 131 525 215
rect 472 115 525 131
rect 579 215 632 243
rect 579 131 587 215
rect 621 131 632 215
rect 579 115 632 131
rect 662 115 704 243
rect 734 215 824 243
rect 734 131 745 215
rect 813 131 824 215
rect 734 115 824 131
rect 854 115 896 243
rect 926 165 982 243
rect 926 131 937 165
rect 971 131 982 165
rect 926 115 982 131
rect 1012 115 1054 243
rect 1084 215 1174 243
rect 1084 131 1095 215
rect 1163 131 1174 215
rect 1084 115 1174 131
rect 1204 115 1246 243
rect 1276 215 1332 243
rect 1276 131 1287 215
rect 1321 131 1332 215
rect 1276 115 1332 131
rect 1362 215 1415 243
rect 1362 131 1373 215
rect 1407 131 1415 215
rect 1362 115 1415 131
rect 1469 215 1522 243
rect 1469 131 1477 215
rect 1511 131 1522 215
rect 1469 115 1522 131
rect 1552 115 1594 243
rect 1624 215 1677 243
rect 1624 131 1635 215
rect 1669 199 1677 215
rect 1831 215 1884 243
rect 1669 131 1692 199
rect 1624 115 1692 131
rect 1722 165 1775 199
rect 1722 131 1733 165
rect 1767 131 1775 165
rect 1722 115 1775 131
rect 1831 131 1839 215
rect 1873 131 1884 215
rect 1831 115 1884 131
rect 1914 215 1970 243
rect 1914 131 1925 215
rect 1959 131 1970 215
rect 1914 115 1970 131
rect 2000 215 2053 243
rect 2000 131 2011 215
rect 2045 131 2053 215
rect 2000 115 2053 131
<< pdiff >>
rect 27 949 80 965
rect 27 741 35 949
rect 69 741 80 949
rect 27 565 80 741
rect 110 949 163 965
rect 110 605 121 949
rect 155 605 163 949
rect 110 565 163 605
rect 217 949 270 965
rect 217 673 225 949
rect 259 673 270 949
rect 217 565 270 673
rect 300 949 356 965
rect 300 673 311 949
rect 345 673 356 949
rect 300 565 356 673
rect 386 949 442 965
rect 386 741 397 949
rect 431 741 442 949
rect 386 565 442 741
rect 472 949 525 965
rect 472 673 483 949
rect 517 673 525 949
rect 472 565 525 673
rect 579 949 632 965
rect 579 673 587 949
rect 621 673 632 949
rect 579 565 632 673
rect 662 565 704 965
rect 734 949 824 965
rect 734 605 745 949
rect 813 605 824 949
rect 734 565 824 605
rect 854 565 896 965
rect 926 949 982 965
rect 926 673 937 949
rect 971 673 982 949
rect 926 565 982 673
rect 1012 565 1054 965
rect 1084 949 1174 965
rect 1084 673 1095 949
rect 1163 673 1174 949
rect 1084 565 1174 673
rect 1204 565 1246 965
rect 1276 949 1332 965
rect 1276 605 1287 949
rect 1321 605 1332 949
rect 1276 565 1332 605
rect 1362 949 1415 965
rect 1362 605 1373 949
rect 1407 605 1415 949
rect 1362 565 1415 605
rect 1469 949 1522 965
rect 1469 673 1477 949
rect 1511 673 1522 949
rect 1469 565 1522 673
rect 1552 949 1608 965
rect 1552 741 1563 949
rect 1597 741 1608 949
rect 1552 565 1608 741
rect 1638 949 1694 965
rect 1638 673 1649 949
rect 1683 673 1694 949
rect 1638 565 1694 673
rect 1724 949 1777 965
rect 1724 673 1735 949
rect 1769 673 1777 949
rect 1724 565 1777 673
rect 1831 949 1884 965
rect 1831 605 1839 949
rect 1873 605 1884 949
rect 1831 565 1884 605
rect 1914 949 1970 965
rect 1914 605 1925 949
rect 1959 605 1970 949
rect 1914 565 1970 605
rect 2000 949 2053 965
rect 2000 605 2011 949
rect 2045 605 2053 949
rect 2000 565 2053 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 227 131 261 165
rect 325 131 359 215
rect 483 131 517 215
rect 587 131 621 215
rect 745 131 813 215
rect 937 131 971 165
rect 1095 131 1163 215
rect 1287 131 1321 215
rect 1373 131 1407 215
rect 1477 131 1511 215
rect 1635 131 1669 215
rect 1733 131 1767 165
rect 1839 131 1873 215
rect 1925 131 1959 215
rect 2011 131 2045 215
<< pdiffc >>
rect 35 741 69 949
rect 121 605 155 949
rect 225 673 259 949
rect 311 673 345 949
rect 397 741 431 949
rect 483 673 517 949
rect 587 673 621 949
rect 745 605 813 949
rect 937 673 971 949
rect 1095 673 1163 949
rect 1287 605 1321 949
rect 1373 605 1407 949
rect 1477 673 1511 949
rect 1563 741 1597 949
rect 1649 673 1683 949
rect 1735 673 1769 949
rect 1839 605 1873 949
rect 1925 605 1959 949
rect 2011 605 2045 949
<< psubdiff >>
rect 26 27 50 61
rect 84 27 108 61
rect 162 27 186 61
rect 220 27 244 61
rect 298 27 322 61
rect 356 27 380 61
rect 434 27 458 61
rect 492 27 516 61
rect 570 27 594 61
rect 628 27 652 61
rect 706 27 730 61
rect 764 27 788 61
rect 842 27 866 61
rect 900 27 924 61
rect 978 27 1002 61
rect 1036 27 1060 61
rect 1114 27 1138 61
rect 1172 27 1196 61
rect 1250 27 1274 61
rect 1308 27 1332 61
rect 1386 27 1410 61
rect 1444 27 1468 61
rect 1522 27 1546 61
rect 1580 27 1604 61
rect 1658 27 1682 61
rect 1716 27 1740 61
rect 1794 27 1818 61
rect 1852 27 1876 61
rect 1930 27 1954 61
rect 1988 27 2012 61
<< nsubdiff >>
rect 26 1049 50 1083
rect 84 1049 108 1083
rect 162 1049 186 1083
rect 220 1049 244 1083
rect 298 1049 322 1083
rect 356 1049 380 1083
rect 434 1049 458 1083
rect 492 1049 516 1083
rect 570 1049 594 1083
rect 628 1049 652 1083
rect 706 1049 730 1083
rect 764 1049 788 1083
rect 842 1049 866 1083
rect 900 1049 924 1083
rect 978 1049 1002 1083
rect 1036 1049 1060 1083
rect 1114 1049 1138 1083
rect 1172 1049 1196 1083
rect 1250 1049 1274 1083
rect 1308 1049 1332 1083
rect 1386 1049 1410 1083
rect 1444 1049 1468 1083
rect 1522 1049 1546 1083
rect 1580 1049 1604 1083
rect 1658 1049 1682 1083
rect 1716 1049 1740 1083
rect 1794 1049 1818 1083
rect 1852 1049 1876 1083
rect 1930 1049 1954 1083
rect 1988 1049 2012 1083
<< psubdiffcont >>
rect 50 27 84 61
rect 186 27 220 61
rect 322 27 356 61
rect 458 27 492 61
rect 594 27 628 61
rect 730 27 764 61
rect 866 27 900 61
rect 1002 27 1036 61
rect 1138 27 1172 61
rect 1274 27 1308 61
rect 1410 27 1444 61
rect 1546 27 1580 61
rect 1682 27 1716 61
rect 1818 27 1852 61
rect 1954 27 1988 61
<< nsubdiffcont >>
rect 50 1049 84 1083
rect 186 1049 220 1083
rect 322 1049 356 1083
rect 458 1049 492 1083
rect 594 1049 628 1083
rect 730 1049 764 1083
rect 866 1049 900 1083
rect 1002 1049 1036 1083
rect 1138 1049 1172 1083
rect 1274 1049 1308 1083
rect 1410 1049 1444 1083
rect 1546 1049 1580 1083
rect 1682 1049 1716 1083
rect 1818 1049 1852 1083
rect 1954 1049 1988 1083
<< poly >>
rect 80 965 110 991
rect 270 965 300 991
rect 356 965 386 991
rect 442 965 472 991
rect 632 965 662 991
rect 704 965 734 991
rect 824 965 854 991
rect 896 965 926 991
rect 982 965 1012 991
rect 1054 965 1084 991
rect 1174 965 1204 991
rect 1246 965 1276 991
rect 1332 965 1362 991
rect 1522 965 1552 991
rect 1608 965 1638 991
rect 1694 965 1724 991
rect 1884 965 1914 991
rect 1970 965 2000 991
rect 80 442 110 565
rect 270 527 300 565
rect 243 497 300 527
rect 79 426 133 442
rect 79 392 89 426
rect 123 392 133 426
rect 79 376 133 392
rect 79 375 110 376
rect 80 243 110 375
rect 243 307 273 497
rect 356 455 386 565
rect 442 534 472 565
rect 432 518 486 534
rect 432 484 442 518
rect 476 484 486 518
rect 432 468 486 484
rect 315 439 386 455
rect 315 405 325 439
rect 359 425 386 439
rect 359 405 400 425
rect 315 389 400 405
rect 219 291 273 307
rect 356 303 400 389
rect 219 257 229 291
rect 263 271 273 291
rect 263 257 302 271
rect 219 241 302 257
rect 370 243 400 303
rect 442 243 472 468
rect 632 425 662 565
rect 704 534 734 565
rect 704 518 758 534
rect 704 484 714 518
rect 748 484 758 518
rect 704 468 758 484
rect 632 409 686 425
rect 824 423 854 565
rect 896 528 926 565
rect 982 528 1012 565
rect 896 518 1012 528
rect 896 484 928 518
rect 962 484 1012 518
rect 896 474 1012 484
rect 1054 423 1084 565
rect 1174 534 1204 565
rect 1150 518 1204 534
rect 1150 484 1160 518
rect 1194 484 1204 518
rect 1150 468 1204 484
rect 632 375 642 409
rect 676 375 686 409
rect 632 359 686 375
rect 728 393 1180 423
rect 632 243 662 359
rect 728 315 758 393
rect 1150 351 1180 393
rect 1246 419 1276 565
rect 1332 534 1362 565
rect 1332 518 1403 534
rect 1522 528 1552 565
rect 1332 504 1359 518
rect 1343 484 1359 504
rect 1393 484 1403 518
rect 1343 468 1403 484
rect 1486 518 1552 528
rect 1486 484 1502 518
rect 1536 484 1552 518
rect 1486 474 1552 484
rect 1246 403 1300 419
rect 1246 369 1256 403
rect 1290 369 1300 403
rect 1246 353 1300 369
rect 704 285 758 315
rect 800 335 854 351
rect 800 301 810 335
rect 844 301 854 335
rect 800 285 854 301
rect 704 243 734 285
rect 824 243 854 285
rect 896 335 1012 345
rect 896 301 928 335
rect 962 301 1012 335
rect 896 291 1012 301
rect 896 243 926 291
rect 982 243 1012 291
rect 1054 335 1108 351
rect 1054 301 1064 335
rect 1098 301 1108 335
rect 1054 285 1108 301
rect 1150 335 1204 351
rect 1150 301 1160 335
rect 1194 301 1204 335
rect 1150 285 1204 301
rect 1054 243 1084 285
rect 1174 243 1204 285
rect 1246 243 1276 353
rect 1343 315 1373 468
rect 1332 285 1373 315
rect 1486 318 1516 474
rect 1608 432 1638 565
rect 1694 527 1724 565
rect 1884 549 1914 565
rect 1694 501 1751 527
rect 1874 519 1914 549
rect 1694 497 1775 501
rect 1721 469 1775 497
rect 1576 416 1638 432
rect 1576 382 1588 416
rect 1622 382 1638 416
rect 1576 366 1638 382
rect 1486 286 1552 318
rect 1332 243 1362 285
rect 1522 243 1552 286
rect 1594 243 1624 366
rect 1745 307 1775 469
rect 1874 419 1904 519
rect 1970 460 2000 565
rect 1849 403 1904 419
rect 1849 369 1859 403
rect 1893 369 1904 403
rect 1946 444 2000 460
rect 1946 410 1956 444
rect 1990 410 2000 444
rect 1946 394 2000 410
rect 1849 353 1904 369
rect 1874 308 1904 353
rect 1745 291 1799 307
rect 1745 271 1755 291
rect 1692 257 1755 271
rect 1789 257 1799 291
rect 1874 258 1914 308
rect 272 199 302 241
rect 1692 241 1799 257
rect 1884 243 1914 258
rect 1970 243 2000 394
rect 1692 199 1722 241
rect 80 89 110 115
rect 272 89 302 115
rect 370 89 400 115
rect 442 89 472 115
rect 632 89 662 115
rect 704 89 734 115
rect 824 89 854 115
rect 896 89 926 115
rect 982 89 1012 115
rect 1054 89 1084 115
rect 1174 89 1204 115
rect 1246 89 1276 115
rect 1332 89 1362 115
rect 1522 89 1552 115
rect 1594 89 1624 115
rect 1692 89 1722 115
rect 1884 89 1914 115
rect 1970 89 2000 115
<< polycont >>
rect 89 392 123 426
rect 442 484 476 518
rect 325 405 359 439
rect 229 257 263 291
rect 714 484 748 518
rect 928 484 962 518
rect 1160 484 1194 518
rect 642 375 676 409
rect 1359 484 1393 518
rect 1502 484 1536 518
rect 1256 369 1290 403
rect 810 301 844 335
rect 928 301 962 335
rect 1064 301 1098 335
rect 1160 301 1194 335
rect 1588 382 1622 416
rect 1859 369 1893 403
rect 1956 410 1990 444
rect 1755 257 1789 291
<< locali >>
rect 0 1089 2090 1110
rect 0 1049 50 1089
rect 84 1049 186 1089
rect 220 1049 322 1089
rect 356 1049 458 1089
rect 492 1049 594 1089
rect 628 1049 730 1089
rect 764 1049 866 1089
rect 900 1049 1002 1089
rect 1036 1049 1138 1089
rect 1172 1049 1274 1089
rect 1308 1049 1410 1089
rect 1444 1049 1546 1089
rect 1580 1049 1682 1089
rect 1716 1049 1818 1089
rect 1852 1049 1954 1089
rect 1988 1049 2090 1089
rect 35 949 69 1049
rect 35 725 69 741
rect 121 949 155 965
rect 47 442 81 597
rect 121 513 155 605
rect 225 949 259 965
rect 121 479 191 513
rect 47 426 123 442
rect 47 392 89 426
rect 89 376 123 392
rect 157 291 191 479
rect 225 369 259 673
rect 311 949 345 965
rect 397 949 431 1049
rect 397 725 431 741
rect 483 949 517 965
rect 345 673 483 691
rect 311 657 517 673
rect 587 949 621 1049
rect 587 657 621 673
rect 745 949 813 965
rect 937 949 971 1049
rect 937 657 971 673
rect 1095 949 1163 965
rect 813 605 816 623
rect 745 602 816 605
rect 1095 602 1163 673
rect 442 568 816 602
rect 996 568 1163 602
rect 1287 949 1321 1049
rect 1287 589 1321 605
rect 1373 949 1407 965
rect 1477 949 1511 965
rect 1563 949 1597 1049
rect 1563 725 1597 741
rect 1649 949 1683 965
rect 1511 673 1649 691
rect 1477 657 1683 673
rect 1735 949 1769 965
rect 1373 602 1407 605
rect 1373 568 1461 602
rect 325 439 359 523
rect 442 518 476 568
rect 309 405 325 439
rect 359 405 375 439
rect 225 335 359 369
rect 121 257 229 291
rect 263 257 279 291
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 257
rect 325 215 359 301
rect 442 318 476 484
rect 714 518 748 534
rect 714 483 748 484
rect 928 518 962 534
rect 748 449 844 483
rect 642 409 676 425
rect 642 359 676 375
rect 810 335 844 449
rect 928 335 962 484
rect 442 284 776 318
rect 810 285 844 301
rect 928 285 962 301
rect 996 335 1030 568
rect 1160 518 1194 534
rect 1160 483 1194 484
rect 742 231 776 284
rect 996 251 1030 301
rect 1064 449 1160 483
rect 1359 518 1393 534
rect 1359 483 1393 484
rect 1064 335 1098 449
rect 1427 403 1461 568
rect 1240 369 1256 403
rect 1290 369 1306 403
rect 1373 369 1461 403
rect 1502 518 1536 534
rect 1373 335 1407 369
rect 1144 301 1160 335
rect 1194 301 1407 335
rect 1502 335 1536 484
rect 1570 432 1604 523
rect 1570 416 1638 432
rect 1570 382 1588 416
rect 1622 382 1638 416
rect 1735 403 1769 673
rect 1839 949 1873 965
rect 1839 557 1873 605
rect 1925 949 1959 1049
rect 1925 589 1959 605
rect 2011 949 2045 965
rect 2011 583 2045 597
rect 2011 549 2068 583
rect 1839 518 1873 523
rect 1839 484 1990 518
rect 1956 444 1990 484
rect 1672 369 1859 403
rect 1893 369 1909 403
rect 1672 347 1706 369
rect 1635 313 1706 347
rect 1956 335 1990 410
rect 1064 285 1098 301
rect 121 115 155 131
rect 227 165 261 181
rect 227 61 261 131
rect 325 115 359 131
rect 483 215 517 231
rect 483 61 517 131
rect 587 215 621 231
rect 742 215 813 231
rect 996 217 1163 251
rect 742 197 745 215
rect 587 61 621 131
rect 1095 215 1163 217
rect 745 115 813 131
rect 937 165 971 181
rect 937 61 971 131
rect 1095 115 1163 131
rect 1287 215 1321 231
rect 1287 61 1321 131
rect 1373 215 1407 301
rect 1373 115 1407 131
rect 1477 215 1511 231
rect 1477 61 1511 131
rect 1635 215 1669 313
rect 1839 301 1990 335
rect 1739 257 1755 291
rect 1789 257 1805 291
rect 1839 215 1873 301
rect 2034 268 2068 549
rect 2011 234 2068 268
rect 1635 115 1669 131
rect 1733 165 1767 181
rect 1733 61 1767 131
rect 1839 115 1873 131
rect 1925 215 1959 231
rect 1925 61 1959 131
rect 2011 215 2045 234
rect 2011 115 2045 131
rect 0 21 50 61
rect 84 21 186 61
rect 220 21 322 61
rect 356 21 458 61
rect 492 21 594 61
rect 628 21 730 61
rect 764 21 866 61
rect 900 21 1002 61
rect 1036 21 1138 61
rect 1172 21 1274 61
rect 1308 21 1410 61
rect 1444 21 1546 61
rect 1580 21 1682 61
rect 1716 21 1818 61
rect 1852 21 1954 61
rect 1988 21 2090 61
rect 0 0 2090 21
<< viali >>
rect 50 1083 84 1089
rect 50 1055 84 1083
rect 186 1083 220 1089
rect 186 1055 220 1083
rect 322 1083 356 1089
rect 322 1055 356 1083
rect 458 1083 492 1089
rect 458 1055 492 1083
rect 594 1083 628 1089
rect 594 1055 628 1083
rect 730 1083 764 1089
rect 730 1055 764 1083
rect 866 1083 900 1089
rect 866 1055 900 1083
rect 1002 1083 1036 1089
rect 1002 1055 1036 1083
rect 1138 1083 1172 1089
rect 1138 1055 1172 1083
rect 1274 1083 1308 1089
rect 1274 1055 1308 1083
rect 1410 1083 1444 1089
rect 1410 1055 1444 1083
rect 1546 1083 1580 1089
rect 1546 1055 1580 1083
rect 1682 1083 1716 1089
rect 1682 1055 1716 1083
rect 1818 1083 1852 1089
rect 1818 1055 1852 1083
rect 1954 1083 1988 1089
rect 1954 1055 1988 1083
rect 47 597 81 631
rect 325 523 359 557
rect 325 301 359 335
rect 229 257 263 261
rect 229 227 263 257
rect 714 449 748 483
rect 642 375 676 409
rect 910 301 928 335
rect 928 301 944 335
rect 996 301 1030 335
rect 1160 449 1194 483
rect 1359 449 1393 483
rect 1256 369 1290 403
rect 1570 523 1604 557
rect 2011 605 2045 631
rect 2011 597 2045 605
rect 1839 523 1873 557
rect 1859 369 1893 403
rect 1502 301 1536 335
rect 1755 257 1789 261
rect 1755 227 1789 257
rect 50 27 84 55
rect 50 21 84 27
rect 186 27 220 55
rect 186 21 220 27
rect 322 27 356 55
rect 322 21 356 27
rect 458 27 492 55
rect 458 21 492 27
rect 594 27 628 55
rect 594 21 628 27
rect 730 27 764 55
rect 730 21 764 27
rect 866 27 900 55
rect 866 21 900 27
rect 1002 27 1036 55
rect 1002 21 1036 27
rect 1138 27 1172 55
rect 1138 21 1172 27
rect 1274 27 1308 55
rect 1274 21 1308 27
rect 1410 27 1444 55
rect 1410 21 1444 27
rect 1546 27 1580 55
rect 1546 21 1580 27
rect 1682 27 1716 55
rect 1682 21 1716 27
rect 1818 27 1852 55
rect 1818 21 1852 27
rect 1954 27 1988 55
rect 1954 21 1988 27
<< metal1 >>
rect 0 1089 2090 1110
rect 0 1055 50 1089
rect 84 1055 186 1089
rect 220 1055 322 1089
rect 356 1055 458 1089
rect 492 1055 594 1089
rect 628 1055 730 1089
rect 764 1055 866 1089
rect 900 1055 1002 1089
rect 1036 1055 1138 1089
rect 1172 1055 1274 1089
rect 1308 1055 1410 1089
rect 1444 1055 1546 1089
rect 1580 1055 1682 1089
rect 1716 1055 1818 1089
rect 1852 1055 1954 1089
rect 1988 1055 2090 1089
rect 0 1049 2090 1055
rect 35 631 93 637
rect 1999 631 2057 637
rect 35 597 47 631
rect 81 597 127 631
rect 1977 597 2011 631
rect 2045 597 2057 631
rect 35 591 93 597
rect 1999 591 2057 597
rect 313 557 371 563
rect 1558 557 1616 563
rect 1827 557 1885 563
rect 313 523 325 557
rect 359 523 1570 557
rect 1604 523 1616 557
rect 1804 523 1839 557
rect 1873 523 1885 557
rect 313 517 371 523
rect 1558 517 1616 523
rect 1827 517 1885 523
rect 702 483 760 489
rect 1148 483 1206 489
rect 1347 483 1405 489
rect 702 449 714 483
rect 748 449 1160 483
rect 1194 449 1359 483
rect 1393 449 1405 483
rect 702 443 760 449
rect 1148 443 1206 449
rect 1347 443 1405 449
rect 630 409 688 415
rect 630 375 642 409
rect 676 375 710 409
rect 1244 403 1302 409
rect 1847 403 1905 409
rect 630 369 688 375
rect 1244 369 1256 403
rect 1290 369 1859 403
rect 1893 369 1905 403
rect 1244 363 1302 369
rect 1847 363 1905 369
rect 313 335 371 341
rect 898 335 956 341
rect 313 301 325 335
rect 359 301 910 335
rect 944 301 956 335
rect 313 295 371 301
rect 898 295 956 301
rect 984 335 1042 341
rect 1490 335 1548 341
rect 984 301 996 335
rect 1030 301 1502 335
rect 1536 301 1548 335
rect 984 295 1042 301
rect 1490 295 1548 301
rect 217 261 275 267
rect 1743 261 1801 267
rect 217 227 229 261
rect 263 227 1755 261
rect 1789 227 1801 261
rect 217 221 275 227
rect 1743 221 1801 227
rect 0 55 2090 61
rect 0 21 50 55
rect 84 21 186 55
rect 220 21 322 55
rect 356 21 458 55
rect 492 21 594 55
rect 628 21 730 55
rect 764 21 866 55
rect 900 21 1002 55
rect 1036 21 1138 55
rect 1172 21 1274 55
rect 1308 21 1410 55
rect 1444 21 1546 55
rect 1580 21 1682 55
rect 1716 21 1818 55
rect 1852 21 1954 55
rect 1988 21 2090 55
rect 0 0 2090 21
<< labels >>
rlabel viali 659 392 659 392 1 D
port 1 n
rlabel viali 1376 466 1376 466 1 CK
port 2 n
rlabel viali 1857 540 1857 540 1 QN
port 3 n
rlabel viali 1587 540 1587 540 1 SN
port 4 n
rlabel viali 65 614 65 614 1 RN
port 5 n
rlabel viali 2028 614 2028 614 1 Q
port 6 n
rlabel viali 67 48 67 48 1 gnd
rlabel viali 67 1062 67 1062 1 vdd
<< end >>
