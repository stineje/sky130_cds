* File: sky130_osu_sc_12T_ms__buf_1.pxi.spice
* Created: Fri Nov 12 15:21:29 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__BUF_1%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_MS__BUF_1%GND
x_PM_SKY130_OSU_SC_12T_MS__BUF_1%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_29_p
+ N_VDD_c_30_p N_VDD_c_39_p VDD N_VDD_c_31_p PM_SKY130_OSU_SC_12T_MS__BUF_1%VDD
x_PM_SKY130_OSU_SC_12T_MS__BUF_1%A N_A_M1002_g N_A_M1001_g N_A_c_54_n N_A_c_55_n
+ A PM_SKY130_OSU_SC_12T_MS__BUF_1%A
x_PM_SKY130_OSU_SC_12T_MS__BUF_1%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_c_103_n
+ N_A_27_115#_M1003_g N_A_27_115#_c_92_n N_A_27_115#_c_93_n N_A_27_115#_c_94_n
+ N_A_27_115#_c_95_n N_A_27_115#_c_98_n N_A_27_115#_c_99_n N_A_27_115#_c_101_n
+ N_A_27_115#_c_102_n PM_SKY130_OSU_SC_12T_MS__BUF_1%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__BUF_1%Y N_Y_M1000_d N_Y_M1003_d N_Y_c_144_n
+ N_Y_c_150_n Y N_Y_c_147_n N_Y_c_149_n PM_SKY130_OSU_SC_12T_MS__BUF_1%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_A_M1002_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.475 $Y2=0.835
cc_4 N_GND_c_4_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.835
cc_5 N_GND_M1002_b N_A_M1001_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_6 N_GND_M1002_b N_A_c_54_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_7 N_GND_M1002_b N_A_c_55_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_8 N_GND_M1002_b N_A_27_115#_M1000_g 0.0337861f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.835
cc_9 N_GND_c_3_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.905
+ $Y2=0.835
cc_10 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=0.835
cc_11 N_GND_M1002_b N_A_27_115#_c_92_n 0.0597491f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.38
cc_12 N_GND_M1002_b N_A_27_115#_c_93_n 0.0562401f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=1.455
cc_13 N_GND_M1002_b N_A_27_115#_c_94_n 0.0168393f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.455
cc_14 N_GND_M1002_b N_A_27_115#_c_95_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_15 N_GND_c_2_p N_A_27_115#_c_95_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_16 N_GND_c_4_p N_A_27_115#_c_95_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_17 N_GND_M1002_b N_A_27_115#_c_98_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.955
cc_18 N_GND_M1002_b N_A_27_115#_c_99_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.455
cc_19 N_GND_c_3_p N_A_27_115#_c_99_n 0.00702738f $X=0.69 $Y=0.755 $X2=0.88
+ $Y2=1.455
cc_20 N_GND_M1002_b N_A_27_115#_c_101_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.455
cc_21 N_GND_M1002_b N_A_27_115#_c_102_n 0.00663593f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.455
cc_22 N_GND_M1002_b N_Y_c_144_n 0.00875894f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.755
cc_23 N_GND_c_4_p N_Y_c_144_n 0.00471849f $X=1.02 $Y=0.19 $X2=1.12 $Y2=0.755
cc_24 N_GND_M1002_b Y 0.0164841f $X=-0.045 $Y=0 $X2=1.065 $Y2=1.795
cc_25 N_GND_M1002_b N_Y_c_147_n 0.0130304f $X=-0.045 $Y=0 $X2=1.12 $Y2=1
cc_26 N_GND_c_3_p N_Y_c_147_n 0.00125659f $X=0.69 $Y=0.755 $X2=1.12 $Y2=1
cc_27 N_GND_M1002_b N_Y_c_149_n 0.00501078f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.48
cc_28 N_VDD_M1001_b N_A_M1001_g 0.0245629f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_29 N_VDD_c_29_p N_A_M1001_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=3.235
cc_30 N_VDD_c_30_p N_A_M1001_g 0.00337744f $X=0.69 $Y=3.635 $X2=0.475 $Y2=3.235
cc_31 N_VDD_c_31_p N_A_M1001_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.235
cc_32 N_VDD_M1001_d N_A_c_55_n 0.00628533f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2
cc_33 N_VDD_M1001_b N_A_c_55_n 0.00328912f $X=-0.045 $Y=2.425 $X2=0.635 $Y2=2
cc_34 N_VDD_c_30_p N_A_c_55_n 0.00264661f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2
cc_35 N_VDD_M1001_d A 0.00797576f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2.85
cc_36 N_VDD_c_30_p A 0.00510982f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2.85
cc_37 N_VDD_M1001_b N_A_27_115#_c_103_n 0.0194495f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.53
cc_38 N_VDD_c_30_p N_A_27_115#_c_103_n 0.00337744f $X=0.69 $Y=3.635 $X2=0.905
+ $Y2=2.53
cc_39 N_VDD_c_39_p N_A_27_115#_c_103_n 0.00606474f $X=1.02 $Y=4.22 $X2=0.905
+ $Y2=2.53
cc_40 N_VDD_c_31_p N_A_27_115#_c_103_n 0.00468827f $X=1.02 $Y=4.25 $X2=0.905
+ $Y2=2.53
cc_41 N_VDD_M1001_b N_A_27_115#_c_94_n 0.0187682f $X=-0.045 $Y=2.425 $X2=1.18
+ $Y2=2.455
cc_42 N_VDD_M1001_b N_A_27_115#_c_98_n 0.00996008f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=2.955
cc_43 N_VDD_c_29_p N_A_27_115#_c_98_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=2.955
cc_44 N_VDD_c_31_p N_A_27_115#_c_98_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26
+ $Y2=2.955
cc_45 N_VDD_M1001_b N_Y_c_150_n 0.00317324f $X=-0.045 $Y=2.425 $X2=1.12 $Y2=2.48
cc_46 N_VDD_c_39_p N_Y_c_150_n 0.00736239f $X=1.02 $Y=4.22 $X2=1.12 $Y2=2.48
cc_47 N_VDD_c_31_p N_Y_c_150_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.12 $Y2=2.48
cc_48 N_VDD_M1001_b N_Y_c_149_n 0.0107503f $X=-0.045 $Y=2.425 $X2=1.12 $Y2=2.48
cc_49 A N_A_27_115#_M1001_s 0.00410657f $X=0.635 $Y=2.85 $X2=0.135 $Y2=2.605
cc_50 N_A_M1002_g N_A_27_115#_M1000_g 0.0340677f $X=0.475 $Y=0.835 $X2=0.905
+ $Y2=0.835
cc_51 A N_A_27_115#_c_103_n 0.00419145f $X=0.635 $Y=2.85 $X2=0.905 $Y2=2.53
cc_52 N_A_M1002_g N_A_27_115#_c_92_n 0.00260138f $X=0.475 $Y=0.835 $X2=1.18
+ $Y2=2.38
cc_53 N_A_M1001_g N_A_27_115#_c_92_n 0.00209773f $X=0.475 $Y=3.235 $X2=1.18
+ $Y2=2.38
cc_54 N_A_c_54_n N_A_27_115#_c_92_n 0.0139096f $X=0.635 $Y=2 $X2=1.18 $Y2=2.38
cc_55 N_A_c_55_n N_A_27_115#_c_92_n 0.00361737f $X=0.635 $Y=2 $X2=1.18 $Y2=2.38
cc_56 N_A_M1001_g N_A_27_115#_c_94_n 0.0482814f $X=0.475 $Y=3.235 $X2=1.18
+ $Y2=2.455
cc_57 N_A_c_55_n N_A_27_115#_c_94_n 0.00468272f $X=0.635 $Y=2 $X2=1.18 $Y2=2.455
cc_58 N_A_M1002_g N_A_27_115#_c_95_n 0.0124465f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.755
cc_59 N_A_M1002_g N_A_27_115#_c_98_n 0.0330322f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=2.955
cc_60 N_A_c_55_n N_A_27_115#_c_98_n 0.0548951f $X=0.635 $Y=2 $X2=0.26 $Y2=2.955
cc_61 A N_A_27_115#_c_98_n 0.0155137f $X=0.635 $Y=2.85 $X2=0.26 $Y2=2.955
cc_62 N_A_M1002_g N_A_27_115#_c_99_n 0.0207696f $X=0.475 $Y=0.835 $X2=0.88
+ $Y2=1.455
cc_63 N_A_c_54_n N_A_27_115#_c_99_n 0.00273049f $X=0.635 $Y=2 $X2=0.88 $Y2=1.455
cc_64 N_A_c_55_n N_A_27_115#_c_99_n 0.00886797f $X=0.635 $Y=2 $X2=0.88 $Y2=1.455
cc_65 N_A_M1002_g N_A_27_115#_c_102_n 6.59135e-19 $X=0.475 $Y=0.835 $X2=0.965
+ $Y2=1.455
cc_66 N_A_c_55_n N_Y_c_150_n 0.0135622f $X=0.635 $Y=2 $X2=1.12 $Y2=2.48
cc_67 A N_Y_c_150_n 0.00731851f $X=0.635 $Y=2.85 $X2=1.12 $Y2=2.48
cc_68 N_A_M1002_g Y 0.00310306f $X=0.475 $Y=0.835 $X2=1.065 $Y2=1.795
cc_69 N_A_c_54_n Y 0.00441844f $X=0.635 $Y=2 $X2=1.065 $Y2=1.795
cc_70 N_A_c_55_n Y 0.0200396f $X=0.635 $Y=2 $X2=1.065 $Y2=1.795
cc_71 N_A_M1002_g N_Y_c_147_n 7.77582e-19 $X=0.475 $Y=0.835 $X2=1.12 $Y2=1
cc_72 N_A_c_55_n N_Y_c_149_n 0.00609526f $X=0.635 $Y=2 $X2=1.12 $Y2=2.48
cc_73 N_A_27_115#_M1000_g N_Y_c_144_n 0.00356431f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_74 N_A_27_115#_c_93_n N_Y_c_144_n 0.00467107f $X=1.18 $Y=1.455 $X2=1.12
+ $Y2=0.755
cc_75 N_A_27_115#_c_102_n N_Y_c_144_n 7.29965e-19 $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=0.755
cc_76 N_A_27_115#_c_103_n N_Y_c_150_n 0.00519491f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_77 N_A_27_115#_c_94_n N_Y_c_150_n 0.0134943f $X=1.18 $Y=2.455 $X2=1.12
+ $Y2=2.48
cc_78 N_A_27_115#_M1000_g Y 0.00406656f $X=0.905 $Y=0.835 $X2=1.065 $Y2=1.795
cc_79 N_A_27_115#_c_92_n Y 0.0310322f $X=1.18 $Y=2.38 $X2=1.065 $Y2=1.795
cc_80 N_A_27_115#_c_93_n Y 0.0161039f $X=1.18 $Y=1.455 $X2=1.065 $Y2=1.795
cc_81 N_A_27_115#_c_99_n Y 8.73078e-19 $X=0.88 $Y=1.455 $X2=1.065 $Y2=1.795
cc_82 N_A_27_115#_c_102_n Y 0.0121742f $X=0.965 $Y=1.455 $X2=1.065 $Y2=1.795
cc_83 N_A_27_115#_M1000_g N_Y_c_147_n 0.00567487f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=1
cc_84 N_A_27_115#_c_93_n N_Y_c_147_n 0.0014753f $X=1.18 $Y=1.455 $X2=1.12 $Y2=1
cc_85 N_A_27_115#_c_102_n N_Y_c_147_n 0.00278861f $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=1
cc_86 N_A_27_115#_c_103_n N_Y_c_149_n 0.0015856f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_87 N_A_27_115#_c_92_n N_Y_c_149_n 0.00226191f $X=1.18 $Y=2.38 $X2=1.12
+ $Y2=2.48
cc_88 N_A_27_115#_c_94_n N_Y_c_149_n 0.00513726f $X=1.18 $Y=2.455 $X2=1.12
+ $Y2=2.48
