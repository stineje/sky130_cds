magic
tech sky130A
magscale 1 2
timestamp 1612371863
<< nwell >>
rect -9 529 462 1119
<< nmoslvt >>
rect 80 115 110 243
rect 152 115 182 243
rect 252 115 282 243
rect 324 115 354 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
rect 338 565 368 965
<< ndiff >>
rect 27 231 80 243
rect 27 131 35 231
rect 69 131 80 231
rect 27 115 80 131
rect 110 115 152 243
rect 182 231 252 243
rect 182 131 200 231
rect 234 131 252 231
rect 182 115 252 131
rect 282 115 324 243
rect 354 231 407 243
rect 354 131 365 231
rect 399 131 407 231
rect 354 115 407 131
<< pdiff >>
rect 27 949 80 965
rect 27 711 35 949
rect 69 711 80 949
rect 27 565 80 711
rect 110 949 166 965
rect 110 779 121 949
rect 155 779 166 949
rect 110 565 166 779
rect 196 949 252 965
rect 196 711 207 949
rect 241 711 252 949
rect 196 565 252 711
rect 282 881 338 965
rect 282 711 293 881
rect 327 711 338 881
rect 282 565 338 711
rect 368 949 421 965
rect 368 711 379 949
rect 413 711 421 949
rect 368 565 421 711
<< ndiffc >>
rect 35 131 69 231
rect 200 131 234 231
rect 365 131 399 231
<< pdiffc >>
rect 35 711 69 949
rect 121 779 155 949
rect 207 711 241 949
rect 293 711 327 881
rect 379 711 413 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 991
rect 338 965 368 991
rect 80 528 110 565
rect 44 518 110 528
rect 44 484 60 518
rect 94 484 110 518
rect 44 474 110 484
rect 44 318 74 474
rect 166 462 196 565
rect 152 432 196 462
rect 116 416 182 432
rect 116 382 128 416
rect 162 382 182 416
rect 116 366 182 382
rect 44 266 110 318
rect 80 243 110 266
rect 152 243 182 366
rect 252 361 282 565
rect 338 426 368 565
rect 338 410 416 426
rect 338 382 370 410
rect 224 345 282 361
rect 224 311 234 345
rect 268 311 282 345
rect 224 295 282 311
rect 252 243 282 295
rect 324 376 370 382
rect 404 376 416 410
rect 324 360 416 376
rect 324 352 368 360
rect 324 243 354 352
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
rect 324 89 354 115
<< polycont >>
rect 60 484 94 518
rect 128 382 162 416
rect 234 311 268 345
rect 370 376 404 410
<< locali >>
rect 0 1089 462 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 462 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 763 155 779
rect 207 950 413 985
rect 207 949 241 950
rect 69 711 207 729
rect 379 949 413 950
rect 35 695 241 711
rect 293 881 327 897
rect 60 518 94 597
rect 293 614 327 711
rect 379 695 413 711
rect 293 580 336 614
rect 60 468 94 484
rect 128 416 162 523
rect 128 366 162 382
rect 216 361 250 449
rect 216 345 268 361
rect 216 311 234 345
rect 234 295 268 311
rect 302 335 336 580
rect 370 410 404 426
rect 370 360 404 376
rect 35 231 69 249
rect 35 61 69 131
rect 200 115 234 131
rect 365 231 399 249
rect 365 61 399 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 462 61
rect 0 0 462 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 60 597 94 631
rect 128 523 162 557
rect 216 449 250 483
rect 370 376 404 410
rect 302 301 336 335
rect 200 231 234 261
rect 200 227 234 231
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
<< metal1 >>
rect 0 1089 462 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 462 1089
rect 0 1049 462 1055
rect 48 631 106 637
rect 48 597 60 631
rect 94 597 128 631
rect 48 591 106 597
rect 116 557 174 563
rect 116 523 128 557
rect 162 523 196 557
rect 116 517 174 523
rect 204 483 262 489
rect 182 449 216 483
rect 250 449 262 483
rect 204 443 262 449
rect 358 410 416 416
rect 336 376 370 410
rect 404 376 416 410
rect 358 370 416 376
rect 290 335 348 341
rect 290 301 302 335
rect 336 301 348 335
rect 290 295 348 301
rect 188 261 246 267
rect 304 261 338 295
rect 188 227 200 261
rect 234 227 338 261
rect 188 221 246 227
rect 0 55 462 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 462 55
rect 0 0 462 21
<< labels >>
rlabel viali 77 614 77 614 1 A0
port 1 n
rlabel viali 233 466 233 466 1 B0
port 2 n
rlabel viali 145 540 145 540 1 A1
port 4 n
rlabel viali 387 393 387 393 1 B1
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
rlabel metal1 321 268 321 268 1 Y
port 3 n
<< end >>
