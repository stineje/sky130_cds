* File: sky130_osu_sc_18T_ms__addf_1.pex.spice
* Created: Thu Oct 29 17:26:53 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%GND 1 2 3 4 5 56 60 62 72 74 81 83 96 98
+ 105 107 120 122
c182 96 0 1.91914e-19 $X=5.31 $Y=0.825
c183 72 0 1.85877e-19 $X=2.34 $Y=0.825
r184 120 122 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r185 114 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=0.152
+ $X2=6.32 $Y2=0.152
r186 107 108 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r187 103 115 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.152
r188 103 105 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.825
r189 99 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.152
+ $X2=5.31 $Y2=0.152
r190 98 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.152
+ $X2=6.32 $Y2=0.152
r191 94 113 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.152
r192 94 96 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.825
r193 84 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0.152
+ $X2=3.2 $Y2=0.152
r194 83 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=0.152
+ $X2=5.31 $Y2=0.152
r195 79 112 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.152
r196 79 81 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.825
r197 74 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.152
+ $X2=3.2 $Y2=0.152
r198 70 72 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.34 $Y=0.305
+ $X2=2.34 $Y2=0.825
r199 63 108 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r200 58 108 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r201 58 60 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r202 56 114 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.46 $Y=0.152
+ $X2=6.405 $Y2=0.152
r203 56 107 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r204 56 122 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.17
+ $X2=6.46 $Y2=0.17
r205 56 120 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r206 56 70 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.34 $Y2=0.305
r207 56 62 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.255 $Y2=0.152
r208 56 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.425 $Y2=0.152
r209 56 98 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.235 $Y2=0.152
r210 56 99 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.395 $Y2=0.152
r211 56 83 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=0.152
+ $X2=5.225 $Y2=0.152
r212 56 84 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.285 $Y2=0.152
r213 56 74 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.115 $Y2=0.152
r214 56 75 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.425 $Y2=0.152
r215 56 62 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.255 $Y2=0.152
r216 56 63 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r217 5 105 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=6.195
+ $Y=0.575 $X2=6.32 $Y2=0.825
r218 4 96 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.17
+ $Y=0.575 $X2=5.31 $Y2=0.825
r219 3 81 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.575 $X2=3.2 $Y2=0.825
r220 2 72 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.2
+ $Y=0.575 $X2=2.34 $Y2=0.825
r221 1 60 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%VDD 1 2 3 4 5 46 50 54 62 66 72 76 86 90
+ 96 100 109 114 121
r109 114 121 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=6.49
+ $X2=6.46 $Y2=6.49
r110 109 114 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=6.46 $Y2=6.507
r111 109 118 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r112 106 121 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.405 $Y=6.507
+ $X2=6.46 $Y2=6.507
r113 106 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=6.507
+ $X2=6.32 $Y2=6.507
r114 100 118 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r115 100 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r116 96 99 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.32 $Y=3.455
+ $X2=6.32 $Y2=5.835
r117 94 107 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.32 $Y=6.355
+ $X2=6.32 $Y2=6.507
r118 94 99 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.32 $Y=6.355
+ $X2=6.32 $Y2=5.835
r119 91 105 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=6.507
+ $X2=5.31 $Y2=6.507
r120 91 93 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.395 $Y=6.507
+ $X2=5.78 $Y2=6.507
r121 90 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=6.507
+ $X2=6.32 $Y2=6.507
r122 90 93 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=6.235 $Y=6.507
+ $X2=5.78 $Y2=6.507
r123 86 89 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=5.31 $Y=4.135
+ $X2=5.31 $Y2=5.835
r124 84 105 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.31 $Y=6.355
+ $X2=5.31 $Y2=6.507
r125 84 89 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.31 $Y=6.355
+ $X2=5.31 $Y2=5.835
r126 81 83 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=4.42 $Y=6.507
+ $X2=5.1 $Y2=6.507
r127 79 81 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.74 $Y=6.507
+ $X2=4.42 $Y2=6.507
r128 77 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=6.507
+ $X2=3.2 $Y2=6.507
r129 77 79 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.285 $Y=6.507
+ $X2=3.74 $Y2=6.507
r130 76 105 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.31 $Y2=6.507
r131 76 83 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.1 $Y2=6.507
r132 72 75 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=3.2 $Y=4.135
+ $X2=3.2 $Y2=5.835
r133 70 104 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.2 $Y=6.355
+ $X2=3.2 $Y2=6.507
r134 70 75 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.2 $Y=6.355
+ $X2=3.2 $Y2=5.835
r135 67 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=6.507
+ $X2=2.34 $Y2=6.507
r136 67 69 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=2.425 $Y=6.507
+ $X2=3.06 $Y2=6.507
r137 66 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=6.507
+ $X2=3.2 $Y2=6.507
r138 66 69 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.115 $Y=6.507
+ $X2=3.06 $Y2=6.507
r139 62 65 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.34 $Y=3.795
+ $X2=2.34 $Y2=5.835
r140 60 103 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.34 $Y=6.355
+ $X2=2.34 $Y2=6.507
r141 60 65 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.34 $Y=6.355
+ $X2=2.34 $Y2=5.835
r142 57 59 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r143 55 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r144 55 57 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r145 54 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=6.507
+ $X2=2.34 $Y2=6.507
r146 54 59 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=2.255 $Y=6.507
+ $X2=1.7 $Y2=6.507
r147 50 53 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r148 48 101 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r149 48 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r150 46 121 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=6.355 $X2=6.46 $Y2=6.44
r151 46 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r152 46 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r153 46 93 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=6.355 $X2=5.78 $Y2=6.44
r154 46 83 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=6.355 $X2=5.1 $Y2=6.44
r155 46 81 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r156 46 79 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r157 46 69 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r158 46 59 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r159 46 57 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r160 5 99 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=6.195
+ $Y=3.085 $X2=6.32 $Y2=5.835
r161 5 96 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=6.195
+ $Y=3.085 $X2=6.32 $Y2=3.455
r162 4 89 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=5.17
+ $Y=3.085 $X2=5.31 $Y2=5.835
r163 4 86 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=5.17
+ $Y=3.085 $X2=5.31 $Y2=4.135
r164 3 75 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.06
+ $Y=3.085 $X2=3.2 $Y2=5.835
r165 3 72 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=3.06
+ $Y=3.085 $X2=3.2 $Y2=4.135
r166 2 65 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.2
+ $Y=3.085 $X2=2.34 $Y2=5.835
r167 2 62 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=2.2
+ $Y=3.085 $X2=2.34 $Y2=3.795
r168 1 53 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r169 1 50 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%A 3 6 8 10 11 13 14 15 16 17 19 22 23 25
+ 28 31 36 38 39 40 41 42 43 45 48 52 54 55 59 60 62 63 70 71
c207 54 0 1.91914e-19 $X=5.155 $Y=1.85
c208 43 0 1.85877e-19 $X=2.64 $Y=1.85
c209 41 0 1.24216e-19 $X=0.63 $Y=1.85
c210 40 0 1.77566e-19 $X=2.35 $Y=1.85
c211 39 0 2.67871e-19 $X=5.13 $Y=2.925
c212 31 0 1.32911e-19 $X=5.095 $Y=4.585
c213 19 0 1.74961e-19 $X=2.435 $Y=2.81
c214 14 0 9.53445e-20 $X=2.36 $Y=1.76
r215 70 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.85
+ $X2=5.155 $Y2=2.015
r216 70 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.85
+ $X2=5.155 $Y2=1.685
r217 66 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.85
+ $X2=2.495 $Y2=2.015
r218 62 66 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.495 $Y=1.76
+ $X2=2.495 $Y2=1.85
r219 62 63 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.495 $Y=1.76
+ $X2=2.495 $Y2=1.685
r220 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=2.015
r221 59 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=1.685
r222 55 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.85 $X2=5.155 $Y2=1.85
r223 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.155 $Y=1.85
+ $X2=5.155 $Y2=1.85
r224 52 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.85 $X2=2.495 $Y2=1.85
r225 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.495 $Y=1.85
+ $X2=2.495 $Y2=1.85
r226 48 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.85 $X2=0.485 $Y2=1.85
r227 45 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=1.85
r228 43 51 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.64 $Y=1.85
+ $X2=2.495 $Y2=1.85
r229 42 54 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.01 $Y=1.85
+ $X2=5.155 $Y2=1.85
r230 42 43 2.28203 $w=1.7e-07 $l=2.37e-06 $layer=MET1_cond $X=5.01 $Y=1.85
+ $X2=2.64 $Y2=1.85
r231 41 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=1.85
+ $X2=0.485 $Y2=1.85
r232 40 51 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.35 $Y=1.85
+ $X2=2.495 $Y2=1.85
r233 40 41 1.65616 $w=1.7e-07 $l=1.72e-06 $layer=MET1_cond $X=2.35 $Y=1.85
+ $X2=0.63 $Y2=1.85
r234 38 39 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=5.13 $Y=2.775
+ $X2=5.13 $Y2=2.925
r235 38 72 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.165 $Y=2.775
+ $X2=5.165 $Y2=2.015
r236 35 36 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.435 $Y=2.885
+ $X2=2.555 $Y2=2.885
r237 31 39 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=5.095 $Y=4.585
+ $X2=5.095 $Y2=2.925
r238 28 71 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.095 $Y=1.075
+ $X2=5.095 $Y2=1.685
r239 23 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.555 $Y=2.96
+ $X2=2.555 $Y2=2.885
r240 23 25 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.555 $Y=2.96
+ $X2=2.555 $Y2=4.585
r241 22 63 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.555 $Y=1.075
+ $X2=2.555 $Y2=1.685
r242 19 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=2.81
+ $X2=2.435 $Y2=2.885
r243 19 67 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.435 $Y=2.81
+ $X2=2.435 $Y2=2.015
r244 16 35 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=2.885
+ $X2=2.435 $Y2=2.885
r245 16 17 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=2.885
+ $X2=2.2 $Y2=2.885
r246 14 62 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.36 $Y=1.76
+ $X2=2.495 $Y2=1.76
r247 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=1.76
+ $X2=2.2 $Y2=1.76
r248 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=2.96
+ $X2=2.2 $Y2=2.885
r249 11 13 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.125 $Y=2.96
+ $X2=2.125 $Y2=4.585
r250 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=1.685
+ $X2=2.2 $Y2=1.76
r251 8 10 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.125 $Y=1.685
+ $X2=2.125 $Y2=1.075
r252 6 61 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.015
r253 3 60 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=1.685
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%B 3 7 11 15 19 22 26 30 34 35 38 39 44
+ 45 47 49 50 51 52 55 59 65 74 75 76 80
c228 59 0 9.53445e-20 $X=2.305 $Y=2.59
c229 55 0 1.26882e-19 $X=0.485 $Y=2.59
c230 52 0 6.46001e-20 $X=3.67 $Y=2.592
r231 80 82 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.59
+ $X2=4.265 $Y2=2.755
r232 80 81 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.59
+ $X2=4.265 $Y2=2.425
r233 75 77 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.85
+ $X2=2.975 $Y2=2.015
r234 75 76 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.85
+ $X2=2.975 $Y2=1.685
r235 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.85 $X2=2.975 $Y2=1.85
r236 65 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=2.59 $X2=4.265 $Y2=2.59
r237 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.265 $Y=2.59
+ $X2=4.265 $Y2=2.59
r238 62 74 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.975 $Y=2.59
+ $X2=2.975 $Y2=1.85
r239 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=2.59
+ $X2=2.975 $Y2=2.59
r240 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.305 $Y=2.59
+ $X2=2.305 $Y2=2.59
r241 55 94 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.485 $Y=2.59
+ $X2=0.485 $Y2=2.76
r242 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=2.59
+ $X2=0.485 $Y2=2.59
r243 52 61 0.459737 $w=1.9e-07 $l=6.95999e-07 $layer=MET1_cond $X=3.67 $Y=2.592
+ $X2=2.975 $Y2=2.59
r244 51 64 0.124897 $w=2.19e-07 $l=2.05998e-07 $layer=MET1_cond $X=4.06 $Y=2.592
+ $X2=4.265 $Y2=2.59
r245 51 52 0.386904 $w=1.65e-07 $l=3.9e-07 $layer=MET1_cond $X=4.06 $Y=2.592
+ $X2=3.67 $Y2=2.592
r246 50 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.45 $Y=2.59
+ $X2=2.305 $Y2=2.59
r247 49 61 0.0970649 $w=1.9e-07 $l=1.45e-07 $layer=MET1_cond $X=2.83 $Y=2.59
+ $X2=2.975 $Y2=2.59
r248 49 50 0.365895 $w=1.7e-07 $l=3.8e-07 $layer=MET1_cond $X=2.83 $Y=2.59
+ $X2=2.45 $Y2=2.59
r249 45 54 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=2.59
+ $X2=0.485 $Y2=2.59
r250 45 47 0.0144432 $w=1.7e-07 $l=1.5e-08 $layer=MET1_cond $X=0.63 $Y=2.59
+ $X2=0.645 $Y2=2.59
r251 44 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.16 $Y=2.59
+ $X2=2.305 $Y2=2.59
r252 44 47 1.45877 $w=1.7e-07 $l=1.515e-06 $layer=MET1_cond $X=2.16 $Y=2.59
+ $X2=0.645 $Y2=2.59
r253 42 59 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.1 $Y=2.59
+ $X2=2.305 $Y2=2.59
r254 41 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=2.59
+ $X2=2.1 $Y2=2.59
r255 39 69 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.015 $Y=2.43
+ $X2=1.765 $Y2=2.43
r256 38 41 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.015 $Y=2.43
+ $X2=2.015 $Y2=2.59
r257 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=2.43 $X2=2.015 $Y2=2.43
r258 35 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.76
+ $X2=0.895 $Y2=2.925
r259 35 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.76
+ $X2=0.895 $Y2=2.595
r260 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=2.76 $X2=0.895 $Y2=2.76
r261 32 94 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=2.76
+ $X2=0.485 $Y2=2.76
r262 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.57 $Y=2.76
+ $X2=0.895 $Y2=2.76
r263 30 82 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=4.275 $Y=4.585
+ $X2=4.275 $Y2=2.755
r264 26 81 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=4.275 $Y=1.075
+ $X2=4.275 $Y2=2.425
r265 22 77 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=2.985 $Y=4.585
+ $X2=2.985 $Y2=2.015
r266 19 76 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.985 $Y=1.075
+ $X2=2.985 $Y2=1.685
r267 13 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.595
+ $X2=1.765 $Y2=2.43
r268 13 15 1020.4 $w=1.5e-07 $l=1.99e-06 $layer=POLY_cond $X=1.765 $Y=2.595
+ $X2=1.765 $Y2=4.585
r269 9 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.265
+ $X2=1.765 $Y2=2.43
r270 9 11 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=1.765 $Y=2.265
+ $X2=1.765 $Y2=1.075
r271 7 68 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.925
r272 3 67 779.404 $w=1.5e-07 $l=1.52e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.595
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%CI 3 7 11 15 19 23 27 28 32 33 34 35 37
+ 39 43 45 46 50 56
c183 33 0 3.15979e-20 $X=1.47 $Y=2.22
c184 11 0 1.47588e-19 $X=3.415 $Y=1.075
c185 7 0 1.26882e-19 $X=1.335 $Y=4.585
r186 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=2.4
+ $X2=4.745 $Y2=2.565
r187 56 57 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=2.4
+ $X2=4.745 $Y2=2.235
r188 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=2.4 $X2=4.745 $Y2=2.4
r189 50 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.22
+ $X2=1.325 $Y2=2.385
r190 50 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.22
+ $X2=1.325 $Y2=2.055
r191 46 55 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.745 $Y=2.22
+ $X2=4.745 $Y2=2.4
r192 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.745 $Y=2.22
+ $X2=4.745 $Y2=2.22
r193 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.415 $Y=2.22
+ $X2=3.415 $Y2=2.22
r194 39 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.22 $X2=1.325 $Y2=2.22
r195 37 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.325 $Y=2.22
+ $X2=1.325 $Y2=2.22
r196 35 42 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.56 $Y=2.22
+ $X2=3.415 $Y2=2.22
r197 34 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.6 $Y=2.22
+ $X2=4.745 $Y2=2.22
r198 34 35 1.0014 $w=1.7e-07 $l=1.04e-06 $layer=MET1_cond $X=4.6 $Y=2.22
+ $X2=3.56 $Y2=2.22
r199 33 37 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.47 $Y=2.22
+ $X2=1.325 $Y2=2.22
r200 32 42 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.27 $Y=2.22
+ $X2=3.415 $Y2=2.22
r201 32 33 1.73319 $w=1.7e-07 $l=1.8e-06 $layer=MET1_cond $X=3.27 $Y=2.22
+ $X2=1.47 $Y2=2.22
r202 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=2.59 $X2=3.415 $Y2=2.59
r203 25 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.415 $Y=2.505
+ $X2=3.415 $Y2=2.22
r204 25 27 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=2.505
+ $X2=3.415 $Y2=2.59
r205 23 58 1035.79 $w=1.5e-07 $l=2.02e-06 $layer=POLY_cond $X=4.685 $Y=4.585
+ $X2=4.685 $Y2=2.565
r206 19 57 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=4.685 $Y=1.075
+ $X2=4.685 $Y2=2.235
r207 13 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.755
+ $X2=3.415 $Y2=2.59
r208 13 15 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.415 $Y=2.755
+ $X2=3.415 $Y2=4.585
r209 9 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.425
+ $X2=3.415 $Y2=2.59
r210 9 11 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=3.415 $Y=2.425
+ $X2=3.415 $Y2=1.075
r211 7 52 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.385
r212 3 51 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%CON 1 2 7 9 12 16 20 24 29 32 33 38 46
+ 48 51 52 53 54 61 63 73 80
c188 73 0 1.77566e-19 $X=1.55 $Y=0.825
c189 54 0 1.47588e-19 $X=4.115 $Y=1.48
c190 46 0 1.22485e-19 $X=3.845 $Y=1.85
c191 38 0 3.15979e-20 $X=1.665 $Y=1.765
c192 33 0 1.71092e-19 $X=6.41 $Y=2.74
c193 29 0 1.74961e-19 $X=1.665 $Y=3.025
r194 65 80 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.14 $Y=1.48
+ $X2=6.41 $Y2=1.48
r195 63 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.14 $Y=1.48
+ $X2=6.14 $Y2=1.48
r196 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.97 $Y=1.48
+ $X2=3.97 $Y2=1.48
r197 57 73 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r198 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r199 54 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.115 $Y=1.48
+ $X2=3.97 $Y2=1.48
r200 53 63 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.995 $Y=1.48
+ $X2=6.14 $Y2=1.48
r201 53 54 1.81022 $w=1.7e-07 $l=1.88e-06 $layer=MET1_cond $X=5.995 $Y=1.48
+ $X2=4.115 $Y2=1.48
r202 52 56 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.48
+ $X2=1.55 $Y2=1.48
r203 51 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.825 $Y=1.48
+ $X2=3.97 $Y2=1.48
r204 51 52 2.05094 $w=1.7e-07 $l=2.13e-06 $layer=MET1_cond $X=3.825 $Y=1.48
+ $X2=1.695 $Y2=1.48
r205 49 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.97 $Y=1.765
+ $X2=3.97 $Y2=1.48
r206 48 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=1.85
+ $X2=3.97 $Y2=1.765
r207 45 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.85
+ $X2=3.97 $Y2=1.85
r208 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.85 $X2=3.845 $Y2=1.85
r209 36 57 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.55 $Y=1.68 $X2=1.55
+ $Y2=1.48
r210 35 38 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=1.765
+ $X2=1.665 $Y2=1.765
r211 35 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.765
+ $X2=1.55 $Y2=1.68
r212 33 71 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.74
+ $X2=6.442 $Y2=2.905
r213 33 70 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.74
+ $X2=6.442 $Y2=2.575
r214 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=2.74 $X2=6.41 $Y2=2.74
r215 30 80 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.565
+ $X2=6.41 $Y2=1.48
r216 30 32 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.41 $Y=1.565
+ $X2=6.41 $Y2=2.74
r217 29 40 6.89435 $w=1.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.665 $Y=3.117
+ $X2=1.55 $Y2=3.117
r218 28 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.85
+ $X2=1.665 $Y2=1.765
r219 28 29 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.665 $Y=1.85
+ $X2=1.665 $Y2=3.025
r220 24 26 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.55 $Y=3.795
+ $X2=1.55 $Y2=5.835
r221 22 40 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.55 $Y=3.21
+ $X2=1.55 $Y2=3.117
r222 22 24 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.55 $Y=3.21
+ $X2=1.55 $Y2=3.795
r223 20 71 861.447 $w=1.5e-07 $l=1.68e-06 $layer=POLY_cond $X=6.535 $Y=4.585
+ $X2=6.535 $Y2=2.905
r224 16 70 769.149 $w=1.5e-07 $l=1.5e-06 $layer=POLY_cond $X=6.535 $Y=1.075
+ $X2=6.535 $Y2=2.575
r225 10 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=2.015
+ $X2=3.845 $Y2=1.85
r226 10 12 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=3.845 $Y=2.015
+ $X2=3.845 $Y2=4.585
r227 7 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.685
+ $X2=3.845 $Y2=1.85
r228 7 9 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.845 $Y=1.685
+ $X2=3.845 $Y2=1.075
r229 2 26 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r230 2 24 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.795
r231 1 73 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%A_784_115# 1 2 9 13 16 17 18 19 22 24 28
+ 31 33 37 39 42
c125 42 0 3.07391e-19 $X=5.585 $Y=2.755
c126 37 0 1.48211e-20 $X=4.31 $Y=0.99
c127 33 0 9.63581e-20 $X=5.415 $Y=3.25
c128 16 0 6.46001e-20 $X=3.845 $Y=3.03
c129 13 0 1.71513e-19 $X=5.585 $Y=4.585
c130 9 0 1.71092e-19 $X=5.585 $Y=1.075
r131 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.585
+ $Y=2.755 $X2=5.585 $Y2=2.755
r132 39 41 7.30282 $w=2.84e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=2.755
+ $X2=5.585 $Y2=2.755
r133 35 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.06 $Y=0.99
+ $X2=4.31 $Y2=0.99
r134 32 39 3.73949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=2.92
+ $X2=5.415 $Y2=2.755
r135 32 33 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.415 $Y=2.92
+ $X2=5.415 $Y2=3.25
r136 30 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=1.075
+ $X2=4.31 $Y2=0.99
r137 30 31 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=4.31 $Y=1.075
+ $X2=4.31 $Y2=2.135
r138 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.33 $Y=3.335
+ $X2=5.415 $Y2=3.25
r139 28 29 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=5.33 $Y=3.335
+ $X2=4.145 $Y2=3.335
r140 24 26 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.06 $Y=3.795
+ $X2=4.06 $Y2=5.835
r141 22 29 5.48216 $w=2.66e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=3.42
+ $X2=4.145 $Y2=3.335
r142 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.06 $Y=3.42
+ $X2=4.06 $Y2=3.795
r143 19 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=0.905
+ $X2=4.06 $Y2=0.99
r144 19 21 5.74118 $w=1.7e-07 $l=8e-08 $layer=LI1_cond $X=4.06 $Y=0.905 $X2=4.06
+ $Y2=0.825
r145 17 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.225 $Y=2.22
+ $X2=4.31 $Y2=2.135
r146 17 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.225 $Y=2.22
+ $X2=3.93 $Y2=2.22
r147 16 29 15.5724 $w=2.66e-07 $l=4.29564e-07 $layer=LI1_cond $X=3.845 $Y=3.03
+ $X2=4.145 $Y2=3.335
r148 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=2.305
+ $X2=3.93 $Y2=2.22
r149 15 16 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.845 $Y=2.305
+ $X2=3.845 $Y2=3.03
r150 11 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.92
+ $X2=5.585 $Y2=2.755
r151 11 13 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=5.585 $Y=2.92
+ $X2=5.585 $Y2=4.585
r152 7 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.59
+ $X2=5.585 $Y2=2.755
r153 7 9 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=5.585 $Y=2.59
+ $X2=5.585 $Y2=1.075
r154 2 26 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.92
+ $Y=3.085 $X2=4.06 $Y2=5.835
r155 2 24 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=3.92
+ $Y=3.085 $X2=4.06 $Y2=3.795
r156 1 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.575 $X2=4.06 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%A_27_617# 1 2 9 13 17
r13 17 19 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r14 15 17 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.12 $Y=3.545
+ $X2=1.12 $Y2=3.795
r15 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.46
+ $X2=1.12 $Y2=3.545
r16 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.46
+ $X2=0.345 $Y2=3.46
r17 9 11 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.26 $Y=3.795
+ $X2=0.26 $Y2=5.835
r18 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.545
+ $X2=0.345 $Y2=3.46
r19 7 9 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.26 $Y=3.545 $X2=0.26
+ $Y2=3.795
r20 2 19 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r21 2 17 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r22 1 11 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r23 1 9 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%A_526_617# 1 2 9 13 17
r12 17 19 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=3.63 $Y=3.795
+ $X2=3.63 $Y2=5.835
r13 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.63 $Y=3.54
+ $X2=3.63 $Y2=3.795
r14 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=3.455
+ $X2=3.63 $Y2=3.54
r15 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=3.455
+ $X2=2.855 $Y2=3.455
r16 9 11 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.77 $Y=3.795
+ $X2=2.77 $Y2=5.835
r17 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=3.54
+ $X2=2.855 $Y2=3.455
r18 7 9 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.77 $Y=3.54 $X2=2.77
+ $Y2=3.795
r19 2 19 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.49
+ $Y=3.085 $X2=3.63 $Y2=5.835
r20 2 17 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=3.49
+ $Y=3.085 $X2=3.63 $Y2=3.795
r21 1 11 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.63
+ $Y=3.085 $X2=2.77 $Y2=5.835
r22 1 9 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=2.63
+ $Y=3.085 $X2=2.77 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%S 1 2 9 12 15 20 23 29
c49 23 0 1.32911e-19 $X=5.8 $Y=3.335
c50 20 0 1.41304e-19 $X=5.925 $Y=3.25
c51 15 0 1.66087e-19 $X=5.925 $Y=2.22
r52 29 31 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=5.8 $Y=3.795
+ $X2=5.8 $Y2=5.835
r53 25 29 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.8 $Y=3.335 $X2=5.8
+ $Y2=3.795
r54 23 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.8 $Y=3.335 $X2=5.8
+ $Y2=3.335
r55 17 20 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=3.25
+ $X2=5.925 $Y2=3.25
r56 17 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=3.25 $X2=5.8
+ $Y2=3.335
r57 13 15 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=2.22
+ $X2=5.925 $Y2=2.22
r58 12 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=3.165
+ $X2=5.925 $Y2=3.25
r59 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=2.305
+ $X2=5.925 $Y2=2.22
r60 11 12 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.925 $Y=2.305
+ $X2=5.925 $Y2=3.165
r61 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.135 $X2=5.8
+ $Y2=2.22
r62 7 9 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=5.8 $Y=2.135 $X2=5.8
+ $Y2=0.825
r63 2 31 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=5.66
+ $Y=3.085 $X2=5.8 $Y2=5.835
r64 2 29 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=5.66
+ $Y=3.085 $X2=5.8 $Y2=3.795
r65 1 9 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=5.66
+ $Y=0.575 $X2=5.8 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%CO 1 2 8 13
r15 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.75 $Y=3.455
+ $X2=6.75 $Y2=5.835
r16 10 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.75 $Y=2.96
+ $X2=6.75 $Y2=3.455
r17 10 13 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=6.75 $Y=2.96
+ $X2=6.75 $Y2=0.825
r18 8 10 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.75 $Y=2.96 $X2=6.75
+ $Y2=2.96
r19 2 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.61
+ $Y=3.085 $X2=6.75 $Y2=5.835
r20 2 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.61
+ $Y=3.085 $X2=6.75 $Y2=3.455
r21 1 13 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.61
+ $Y=0.575 $X2=6.75 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%A_27_115# 1 2 9 11 12 15
c21 12 0 1.24216e-19 $X=0.345 $Y=1.345
r22 13 15 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.12 $Y=1.26
+ $X2=1.12 $Y2=0.825
r23 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.345
+ $X2=1.12 $Y2=1.26
r24 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.345
+ $X2=0.345 $Y2=1.345
r25 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.26
+ $X2=0.345 $Y2=1.345
r26 7 9 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=1.26 $X2=0.26
+ $Y2=0.825
r27 2 15 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r28 1 9 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__ADDF_1%A_526_115# 1 2 9 11 12 15
c33 11 0 1.07664e-19 $X=3.545 $Y=1.345
r34 13 15 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.63 $Y=1.26
+ $X2=3.63 $Y2=0.825
r35 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=1.345
+ $X2=3.63 $Y2=1.26
r36 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=1.345
+ $X2=2.855 $Y2=1.345
r37 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.26
+ $X2=2.855 $Y2=1.345
r38 7 9 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.77 $Y=1.26 $X2=2.77
+ $Y2=0.825
r39 2 15 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.49
+ $Y=0.575 $X2=3.63 $Y2=0.825
r40 1 9 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.63
+ $Y=0.575 $X2=2.77 $Y2=0.825
.ends

