* File: sky130_osu_sc_12T_hs__dff_l.spice
* Created: Fri Nov 12 15:09:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__dff_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__dff_l  GND VDD D CK ON Q
* 
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1009 N_GND_M1009_d N_A_75_248#_M1009_g N_A_32_115#_M1009_s N_GND_M1009_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1008 A_201_115# N_D_M1008_g N_GND_M1009_d N_GND_M1009_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1025 N_A_75_248#_M1025_d N_A_243_89#_M1025_g A_201_115# N_GND_M1009_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75001 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1020 A_393_115# N_CK_M1020_g N_A_75_248#_M1025_d N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.6 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1014 N_GND_M1014_d N_A_32_115#_M1014_g A_393_115# N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.9 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1016 A_551_115# N_A_32_115#_M1016_g N_GND_M1014_d N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75002.4 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1013 N_A_623_115#_M1013_d N_CK_M1013_g A_551_115# N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1005 A_743_115# N_A_243_89#_M1005_g N_A_623_115#_M1013_d N_GND_M1009_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75003.3 SB=75001 A=0.0825 P=1.4 MULT=1
MM1000 N_GND_M1000_d N_A_785_89#_M1000_g A_743_115# N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75003.7 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1001 N_A_243_89#_M1001_d N_CK_M1001_g N_GND_M1000_d N_GND_M1009_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75004.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1010 N_A_785_89#_M1010_d N_A_623_115#_M1010_g N_GND_M1010_s N_GND_M1009_b
+ NLOWVT L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1011 N_GND_M1011_d N_A_785_89#_M1011_g N_ON_M1011_s N_GND_M1009_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_Q_M1002_d N_ON_M1002_g N_GND_M1011_d N_GND_M1009_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1022 N_VDD_M1022_d N_A_75_248#_M1022_g N_A_32_115#_M1022_s N_VDD_M1022_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1021 A_201_521# N_D_M1021_g N_VDD_M1022_d N_VDD_M1022_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1015 N_A_75_248#_M1015_d N_CK_M1015_g A_201_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1012 A_393_521# N_A_243_89#_M1012_g N_A_75_248#_M1015_d N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.6 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_32_115#_M1004_g A_393_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 A_551_521# N_A_32_115#_M1006_g N_VDD_M1004_d N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_623_115#_M1003_d N_A_243_89#_M1003_g A_551_521# N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.7 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1019 A_743_521# N_CK_M1019_g N_A_623_115#_M1003_d N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75003.3 SB=75001 A=0.189 P=2.82 MULT=1
MM1017 N_VDD_M1017_d N_A_785_89#_M1017_g A_743_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_A_243_89#_M1018_d N_CK_M1018_g N_VDD_M1017_d N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1024 N_A_785_89#_M1024_d N_A_623_115#_M1024_g N_VDD_M1024_s N_VDD_M1022_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_VDD_M1007_d N_A_785_89#_M1007_g N_ON_M1007_s N_VDD_M1022_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_Q_M1023_d N_ON_M1023_g N_VDD_M1007_d N_VDD_M1022_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX26_noxref N_GND_M1009_b N_VDD_M1022_b NWDIODE A=15.0895 P=18.77
pX27_noxref noxref_20 D D PROBETYPE=1
pX28_noxref noxref_21 CK CK PROBETYPE=1
pX29_noxref noxref_22 ON ON PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
c_1323 A_551_521# 0 1.57671e-19 $X=2.755 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dff_l.pxi.spice"
*
.ends
*
*
