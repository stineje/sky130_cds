* File: sky130_osu_sc_15T_hs__addh_1.spice
* Created: Fri Nov 12 14:26:25 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_hs__addh_1.pex.spice"
.subckt sky130_osu_sc_15T_hs__addh_1  GND VDD CON B A S CO
* 
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_CON_M1006_g N_S_M1006_s N_GND_M1006_b NLOWVT L=0.15
+ W=0.64 AD=0.1088 AS=0.1696 PD=0.98 PS=1.81 NRD=11.244 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1007 A_208_115# N_B_M1007_g N_GND_M1006_d N_GND_M1006_b NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1088 PD=0.85 PS=0.98 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_208_565#_M1008_d N_A_M1008_g A_208_115# N_GND_M1006_b NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75001 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_GND_M1001_d N_A_208_565#_M1001_g N_CO_M1001_s N_GND_M1006_b NLOWVT
+ L=0.15 W=0.84 AD=0.1428 AS=0.2226 PD=1.18 PS=2.21 NRD=8.568 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_A_570_115#_M1010_d N_A_208_565#_M1010_g N_GND_M1001_d N_GND_M1006_b
+ NLOWVT L=0.15 W=0.84 AD=0.1176 AS=0.1428 PD=1.12 PS=1.18 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_CON_M1004_d N_B_M1004_g N_A_570_115#_M1010_d N_GND_M1006_b NLOWVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.1 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_A_570_115#_M1005_d N_A_M1005_g N_CON_M1004_d N_GND_M1006_b NLOWVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VDD_M1009_d N_CON_M1009_g N_S_M1009_s N_VDD_M1009_b PSHORT L=0.15 W=2
+ AD=0.34 AS=0.53 PD=2.34 PS=4.53 NRD=5.8903 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001.6 A=0.3 P=4.3 MULT=1
MM1011 N_A_208_565#_M1011_d N_B_M1011_g N_VDD_M1009_d N_VDD_M1009_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.34 PD=2.28 PS=2.34 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.7 SB=75001.1 A=0.3 P=4.3 MULT=1
MM1012 N_VDD_M1012_d N_A_M1012_g N_A_208_565#_M1011_d N_VDD_M1009_b PSHORT
+ L=0.15 W=2 AD=0.34 AS=0.28 PD=2.34 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001.1 SB=75000.7 A=0.3 P=4.3 MULT=1
MM1002 N_CO_M1002_d N_A_208_565#_M1002_g N_VDD_M1012_d N_VDD_M1009_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.34 PD=4.53 PS=2.34 NRD=0 NRS=5.8903 M=1 R=13.3333
+ SA=75001.6 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1003 N_VDD_M1003_d N_A_208_565#_M1003_g N_CON_M1003_s N_VDD_M1009_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75001 A=0.3 P=4.3 MULT=1
MM1013 A_668_565# N_B_M1013_g N_VDD_M1003_d N_VDD_M1009_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1000 N_CON_M1000_d N_A_M1000_g A_668_565# N_VDD_M1009_b PSHORT L=0.15 W=2
+ AD=0.56 AS=0.21 PD=4.56 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX14_noxref N_GND_M1006_b N_VDD_M1009_b NWDIODE A=12.4785 P=14.36
pX15_noxref noxref_12 S S PROBETYPE=1
pX16_noxref noxref_13 CO CO PROBETYPE=1
pX17_noxref noxref_14 B B PROBETYPE=1
pX18_noxref noxref_15 CON CON PROBETYPE=1
pX19_noxref noxref_16 A A PROBETYPE=1
*
.include "sky130_osu_sc_15T_hs__addh_1.pxi.spice"
*
.ends
*
*
