* File: sky130_osu_sc_15T_hs__nand2_1.pex.spice
* Created: Fri Nov 12 14:31:41 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__NAND2_1%GND 1 17 19 26 33 36
r26 33 36 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r27 24 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.865
r28 17 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r29 17 24 4.26217 $w=1.7e-07 $l=2.14243e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=1.05 $Y2=0.305
r30 17 19 3.29607 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=0.965 $Y2=0.152
r31 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r32 1 26 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NAND2_1%VDD 1 2 17 21 25 32 39 42
r20 39 42 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r21 32 35 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=3.545
+ $X2=1.12 $Y2=4.565
r22 30 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r23 28 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r24 26 37 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r25 26 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r26 25 30 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.245
r27 25 28 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r28 21 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r29 19 37 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r30 19 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r31 17 28 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r32 17 37 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r33 2 35 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r34 2 32 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.545
r35 1 24 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r36 1 21 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NAND2_1%A 3 7 10 14 20
r31 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r32 14 17 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.32 $Y=2.425
+ $X2=0.32 $Y2=3.07
r33 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.425 $X2=0.32 $Y2=2.425
r34 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.425
+ $X2=0.367 $Y2=2.59
r35 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.425
+ $X2=0.367 $Y2=2.26
r36 7 12 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.59
r37 3 11 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NAND2_1%B 3 7 10 14 19 22
c38 3 0 1.57512e-19 $X=0.835 $Y=0.895
r39 17 19 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.915 $Y=1.96
+ $X2=1.06 $Y2=1.96
r40 14 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.06 $Y=2.7 $X2=1.06
+ $Y2=2.7
r41 12 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=2.045
+ $X2=1.06 $Y2=1.96
r42 12 14 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.06 $Y=2.045
+ $X2=1.06 $Y2=2.7
r43 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=1.96 $X2=0.915 $Y2=1.96
r44 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=1.795
r45 5 10 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.125
+ $X2=0.905 $Y2=1.96
r46 5 7 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=0.905 $Y=2.125
+ $X2=0.905 $Y2=3.825
r47 3 11 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.835 $Y=0.895
+ $X2=0.835 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__NAND2_1%Y 1 3 10 16 23 24 28 34
c42 24 0 1.57512e-19 $X=0.405 $Y=1.22
r43 26 34 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.215
+ $X2=0.69 $Y2=2.33
r44 26 28 0.12036 $w=1.7e-07 $l=1.25e-07 $layer=MET1_cond $X=0.69 $Y=2.215
+ $X2=0.69 $Y2=2.09
r45 25 28 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=0.69 $Y=1.305
+ $X2=0.69 $Y2=2.09
r46 24 31 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=1.22
+ $X2=0.26 $Y2=1.22
r47 23 25 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=1.22
+ $X2=0.69 $Y2=1.305
r48 23 24 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=1.22
+ $X2=0.405 $Y2=1.22
r49 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r50 16 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.33
+ $X2=0.69 $Y2=2.33
r51 16 19 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.69 $Y=2.33
+ $X2=0.69 $Y2=3.205
r52 13 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.22
+ $X2=0.26 $Y2=1.22
r53 10 13 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.26 $Y=0.865
+ $X2=0.26 $Y2=1.22
r54 3 21 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r55 3 19 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r56 1 10 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

