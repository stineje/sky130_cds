* File: sky130_osu_sc_18T_ls__addh_1.pex.spice
* Created: Thu Oct 29 17:33:25 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%GND 1 2 31 35 37 50 52 60 62
r94 60 62 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r95 54 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r96 52 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r97 48 55 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r98 48 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.825
r99 38 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r100 37 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r101 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r102 33 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.825
r103 31 54 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r104 31 52 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r105 31 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.17
+ $X2=3.74 $Y2=0.17
r106 31 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r107 31 37 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r108 31 38 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r109 2 50 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.825
r110 1 35 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%VDD 1 2 3 28 32 36 42 46 54 58 65 70 77
r57 70 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=6.49
+ $X2=3.74 $Y2=6.49
r58 65 70 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.74 $Y2=6.507
r59 65 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r60 61 77 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.74 $Y2=6.507
r61 61 63 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.05 $Y2=6.507
r62 58 74 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.34 $Y2=6.507
r63 58 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.75 $Y2=6.507
r64 54 57 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.05 $Y=3.455
+ $X2=3.05 $Y2=5.835
r65 52 63 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=6.507
r66 52 57 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=5.835
r67 49 51 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=6.507
+ $X2=2.38 $Y2=6.507
r68 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.61 $Y2=6.507
r69 47 49 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.7 $Y2=6.507
r70 46 63 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=3.05 $Y2=6.507
r71 46 51 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=2.38 $Y2=6.507
r72 42 45 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.61 $Y=3.795
+ $X2=1.61 $Y2=5.835
r73 40 60 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=6.507
r74 40 45 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=5.835
r75 37 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=0.75 $Y2=6.507
r76 37 39 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=1.02 $Y2=6.507
r77 36 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.61 $Y2=6.507
r78 36 39 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.02 $Y2=6.507
r79 32 35 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.75 $Y=3.455
+ $X2=0.75 $Y2=5.835
r80 30 59 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=6.507
r81 30 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=5.835
r82 28 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r83 28 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r84 28 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r85 28 51 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r86 28 49 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r87 28 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r88 3 57 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=5.835
r89 3 54 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=3.455
r90 2 45 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=5.835
r91 2 42 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=3.795
r92 1 35 150 $w=1.7e-07 $l=2.84825e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.75 $Y2=5.835
r93 1 32 150 $w=1.7e-07 $l=4.59238e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.75 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%CON 1 2 3 12 15 17 18 21 25 27 29 31 35
+ 39 40 41 44 47 51 57 58
c128 51 0 2.7119e-19 $X=3.42 $Y=1.85
c129 41 0 1.57622e-19 $X=0.78 $Y=1.85
c130 29 0 1.92558e-19 $X=3.42 $Y=1.765
r131 57 59 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=2.015
r132 57 58 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=1.685
r133 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.85 $X2=0.35 $Y2=1.85
r134 51 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.85
+ $X2=3.42 $Y2=1.85
r135 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.85
+ $X2=2.62 $Y2=1.85
r136 44 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.635 $Y=1.85
+ $X2=0.35 $Y2=1.85
r137 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.85
+ $X2=0.635 $Y2=1.85
r138 41 43 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.85
+ $X2=0.635 $Y2=1.85
r139 40 47 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=2.62 $Y2=1.85
r140 40 41 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=0.78 $Y2=1.85
r141 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.84 $Y=3.455
+ $X2=3.84 $Y2=5.835
r142 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.84 $Y=3.035
+ $X2=3.84 $Y2=3.455
r143 29 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.85
r144 29 31 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.165
r145 28 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.95
+ $X2=2.62 $Y2=2.95
r146 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=3.84 $Y2=3.035
r147 27 28 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=2.705 $Y2=2.95
r148 26 48 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.85
+ $X2=2.62 $Y2=1.85
r149 25 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=3.42 $Y2=1.85
r150 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=2.705 $Y2=1.85
r151 21 23 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.62 $Y=3.455
+ $X2=2.62 $Y2=5.835
r152 19 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=2.95
r153 19 21 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=3.455
r154 18 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.865
+ $X2=2.62 $Y2=2.95
r155 17 48 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=1.85
r156 17 18 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=2.865
r157 15 59 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.015
r158 12 58 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=1.685
r159 3 37 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=5.835
r160 3 35 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=3.455
r161 2 23 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=5.835
r162 2 21 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=3.455
r163 1 31 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=1.165
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%B 3 7 11 15 21 23 26 27 28 33 38
c101 38 0 1.42567e-19 $X=3.205 $Y=2.22
c102 33 0 1.57622e-19 $X=0.905 $Y=2.22
c103 28 0 4.99902e-20 $X=3.21 $Y=2.22
r104 38 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.385
r105 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.385
r106 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.055
r107 27 28 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.06 $Y=2.22
+ $X2=3.205 $Y2=2.22
r108 26 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=2.22 $X2=3.205 $Y2=2.22
r109 26 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.22
r110 23 27 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=2.222
+ $X2=3.06 $Y2=2.222
r111 21 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=2.22 $X2=0.905 $Y2=2.22
r112 20 23 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=2.22
+ $X2=1.05 $Y2=2.22
r113 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.22
r114 15 39 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=3.265 $Y=4.585
+ $X2=3.265 $Y2=2.385
r115 9 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=2.22
r116 9 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=1.075
r117 7 35 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.965 $Y=4.585
+ $X2=0.965 $Y2=2.385
r118 3 34 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.965 $Y=1.075
+ $X2=0.965 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%A 3 7 11 15 21 23 25 26 28 33 38
c87 38 0 1.74252e-19 $X=3.685 $Y=2.59
r88 38 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.755
r89 38 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.425
r90 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.755
r91 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.425
r92 28 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.59 $X2=3.685 $Y2=2.59
r93 25 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.59
r94 25 26 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.59
+ $X2=3.54 $Y2=2.59
r95 23 26 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.587
+ $X2=3.54 $Y2=2.587
r96 21 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.59 $X2=1.385 $Y2=2.59
r97 20 23 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.59
+ $X2=1.53 $Y2=2.59
r98 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.59
r99 15 39 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=3.635 $Y=1.075
+ $X2=3.635 $Y2=2.425
r100 11 40 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.625 $Y=4.585
+ $X2=3.625 $Y2=2.755
r101 7 35 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=1.395 $Y=4.585
+ $X2=1.395 $Y2=2.755
r102 3 34 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=1.325 $Y=1.075
+ $X2=1.325 $Y2=2.425
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%A_208_617# 1 2 8 11 13 15 19 21 25 29 31
+ 32 35 39 40 43 46 48 52
c113 29 0 2.52869e-20 $X=2.835 $Y=4.585
c114 21 0 9.69384e-20 $X=2.7 $Y=1.8
r115 51 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.955
+ $X2=1.825 $Y2=2.12
r116 51 52 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.955
+ $X2=1.825 $Y2=1.8
r117 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.955 $X2=1.825 $Y2=1.955
r118 48 50 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.955
+ $X2=1.825 $Y2=1.955
r119 47 48 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.955
+ $X2=1.725 $Y2=1.955
r120 45 48 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=1.955
r121 45 46 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=2.925
r122 41 47 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=1.955
r123 41 43 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=0.825
r124 39 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.725 $Y2=2.925
r125 39 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.265 $Y2=3.01
r126 35 37 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.18 $Y=3.795
+ $X2=1.18 $Y2=5.835
r127 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.265 $Y2=3.01
r128 33 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.18 $Y2=3.795
r129 27 29 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=2.835 $Y=2.745
+ $X2=2.835 $Y2=4.585
r130 23 25 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=1.075
r131 22 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.8
+ $X2=2.285 $Y2=1.8
r132 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.8
+ $X2=2.775 $Y2=1.725
r133 21 22 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.8 $X2=2.36
+ $Y2=1.8
r134 17 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=1.8
r135 17 19 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=1.075
r136 16 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.67
+ $X2=1.885 $Y2=2.67
r137 15 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.67
+ $X2=2.835 $Y2=2.745
r138 15 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.67 $X2=1.96
+ $Y2=2.67
r139 14 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.8
+ $X2=1.825 $Y2=1.8
r140 13 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=2.285 $Y2=1.8
r141 13 14 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=1.96 $Y2=1.8
r142 9 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=2.67
r143 9 11 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=4.585
r144 8 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.67
r145 8 55 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.12
r146 2 37 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=5.835
r147 2 35 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=3.795
r148 1 43 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%S 1 2 10 13 17 18 21
r32 18 29 163.428 $w=1.68e-07 $l=2.505e-06 $layer=LI1_cond $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=5.835
r33 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=3.33
r34 14 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.26 $Y=1.475
+ $X2=0.26 $Y2=0.825
r35 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.475
+ $X2=0.26 $Y2=1.475
r36 8 17 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=3.33
r37 8 10 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=2.385
r38 7 13 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=1.475
r39 7 10 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=2.385
r40 2 29 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r41 2 18 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r42 1 21 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%CO 1 2 9 13 21 24 26 29
c51 26 0 2.52869e-20 $X=2.175 $Y=2.96
r52 26 30 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=3.045
r53 26 29 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=2.875
r54 24 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.96
+ $X2=2.175 $Y2=2.96
r55 17 21 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=1.472
r56 17 29 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=2.875
r57 13 15 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.1 $Y=3.455
+ $X2=2.1 $Y2=5.835
r58 13 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.1 $Y=3.455 $X2=2.1
+ $Y2=3.045
r59 7 21 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.472
+ $X2=2.175 $Y2=1.472
r60 7 9 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.07 $Y=1.385 $X2=2.07
+ $Y2=0.825
r61 2 15 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.96
+ $Y=3.085 $X2=2.1 $Y2=5.835
r62 2 13 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.96
+ $Y=3.085 $X2=2.1 $Y2=3.455
r63 1 9 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_1%A_570_115# 1 2 9 11 12
r11 13 15 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.85 $Y=0.72
+ $X2=3.85 $Y2=0.825
r12 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.85 $Y2=0.72
r13 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.075 $Y2=0.635
r14 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.72
+ $X2=3.075 $Y2=0.635
r15 7 9 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.72 $X2=2.99
+ $Y2=0.825
r16 2 15 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.825
r17 1 9 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.825
.ends

