magic
tech sky130A
magscale 1 2
timestamp 1606864597
<< checkpaint >>
rect -1209 -1243 1345 2575
<< nwell >>
rect -9 581 199 1341
<< nmos >>
rect 80 115 110 263
<< pmoshvt >>
rect 80 817 110 1217
<< ndiff >>
rect 27 199 80 263
rect 27 131 35 199
rect 69 131 80 199
rect 27 115 80 131
rect 110 199 163 263
rect 110 131 121 199
rect 155 131 163 199
rect 110 115 163 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 929 35 1201
rect 69 929 80 1201
rect 27 817 80 929
rect 110 1201 163 1217
rect 110 929 121 1201
rect 155 929 163 1201
rect 110 817 163 929
<< ndiffc >>
rect 35 131 69 199
rect 121 131 155 199
<< pdiffc >>
rect 35 929 69 1201
rect 121 929 155 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1271 85 1305
<< poly >>
rect 80 1217 110 1243
rect 80 494 110 817
rect 80 478 134 494
rect 80 444 90 478
rect 124 444 134 478
rect 80 428 134 444
rect 80 263 110 428
rect 80 89 110 115
<< polycont >>
rect 90 444 124 478
<< locali >>
rect 0 1311 198 1332
rect 0 1271 51 1311
rect 85 1271 198 1311
rect 35 1201 69 1271
rect 35 913 69 929
rect 121 1201 155 1217
rect 47 478 81 649
rect 121 609 155 929
rect 47 444 90 478
rect 124 444 140 478
rect 35 199 69 215
rect 35 61 69 131
rect 121 199 155 279
rect 121 115 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 47 649 81 683
rect 121 575 155 609
rect 121 279 155 313
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1311 198 1332
rect 0 1277 51 1311
rect 85 1277 198 1311
rect 0 1271 198 1277
rect 35 683 93 689
rect 35 649 47 683
rect 81 649 127 683
rect 35 643 93 649
rect 109 609 167 615
rect 109 575 121 609
rect 155 575 167 609
rect 109 569 167 575
rect 121 319 155 569
rect 109 313 167 319
rect 109 279 121 313
rect 155 279 167 313
rect 109 273 167 279
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel metal1 64 666 64 666 1 A
port 1 n
rlabel metal1 151 441 151 441 1 Y
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
