* File: sky130_osu_sc_12T_ls__tbufi_l.pxi.spice
* Created: Fri Nov 12 15:40:22 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__TBUFI_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_3_p
+ N_GND_c_4_p GND N_GND_c_5_p PM_SKY130_OSU_SC_12T_LS__TBUFI_L%GND
x_PM_SKY130_OSU_SC_12T_LS__TBUFI_L%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_38_p
+ N_VDD_c_39_p N_VDD_c_45_p VDD N_VDD_c_40_p
+ PM_SKY130_OSU_SC_12T_LS__TBUFI_L%VDD
x_PM_SKY130_OSU_SC_12T_LS__TBUFI_L%OE N_OE_c_61_n N_OE_M1002_g N_OE_c_75_n
+ N_OE_M1001_g N_OE_M1000_g N_OE_c_69_n N_OE_c_70_n N_OE_c_72_n N_OE_c_73_n OE
+ PM_SKY130_OSU_SC_12T_LS__TBUFI_L%OE
x_PM_SKY130_OSU_SC_12T_LS__TBUFI_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1003_g N_A_27_115#_c_124_n
+ N_A_27_115#_c_125_n N_A_27_115#_c_128_n N_A_27_115#_c_129_n
+ N_A_27_115#_c_130_n N_A_27_115#_c_131_n
+ PM_SKY130_OSU_SC_12T_LS__TBUFI_L%A_27_115#
x_PM_SKY130_OSU_SC_12T_LS__TBUFI_L%A N_A_M1004_g N_A_M1005_g N_A_c_179_n
+ N_A_c_180_n N_A_c_181_n A PM_SKY130_OSU_SC_12T_LS__TBUFI_L%A
x_PM_SKY130_OSU_SC_12T_LS__TBUFI_L%Y N_Y_M1004_d N_Y_M1005_d N_Y_c_223_n
+ N_Y_c_225_n Y N_Y_c_227_n N_Y_c_228_n PM_SKY130_OSU_SC_12T_LS__TBUFI_L%Y
cc_1 N_GND_M1002_b N_OE_c_61_n 0.0680263f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.75
cc_2 N_GND_M1002_b N_OE_M1002_g 0.0473001f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.755
cc_3 N_GND_c_3_p N_OE_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.755
cc_4 N_GND_c_4_p N_OE_M1002_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.755
cc_5 N_GND_c_5_p N_OE_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.755
cc_6 N_GND_M1002_b N_OE_M1000_g 0.04636f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.755
cc_7 N_GND_c_4_p N_OE_M1000_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.755
cc_8 N_GND_c_5_p N_OE_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=0.755
cc_9 N_GND_M1002_b N_OE_c_69_n 0.0094682f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.825
cc_10 N_GND_M1002_b N_OE_c_70_n 0.0555158f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.74
cc_11 N_GND_c_4_p N_OE_c_70_n 0.00277624f $X=0.69 $Y=0.74 $X2=0.69 $Y2=1.74
cc_12 N_GND_M1002_b N_OE_c_72_n 0.0025915f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.74
cc_13 N_GND_M1002_b N_OE_c_73_n 6.32202e-19 $X=-0.045 $Y=0 $X2=0.69 $Y2=1.74
cc_14 N_GND_M1002_b OE 0.0132975f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.48
cc_15 N_GND_M1002_b N_A_27_115#_M1003_g 0.0144187f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=3.445
cc_16 N_GND_M1002_b N_A_27_115#_c_124_n 0.0326306f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=2.37
cc_17 N_GND_M1002_b N_A_27_115#_c_125_n 0.0560297f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_18 N_GND_c_3_p N_A_27_115#_c_125_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_19 N_GND_c_5_p N_A_27_115#_c_125_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_20 N_GND_M1002_b N_A_27_115#_c_128_n 0.0116459f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.275
cc_21 N_GND_M1002_b N_A_27_115#_c_129_n 0.0100002f $X=-0.045 $Y=0 $X2=0.715
+ $Y2=2.37
cc_22 N_GND_M1002_b N_A_27_115#_c_130_n 0.00665288f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.37
cc_23 N_GND_M1002_b N_A_27_115#_c_131_n 0.00261804f $X=-0.045 $Y=0 $X2=0.8
+ $Y2=2.37
cc_24 N_GND_M1002_b N_A_M1004_g 0.0747634f $X=-0.045 $Y=0 $X2=1.265 $Y2=0.755
cc_25 N_GND_c_5_p N_A_M1004_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.265 $Y2=0.755
cc_26 N_GND_M1002_b N_A_M1005_g 0.0372976f $X=-0.045 $Y=0 $X2=1.265 $Y2=3.445
cc_27 N_GND_M1002_b N_A_c_179_n 0.0369358f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.98
cc_28 N_GND_M1002_b N_A_c_180_n 0.00592636f $X=-0.045 $Y=0 $X2=1.14 $Y2=2.85
cc_29 N_GND_M1002_b N_A_c_181_n 0.00983127f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.98
cc_30 N_GND_M1002_b A 0.00325554f $X=-0.045 $Y=0 $X2=1.14 $Y2=2.85
cc_31 N_GND_M1002_b N_Y_c_223_n 0.0330276f $X=-0.045 $Y=0 $X2=1.48 $Y2=0.74
cc_32 N_GND_c_5_p N_Y_c_223_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.48 $Y2=0.74
cc_33 N_GND_M1002_b N_Y_c_225_n 0.0150859f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.48
cc_34 N_GND_M1002_b Y 0.0383474f $X=-0.045 $Y=0 $X2=1.525 $Y2=1.71
cc_35 N_GND_M1002_b N_Y_c_227_n 0.0157993f $X=-0.045 $Y=0 $X2=1.48 $Y2=1.37
cc_36 N_GND_M1002_b N_Y_c_228_n 0.0157299f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.48
cc_37 N_VDD_M1001_b N_OE_c_75_n 0.0214886f $X=-0.045 $Y=2.795 $X2=0.475 $Y2=2.9
cc_38 N_VDD_c_38_p N_OE_c_75_n 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=2.9
cc_39 N_VDD_c_39_p N_OE_c_75_n 0.00354579f $X=0.69 $Y=3.275 $X2=0.475 $Y2=2.9
cc_40 N_VDD_c_40_p N_OE_c_75_n 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=2.9
cc_41 N_VDD_M1001_b N_OE_c_69_n 0.015858f $X=-0.045 $Y=2.795 $X2=0.475 $Y2=2.825
cc_42 N_VDD_c_39_p OE 0.00511329f $X=0.69 $Y=3.275 $X2=0.69 $Y2=2.48
cc_43 N_VDD_M1001_b N_A_27_115#_M1003_g 0.0215533f $X=-0.045 $Y=2.795 $X2=0.905
+ $Y2=3.445
cc_44 N_VDD_c_39_p N_A_27_115#_M1003_g 0.00354579f $X=0.69 $Y=3.275 $X2=0.905
+ $Y2=3.445
cc_45 N_VDD_c_45_p N_A_27_115#_M1003_g 0.00606474f $X=1.02 $Y=4.22 $X2=0.905
+ $Y2=3.445
cc_46 N_VDD_c_40_p N_A_27_115#_M1003_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.905
+ $Y2=3.445
cc_47 N_VDD_c_39_p N_A_27_115#_c_124_n 0.00108454f $X=0.69 $Y=3.275 $X2=0.905
+ $Y2=2.37
cc_48 N_VDD_M1001_b N_A_27_115#_c_128_n 0.0104218f $X=-0.045 $Y=2.795 $X2=0.26
+ $Y2=3.275
cc_49 N_VDD_c_38_p N_A_27_115#_c_128_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=3.275
cc_50 N_VDD_c_40_p N_A_27_115#_c_128_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26
+ $Y2=3.275
cc_51 N_VDD_c_39_p N_A_27_115#_c_129_n 0.0018576f $X=0.69 $Y=3.275 $X2=0.715
+ $Y2=2.37
cc_52 N_VDD_c_39_p N_A_27_115#_c_131_n 0.00113537f $X=0.69 $Y=3.275 $X2=0.8
+ $Y2=2.37
cc_53 N_VDD_M1001_b N_A_M1005_g 0.0254661f $X=-0.045 $Y=2.795 $X2=1.265
+ $Y2=3.445
cc_54 N_VDD_c_45_p N_A_M1005_g 0.00606474f $X=1.02 $Y=4.22 $X2=1.265 $Y2=3.445
cc_55 N_VDD_c_40_p N_A_M1005_g 0.00468827f $X=1.02 $Y=4.25 $X2=1.265 $Y2=3.445
cc_56 N_VDD_M1001_b N_A_c_180_n 0.00352748f $X=-0.045 $Y=2.795 $X2=1.14 $Y2=2.85
cc_57 N_VDD_M1001_b A 0.00824251f $X=-0.045 $Y=2.795 $X2=1.14 $Y2=2.85
cc_58 N_VDD_M1001_b N_Y_c_225_n 0.0120833f $X=-0.045 $Y=2.795 $X2=1.48 $Y2=2.48
cc_59 N_VDD_c_45_p N_Y_c_225_n 0.00757793f $X=1.02 $Y=4.22 $X2=1.48 $Y2=2.48
cc_60 N_VDD_c_40_p N_Y_c_225_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.48 $Y2=2.48
cc_61 N_OE_c_61_n N_A_27_115#_M1003_g 0.00310233f $X=0.27 $Y=2.75 $X2=0.905
+ $Y2=3.445
cc_62 N_OE_c_69_n N_A_27_115#_M1003_g 0.0207125f $X=0.475 $Y=2.825 $X2=0.905
+ $Y2=3.445
cc_63 OE N_A_27_115#_M1003_g 0.0035347f $X=0.69 $Y=2.48 $X2=0.905 $Y2=3.445
cc_64 N_OE_c_61_n N_A_27_115#_c_124_n 0.0126749f $X=0.27 $Y=2.75 $X2=0.905
+ $Y2=2.37
cc_65 N_OE_c_70_n N_A_27_115#_c_124_n 0.0119465f $X=0.69 $Y=1.74 $X2=0.905
+ $Y2=2.37
cc_66 N_OE_c_72_n N_A_27_115#_c_124_n 4.88301e-19 $X=0.69 $Y=1.74 $X2=0.905
+ $Y2=2.37
cc_67 OE N_A_27_115#_c_124_n 0.00530013f $X=0.69 $Y=2.48 $X2=0.905 $Y2=2.37
cc_68 N_OE_c_61_n N_A_27_115#_c_125_n 0.0232517f $X=0.27 $Y=2.75 $X2=0.26
+ $Y2=0.74
cc_69 N_OE_M1002_g N_A_27_115#_c_125_n 0.0234423f $X=0.475 $Y=0.755 $X2=0.26
+ $Y2=0.74
cc_70 N_OE_c_70_n N_A_27_115#_c_125_n 0.0135784f $X=0.69 $Y=1.74 $X2=0.26
+ $Y2=0.74
cc_71 N_OE_c_72_n N_A_27_115#_c_125_n 0.0116068f $X=0.69 $Y=1.74 $X2=0.26
+ $Y2=0.74
cc_72 N_OE_c_73_n N_A_27_115#_c_125_n 0.00367353f $X=0.69 $Y=1.74 $X2=0.26
+ $Y2=0.74
cc_73 OE N_A_27_115#_c_125_n 0.015341f $X=0.69 $Y=2.48 $X2=0.26 $Y2=0.74
cc_74 N_OE_c_61_n N_A_27_115#_c_128_n 0.0119128f $X=0.27 $Y=2.75 $X2=0.26
+ $Y2=3.275
cc_75 N_OE_c_75_n N_A_27_115#_c_128_n 0.00691971f $X=0.475 $Y=2.9 $X2=0.26
+ $Y2=3.275
cc_76 N_OE_c_69_n N_A_27_115#_c_128_n 0.00937784f $X=0.475 $Y=2.825 $X2=0.26
+ $Y2=3.275
cc_77 OE N_A_27_115#_c_128_n 0.00515602f $X=0.69 $Y=2.48 $X2=0.26 $Y2=3.275
cc_78 N_OE_c_69_n N_A_27_115#_c_129_n 0.00705846f $X=0.475 $Y=2.825 $X2=0.715
+ $Y2=2.37
cc_79 N_OE_c_70_n N_A_27_115#_c_129_n 0.00292172f $X=0.69 $Y=1.74 $X2=0.715
+ $Y2=2.37
cc_80 N_OE_c_72_n N_A_27_115#_c_129_n 0.00456286f $X=0.69 $Y=1.74 $X2=0.715
+ $Y2=2.37
cc_81 N_OE_c_73_n N_A_27_115#_c_129_n 5.35002e-19 $X=0.69 $Y=1.74 $X2=0.715
+ $Y2=2.37
cc_82 OE N_A_27_115#_c_129_n 0.0132193f $X=0.69 $Y=2.48 $X2=0.715 $Y2=2.37
cc_83 N_OE_c_61_n N_A_27_115#_c_130_n 0.00700951f $X=0.27 $Y=2.75 $X2=0.26
+ $Y2=2.37
cc_84 N_OE_c_61_n N_A_27_115#_c_131_n 7.28522e-19 $X=0.27 $Y=2.75 $X2=0.8
+ $Y2=2.37
cc_85 N_OE_c_70_n N_A_27_115#_c_131_n 7.06691e-19 $X=0.69 $Y=1.74 $X2=0.8
+ $Y2=2.37
cc_86 N_OE_c_72_n N_A_27_115#_c_131_n 0.00365965f $X=0.69 $Y=1.74 $X2=0.8
+ $Y2=2.37
cc_87 N_OE_c_73_n N_A_27_115#_c_131_n 5.50959e-19 $X=0.69 $Y=1.74 $X2=0.8
+ $Y2=2.37
cc_88 OE N_A_27_115#_c_131_n 0.0147957f $X=0.69 $Y=2.48 $X2=0.8 $Y2=2.37
cc_89 N_OE_M1000_g N_A_M1004_g 0.0777378f $X=0.905 $Y=0.755 $X2=1.265 $Y2=0.755
cc_90 N_OE_c_70_n N_A_M1004_g 0.00693622f $X=0.69 $Y=1.74 $X2=1.265 $Y2=0.755
cc_91 N_OE_c_72_n N_A_M1004_g 0.00287993f $X=0.69 $Y=1.74 $X2=1.265 $Y2=0.755
cc_92 OE N_A_c_179_n 2.30744e-19 $X=0.69 $Y=2.48 $X2=1.325 $Y2=1.98
cc_93 OE N_A_c_180_n 0.0100867f $X=0.69 $Y=2.48 $X2=1.14 $Y2=2.85
cc_94 N_OE_c_70_n N_A_c_181_n 2.20759e-19 $X=0.69 $Y=1.74 $X2=1.325 $Y2=1.98
cc_95 OE N_A_c_181_n 0.00765298f $X=0.69 $Y=2.48 $X2=1.325 $Y2=1.98
cc_96 N_OE_c_69_n A 9.14085e-19 $X=0.475 $Y=2.825 $X2=1.14 $Y2=2.85
cc_97 OE A 0.004991f $X=0.69 $Y=2.48 $X2=1.14 $Y2=2.85
cc_98 N_OE_c_70_n Y 2.15427e-19 $X=0.69 $Y=1.74 $X2=1.525 $Y2=1.71
cc_99 N_OE_c_72_n Y 0.00375884f $X=0.69 $Y=1.74 $X2=1.525 $Y2=1.71
cc_100 N_OE_c_73_n Y 0.0105247f $X=0.69 $Y=1.74 $X2=1.525 $Y2=1.71
cc_101 N_OE_M1000_g N_Y_c_227_n 0.00101819f $X=0.905 $Y=0.755 $X2=1.48 $Y2=1.37
cc_102 OE N_Y_c_228_n 0.013635f $X=0.69 $Y=2.48 $X2=1.48 $Y2=2.48
cc_103 N_A_27_115#_c_124_n N_A_M1005_g 0.107584f $X=0.905 $Y=2.37 $X2=1.265
+ $Y2=3.445
cc_104 N_A_27_115#_c_131_n N_A_M1005_g 3.3797e-19 $X=0.8 $Y=2.37 $X2=1.265
+ $Y2=3.445
cc_105 N_A_27_115#_c_124_n N_A_c_180_n 0.0103346f $X=0.905 $Y=2.37 $X2=1.14
+ $Y2=2.85
cc_106 N_A_27_115#_c_131_n N_A_c_180_n 0.0207737f $X=0.8 $Y=2.37 $X2=1.14
+ $Y2=2.85
cc_107 N_A_27_115#_M1003_g A 0.01062f $X=0.905 $Y=3.445 $X2=1.14 $Y2=2.85
cc_108 N_A_27_115#_c_128_n A 0.00493371f $X=0.26 $Y=3.275 $X2=1.14 $Y2=2.85
cc_109 N_A_M1004_g N_Y_c_223_n 0.0190376f $X=1.265 $Y=0.755 $X2=1.48 $Y2=0.74
cc_110 N_A_c_179_n N_Y_c_223_n 8.70049e-19 $X=1.325 $Y=1.98 $X2=1.48 $Y2=0.74
cc_111 N_A_c_181_n N_Y_c_223_n 0.00231567f $X=1.325 $Y=1.98 $X2=1.48 $Y2=0.74
cc_112 N_A_M1005_g N_Y_c_225_n 0.0168059f $X=1.265 $Y=3.445 $X2=1.48 $Y2=2.48
cc_113 N_A_c_179_n N_Y_c_225_n 0.00102058f $X=1.325 $Y=1.98 $X2=1.48 $Y2=2.48
cc_114 N_A_c_180_n N_Y_c_225_n 0.0348659f $X=1.14 $Y=2.85 $X2=1.48 $Y2=2.48
cc_115 N_A_c_181_n N_Y_c_225_n 0.00330615f $X=1.325 $Y=1.98 $X2=1.48 $Y2=2.48
cc_116 A N_Y_c_225_n 0.00706656f $X=1.14 $Y=2.85 $X2=1.48 $Y2=2.48
cc_117 N_A_M1004_g Y 0.00631192f $X=1.265 $Y=0.755 $X2=1.525 $Y2=1.71
cc_118 N_A_M1005_g Y 0.00511826f $X=1.265 $Y=3.445 $X2=1.525 $Y2=1.71
cc_119 N_A_c_179_n Y 0.0051471f $X=1.325 $Y=1.98 $X2=1.525 $Y2=1.71
cc_120 N_A_c_180_n Y 0.012418f $X=1.14 $Y=2.85 $X2=1.525 $Y2=1.71
cc_121 N_A_c_181_n Y 0.0167787f $X=1.325 $Y=1.98 $X2=1.525 $Y2=1.71
cc_122 N_A_M1004_g N_Y_c_227_n 0.00707709f $X=1.265 $Y=0.755 $X2=1.48 $Y2=1.37
cc_123 N_A_c_179_n N_Y_c_227_n 0.00129509f $X=1.325 $Y=1.98 $X2=1.48 $Y2=1.37
cc_124 N_A_c_181_n N_Y_c_227_n 0.00203451f $X=1.325 $Y=1.98 $X2=1.48 $Y2=1.37
cc_125 N_A_M1005_g N_Y_c_228_n 0.00423438f $X=1.265 $Y=3.445 $X2=1.48 $Y2=2.48
cc_126 N_A_c_179_n N_Y_c_228_n 0.00138163f $X=1.325 $Y=1.98 $X2=1.48 $Y2=2.48
cc_127 N_A_c_180_n N_Y_c_228_n 0.0027663f $X=1.14 $Y=2.85 $X2=1.48 $Y2=2.48
cc_128 N_A_c_181_n N_Y_c_228_n 0.00227834f $X=1.325 $Y=1.98 $X2=1.48 $Y2=2.48
