* File: sky130_osu_sc_18T_ms__dff_1.spice
* Created: Thu Oct 29 17:28:47 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ms__dff_1.pex.spice"
.subckt sky130_osu_sc_18T_ms__dff_1  GND VDD D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_A_75_344#_M1006_g N_A_32_115#_M1006_s N_GND_M1006_b
+ NSHORT L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1004 A_201_115# N_D_M1004_g N_GND_M1006_d N_GND_M1006_b NSHORT L=0.15 W=1
+ AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1020 N_A_75_344#_M1020_d N_A_243_89#_M1020_g A_201_115# N_GND_M1006_b NSHORT
+ L=0.15 W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1
+ R=6.66667 SA=75001 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1018 A_393_115# N_CK_M1018_g N_A_75_344#_M1020_d N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.6 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1014 N_GND_M1014_d N_A_32_115#_M1014_g A_393_115# N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.9
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1016 A_551_115# N_A_32_115#_M1016_g N_GND_M1014_d N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1012 N_A_623_115#_M1012_d N_CK_M1012_g A_551_115# N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1 R=6.66667
+ SA=75002.7 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1002 A_743_115# N_A_243_89#_M1002_g N_A_623_115#_M1012_d N_GND_M1006_b NSHORT
+ L=0.15 W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1
+ R=6.66667 SA=75003.3 SB=75001 A=0.15 P=2.3 MULT=1
MM1022 N_GND_M1022_d N_A_785_89#_M1022_g A_743_115# N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75003.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1024 N_A_243_89#_M1024_d N_CK_M1024_g N_GND_M1022_d N_GND_M1006_b NSHORT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75004.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1008 N_A_785_89#_M1008_d N_A_623_115#_M1008_g N_GND_M1008_s N_GND_M1006_b
+ NSHORT L=0.15 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1010 N_GND_M1010_d N_A_785_89#_M1010_g N_QN_M1010_s N_GND_M1006_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1025 N_Q_M1025_d N_QN_M1025_g N_GND_M1010_d N_GND_M1006_b NSHORT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_VDD_M1007_d N_A_75_344#_M1007_g N_A_32_115#_M1007_s N_VDD_M1007_b
+ PSHORT L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20
+ SA=75000.2 SB=75004.1 A=0.45 P=6.3 MULT=1
MM1005 A_201_617# N_D_M1005_g N_VDD_M1007_d N_VDD_M1007_b PSHORT L=0.15 W=3
+ AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.6
+ SB=75003.7 A=0.45 P=6.3 MULT=1
MM1021 N_A_75_344#_M1021_d N_CK_M1021_g A_201_617# N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20 SA=75001
+ SB=75003.3 A=0.45 P=6.3 MULT=1
MM1019 A_393_617# N_A_243_89#_M1019_g N_A_75_344#_M1021_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75001.6 SB=75002.7 A=0.45 P=6.3 MULT=1
MM1015 N_VDD_M1015_d N_A_32_115#_M1015_g A_393_617# N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.9
+ SB=75002.4 A=0.45 P=6.3 MULT=1
MM1017 A_551_617# N_A_32_115#_M1017_g N_VDD_M1015_d N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75002.4
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1013 N_A_623_115#_M1013_d N_A_243_89#_M1013_g A_551_617# N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75002.7 SB=75001.6 A=0.45 P=6.3 MULT=1
MM1003 A_743_617# N_CK_M1003_g N_A_623_115#_M1013_d N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75003.3 SB=75001 A=0.45 P=6.3 MULT=1
MM1023 N_VDD_M1023_d N_A_785_89#_M1023_g A_743_617# N_VDD_M1007_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75003.7
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1000 N_A_243_89#_M1000_d N_CK_M1000_g N_VDD_M1023_d N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75004.1
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1009 N_A_785_89#_M1009_d N_A_623_115#_M1009_g N_VDD_M1009_s N_VDD_M1007_b
+ PSHORT L=0.15 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20
+ SA=75000.2 SB=75000.2 A=0.45 P=6.3 MULT=1
MM1011 N_VDD_M1011_d N_A_785_89#_M1011_g N_QN_M1011_s N_VDD_M1007_b PSHORT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1001 N_Q_M1001_d N_QN_M1001_g N_VDD_M1011_d N_VDD_M1007_b PSHORT L=0.15 W=3
+ AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX26_noxref N_GND_M1006_b N_VDD_M1007_b NWDIODE A=27.835 P=22.25
pX27_noxref noxref_20 D D PROBETYPE=1
pX28_noxref noxref_21 CK CK PROBETYPE=1
pX29_noxref noxref_22 QN QN PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
c_1226 A_551_617# 0 1.57671e-19 $X=2.755 $Y=3.085
*
.include "sky130_osu_sc_18T_ms__dff_1.pxi.spice"
*
.ends
*
*
