* File: sky130_osu_sc_18T_ls__ant.pex.spice
* Created: Fri Nov 12 14:14:14 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__ANT%GND 7 10 17 20
r16 17 20 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=0.19
+ $X2=0.495 $Y2=0.24
r17 10 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r18 7 10 0.369697 $w=9.88e-07 $l=3e-08 $layer=LI1_cond $X=0.495 $Y=0.22
+ $X2=0.495 $Y2=0.19
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ANT%VDD 1 9 11 18 23
r7 23 26 0.0066304 $w=9.9e-07 $l=5e-08 $layer=MET1_cond $X=0.495 $Y=6.42
+ $X2=0.495 $Y2=6.47
r8 18 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r9 16 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r10 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r11 11 16 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.355
r12 11 13 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r13 9 13 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r14 1 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r15 1 18 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ANT%A 1 5 15 19 22 27 30 33 37 41 46 49 51
r23 46 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.59
+ $X2=0.32 $Y2=2.59
r24 43 46 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.26 $Y=2.59 $X2=0.32
+ $Y2=2.59
r25 39 41 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.69 $Y=1.915
+ $X2=0.69 $Y2=0.825
r26 38 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.26
+ $Y2=2
r27 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=2
+ $X2=0.69 $Y2=1.915
r28 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=2 $X2=0.345
+ $Y2=2
r29 33 35 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r30 31 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=2.59
r31 31 33 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=3.455
r32 30 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.505
+ $X2=0.26 $Y2=2.59
r33 29 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2
r34 29 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2.505
r35 25 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.915
+ $X2=0.26 $Y2=2
r36 25 27 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.26 $Y=1.915
+ $X2=0.26 $Y2=0.825
r37 22 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.59 $X2=0.32 $Y2=2.59
r38 22 24 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=2.59
+ $X2=0.362 $Y2=2.755
r39 22 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=2.59
+ $X2=0.362 $Y2=2.425
r40 19 24 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.755
r41 15 23 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.425
r42 5 35 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r43 5 33 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r44 1 41 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
r45 1 27 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

