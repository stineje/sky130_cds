* File: sky130_osu_sc_12T_ms__xor2_l.pxi.spice
* Created: Fri Nov 12 15:27:44 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%GND N_GND_M1005_d N_GND_M1009_d N_GND_M1005_b
+ N_GND_c_9_p N_GND_c_2_p N_GND_c_3_p N_GND_c_39_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_MS__XOR2_L%GND
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%VDD N_VDD_M1001_d N_VDD_M1004_d N_VDD_M1001_b
+ N_VDD_c_73_p N_VDD_c_78_p N_VDD_c_69_p N_VDD_c_100_p N_VDD_c_96_p VDD
+ N_VDD_c_70_p PM_SKY130_OSU_SC_12T_MS__XOR2_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_M1003_g
+ N_A_27_115#_c_117_n N_A_27_115#_c_119_n N_A_27_115#_c_120_n
+ N_A_27_115#_c_123_n N_A_27_115#_c_124_n N_A_27_115#_c_125_n
+ N_A_27_115#_c_126_n PM_SKY130_OSU_SC_12T_MS__XOR2_L%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%A N_A_c_189_n N_A_M1005_g N_A_c_207_n
+ N_A_M1001_g N_A_c_190_n N_A_M1010_g N_A_M1008_g N_A_c_194_n N_A_c_195_n
+ N_A_c_196_n N_A_c_200_n N_A_c_201_n N_A_c_202_n N_A_c_214_n N_A_c_203_n
+ N_A_c_218_n N_A_c_204_n N_A_c_205_n N_A_c_221_n N_A_c_206_n N_A_c_247_n
+ N_A_c_249_n A N_A_c_250_n PM_SKY130_OSU_SC_12T_MS__XOR2_L%A
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%A_238_89# N_A_238_89#_M1006_d
+ N_A_238_89#_M1002_d N_A_238_89#_M1011_g N_A_238_89#_M1007_g
+ N_A_238_89#_c_312_n N_A_238_89#_c_313_n N_A_238_89#_c_316_n
+ N_A_238_89#_c_318_n N_A_238_89#_c_320_n N_A_238_89#_c_321_n
+ PM_SKY130_OSU_SC_12T_MS__XOR2_L%A_238_89#
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%B N_B_c_375_n N_B_M1009_g N_B_c_390_n
+ N_B_M1004_g N_B_c_379_n N_B_c_381_n N_B_c_382_n N_B_M1006_g N_B_c_385_n
+ N_B_c_394_n N_B_M1002_g N_B_c_386_n N_B_c_387_n N_B_c_388_n B
+ PM_SKY130_OSU_SC_12T_MS__XOR2_L%B
x_PM_SKY130_OSU_SC_12T_MS__XOR2_L%Y N_Y_M1011_d N_Y_M1007_d N_Y_c_433_n
+ N_Y_c_443_n N_Y_c_450_n N_Y_c_434_n Y N_Y_c_438_n N_Y_c_439_n
+ PM_SKY130_OSU_SC_12T_MS__XOR2_L%Y
cc_1 N_GND_M1005_b N_A_27_115#_M1000_g 0.0358816f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.835
cc_2 N_GND_c_2_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.905
+ $Y2=0.835
cc_3 N_GND_c_3_p N_A_27_115#_M1000_g 0.00606474f $X=2.355 $Y=0.152 $X2=0.905
+ $Y2=0.835
cc_4 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.905
+ $Y2=0.835
cc_5 N_GND_M1005_b N_A_27_115#_c_117_n 0.0277843f $X=-0.045 $Y=0 $X2=0.845
+ $Y2=1.745
cc_6 N_GND_c_2_p N_A_27_115#_c_117_n 0.00172615f $X=0.69 $Y=0.755 $X2=0.845
+ $Y2=1.745
cc_7 N_GND_M1005_b N_A_27_115#_c_119_n 0.0287684f $X=-0.045 $Y=0 $X2=1.805
+ $Y2=2.285
cc_8 N_GND_M1005_b N_A_27_115#_c_120_n 0.028416f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_9 N_GND_c_9_p N_A_27_115#_c_120_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_10 N_GND_c_4_p N_A_27_115#_c_120_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_11 N_GND_M1005_b N_A_27_115#_c_123_n 0.0279827f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.955
cc_12 N_GND_M1005_b N_A_27_115#_c_124_n 0.0351362f $X=-0.045 $Y=0 $X2=1.72
+ $Y2=1.745
cc_13 N_GND_M1005_b N_A_27_115#_c_125_n 0.00402941f $X=-0.045 $Y=0 $X2=1.805
+ $Y2=2.285
cc_14 N_GND_M1005_b N_A_27_115#_c_126_n 0.00692367f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.745
cc_15 N_GND_M1005_b N_A_c_189_n 0.0619806f $X=-0.045 $Y=0 $X2=0.425 $Y2=2.38
cc_16 N_GND_M1005_b N_A_c_190_n 0.00178356f $X=-0.045 $Y=0 $X2=0.71 $Y2=2.455
cc_17 N_GND_M1005_b N_A_M1008_g 0.0361289f $X=-0.045 $Y=0 $X2=1.865 $Y2=0.835
cc_18 N_GND_c_3_p N_A_M1008_g 0.00606474f $X=2.355 $Y=0.152 $X2=1.865 $Y2=0.835
cc_19 N_GND_c_4_p N_A_M1008_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.865 $Y2=0.835
cc_20 N_GND_M1005_b N_A_c_194_n 0.0125853f $X=-0.045 $Y=0 $X2=2.1 $Y2=1.605
cc_21 N_GND_M1005_b N_A_c_195_n 0.00928792f $X=-0.045 $Y=0 $X2=1.94 $Y2=1.605
cc_22 N_GND_M1005_b N_A_c_196_n 0.0186719f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.17
cc_23 N_GND_c_9_p N_A_c_196_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.45 $Y2=1.17
cc_24 N_GND_c_2_p N_A_c_196_n 0.00308284f $X=0.69 $Y=0.755 $X2=0.45 $Y2=1.17
cc_25 N_GND_c_4_p N_A_c_196_n 0.00468827f $X=2.38 $Y=0.19 $X2=0.45 $Y2=1.17
cc_26 N_GND_M1005_b N_A_c_200_n 0.012055f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.295
cc_27 N_GND_M1005_b N_A_c_201_n 0.00205699f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.455
cc_28 N_GND_M1005_b N_A_c_202_n 0.0203167f $X=-0.045 $Y=0 $X2=0.845 $Y2=2.285
cc_29 N_GND_M1005_b N_A_c_203_n 0.0338763f $X=-0.045 $Y=0 $X2=2.235 $Y2=1.605
cc_30 N_GND_M1005_b N_A_c_204_n 0.00930883f $X=-0.045 $Y=0 $X2=2.145 $Y2=2.85
cc_31 N_GND_M1005_b N_A_c_205_n 0.00457153f $X=-0.045 $Y=0 $X2=0.845 $Y2=2.285
cc_32 N_GND_M1005_b N_A_c_206_n 0.00312742f $X=-0.045 $Y=0 $X2=2.235 $Y2=1.74
cc_33 N_GND_M1005_b N_A_238_89#_M1007_g 0.053375f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=3.235
cc_34 N_GND_M1005_b N_A_238_89#_c_312_n 0.0270758f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=1.37
cc_35 N_GND_M1005_b N_A_238_89#_c_313_n 0.0169421f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=1.205
cc_36 N_GND_c_3_p N_A_238_89#_c_313_n 0.00606474f $X=2.355 $Y=0.152 $X2=1.325
+ $Y2=1.205
cc_37 N_GND_c_4_p N_A_238_89#_c_313_n 0.00468827f $X=2.38 $Y=0.19 $X2=1.325
+ $Y2=1.205
cc_38 N_GND_M1005_b N_A_238_89#_c_316_n 0.026678f $X=-0.045 $Y=0 $X2=2.785
+ $Y2=1.37
cc_39 N_GND_c_39_p N_A_238_89#_c_316_n 0.00756829f $X=2.44 $Y=0.755 $X2=2.785
+ $Y2=1.37
cc_40 N_GND_M1005_b N_A_238_89#_c_318_n 0.0176967f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=0.755
cc_41 N_GND_c_4_p N_A_238_89#_c_318_n 0.00476261f $X=2.38 $Y=0.19 $X2=2.87
+ $Y2=0.755
cc_42 N_GND_M1005_b N_A_238_89#_c_320_n 0.045758f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=2.955
cc_43 N_GND_M1005_b N_A_238_89#_c_321_n 0.00720662f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=1.37
cc_44 N_GND_M1005_b N_B_c_375_n 0.0139689f $X=-0.045 $Y=0 $X2=2.225 $Y2=1.17
cc_45 N_GND_c_3_p N_B_c_375_n 0.00606474f $X=2.355 $Y=0.152 $X2=2.225 $Y2=1.17
cc_46 N_GND_c_39_p N_B_c_375_n 0.00308284f $X=2.44 $Y=0.755 $X2=2.225 $Y2=1.17
cc_47 N_GND_c_4_p N_B_c_375_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.225 $Y2=1.17
cc_48 N_GND_M1005_b N_B_c_379_n 0.0134223f $X=-0.045 $Y=0 $X2=2.58 $Y2=1.245
cc_49 N_GND_c_39_p N_B_c_379_n 0.00209358f $X=2.44 $Y=0.755 $X2=2.58 $Y2=1.245
cc_50 N_GND_M1005_b N_B_c_381_n 0.00622799f $X=-0.045 $Y=0 $X2=2.3 $Y2=1.245
cc_51 N_GND_M1005_b N_B_c_382_n 0.0243938f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.17
cc_52 N_GND_c_39_p N_B_c_382_n 0.00308284f $X=2.44 $Y=0.755 $X2=2.655 $Y2=1.17
cc_53 N_GND_c_4_p N_B_c_382_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.655 $Y2=1.17
cc_54 N_GND_M1005_b N_B_c_385_n 0.0434452f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.12
cc_55 N_GND_M1005_b N_B_c_386_n 0.0377483f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.325
cc_56 N_GND_M1005_b N_B_c_387_n 0.0061678f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.245
cc_57 N_GND_M1005_b N_B_c_388_n 0.00229251f $X=-0.045 $Y=0 $X2=2.53 $Y2=2.285
cc_58 N_GND_M1005_b B 2.21435e-19 $X=-0.045 $Y=0 $X2=2.53 $Y2=2.48
cc_59 N_GND_M1005_b N_Y_c_433_n 0.00910143f $X=-0.045 $Y=0 $X2=1.425 $Y2=2.11
cc_60 N_GND_M1005_b N_Y_c_434_n 0.00311329f $X=-0.045 $Y=0 $X2=1.565 $Y2=0.755
cc_61 N_GND_c_3_p N_Y_c_434_n 0.0144921f $X=2.355 $Y=0.152 $X2=1.565 $Y2=0.755
cc_62 N_GND_c_4_p N_Y_c_434_n 0.00949033f $X=2.38 $Y=0.19 $X2=1.565 $Y2=0.755
cc_63 N_GND_M1005_b Y 0.00678007f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.95
cc_64 N_GND_M1005_b N_Y_c_438_n 0.00252706f $X=-0.045 $Y=0 $X2=1.425 $Y2=2.11
cc_65 N_GND_M1005_b N_Y_c_439_n 0.00176349f $X=-0.045 $Y=0 $X2=1.425 $Y2=1
cc_66 N_GND_c_2_p N_Y_c_439_n 3.91112e-19 $X=0.69 $Y=0.755 $X2=1.425 $Y2=1
cc_67 N_GND_c_3_p N_Y_c_439_n 0.00186144f $X=2.355 $Y=0.152 $X2=1.425 $Y2=1
cc_68 N_VDD_M1001_b N_A_27_115#_M1003_g 0.020026f $X=-0.045 $Y=2.425 $X2=1.865
+ $Y2=3.235
cc_69 N_VDD_c_69_p N_A_27_115#_M1003_g 0.00606474f $X=2.355 $Y=4.287 $X2=1.865
+ $Y2=3.235
cc_70 N_VDD_c_70_p N_A_27_115#_M1003_g 0.00468827f $X=2.38 $Y=4.25 $X2=1.865
+ $Y2=3.235
cc_71 N_VDD_M1001_b N_A_27_115#_c_119_n 0.00494544f $X=-0.045 $Y=2.425 $X2=1.805
+ $Y2=2.285
cc_72 N_VDD_M1001_b N_A_27_115#_c_123_n 0.0102731f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=2.955
cc_73 N_VDD_c_73_p N_A_27_115#_c_123_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=2.955
cc_74 N_VDD_c_70_p N_A_27_115#_c_123_n 0.00476261f $X=2.38 $Y=4.25 $X2=0.26
+ $Y2=2.955
cc_75 N_VDD_M1001_b N_A_27_115#_c_125_n 9.80914e-19 $X=-0.045 $Y=2.425 $X2=1.805
+ $Y2=2.285
cc_76 N_VDD_M1001_b N_A_c_207_n 0.0183137f $X=-0.045 $Y=2.425 $X2=0.475 $Y2=2.53
cc_77 N_VDD_c_73_p N_A_c_207_n 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=2.53
cc_78 N_VDD_c_78_p N_A_c_207_n 0.00337744f $X=0.69 $Y=3.635 $X2=0.475 $Y2=2.53
cc_79 N_VDD_c_70_p N_A_c_207_n 0.00468827f $X=2.38 $Y=4.25 $X2=0.475 $Y2=2.53
cc_80 N_VDD_M1001_b N_A_c_190_n 0.00557443f $X=-0.045 $Y=2.425 $X2=0.71
+ $Y2=2.455
cc_81 N_VDD_M1001_b N_A_c_201_n 0.00756323f $X=-0.045 $Y=2.425 $X2=0.45
+ $Y2=2.455
cc_82 N_VDD_M1001_b N_A_c_202_n 0.00635728f $X=-0.045 $Y=2.425 $X2=0.845
+ $Y2=2.285
cc_83 N_VDD_M1001_b N_A_c_214_n 0.0136345f $X=-0.045 $Y=2.425 $X2=0.845 $Y2=2.53
cc_84 N_VDD_c_78_p N_A_c_214_n 0.00337744f $X=0.69 $Y=3.635 $X2=0.845 $Y2=2.53
cc_85 N_VDD_c_69_p N_A_c_214_n 0.00606474f $X=2.355 $Y=4.287 $X2=0.845 $Y2=2.53
cc_86 N_VDD_c_70_p N_A_c_214_n 0.00468827f $X=2.38 $Y=4.25 $X2=0.845 $Y2=2.53
cc_87 N_VDD_M1001_d N_A_c_218_n 0.00200838f $X=0.55 $Y=2.605 $X2=0.845 $Y2=2.765
cc_88 N_VDD_M1001_b N_A_c_218_n 6.29066e-19 $X=-0.045 $Y=2.425 $X2=0.845
+ $Y2=2.765
cc_89 N_VDD_M1001_b N_A_c_204_n 0.00153939f $X=-0.045 $Y=2.425 $X2=2.145
+ $Y2=2.85
cc_90 N_VDD_M1001_d N_A_c_221_n 0.00237538f $X=0.55 $Y=2.605 $X2=1.085 $Y2=2.85
cc_91 N_VDD_c_78_p N_A_c_221_n 4.80344e-19 $X=0.69 $Y=3.635 $X2=1.085 $Y2=2.85
cc_92 N_VDD_M1001_b N_A_238_89#_M1007_g 0.0213207f $X=-0.045 $Y=2.425 $X2=1.265
+ $Y2=3.235
cc_93 N_VDD_c_69_p N_A_238_89#_M1007_g 0.00606474f $X=2.355 $Y=4.287 $X2=1.265
+ $Y2=3.235
cc_94 N_VDD_c_70_p N_A_238_89#_M1007_g 0.00468827f $X=2.38 $Y=4.25 $X2=1.265
+ $Y2=3.235
cc_95 N_VDD_M1001_b N_A_238_89#_c_320_n 0.00972264f $X=-0.045 $Y=2.425 $X2=2.87
+ $Y2=2.955
cc_96 N_VDD_c_96_p N_A_238_89#_c_320_n 0.00757793f $X=2.38 $Y=4.25 $X2=2.87
+ $Y2=2.955
cc_97 N_VDD_c_70_p N_A_238_89#_c_320_n 0.00476261f $X=2.38 $Y=4.25 $X2=2.87
+ $Y2=2.955
cc_98 N_VDD_M1001_b N_B_c_390_n 0.0133577f $X=-0.045 $Y=2.425 $X2=2.225 $Y2=2.53
cc_99 N_VDD_c_69_p N_B_c_390_n 0.00606474f $X=2.355 $Y=4.287 $X2=2.225 $Y2=2.53
cc_100 N_VDD_c_100_p N_B_c_390_n 0.00337744f $X=2.44 $Y=3.635 $X2=2.225 $Y2=2.53
cc_101 N_VDD_c_70_p N_B_c_390_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.225 $Y2=2.53
cc_102 N_VDD_M1001_b N_B_c_394_n 0.0180645f $X=-0.045 $Y=2.425 $X2=2.655
+ $Y2=2.53
cc_103 N_VDD_c_100_p N_B_c_394_n 0.00337744f $X=2.44 $Y=3.635 $X2=2.655 $Y2=2.53
cc_104 N_VDD_c_96_p N_B_c_394_n 0.00606474f $X=2.38 $Y=4.25 $X2=2.655 $Y2=2.53
cc_105 N_VDD_c_70_p N_B_c_394_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.655 $Y2=2.53
cc_106 N_VDD_M1001_b N_B_c_386_n 0.0132516f $X=-0.045 $Y=2.425 $X2=2.655
+ $Y2=2.325
cc_107 N_VDD_M1001_b N_B_c_388_n 0.00187626f $X=-0.045 $Y=2.425 $X2=2.53
+ $Y2=2.285
cc_108 N_VDD_M1001_b B 0.0105467f $X=-0.045 $Y=2.425 $X2=2.53 $Y2=2.48
cc_109 N_VDD_M1001_b N_Y_c_433_n 0.00419006f $X=-0.045 $Y=2.425 $X2=1.425
+ $Y2=2.11
cc_110 N_VDD_M1001_b N_Y_c_443_n 0.00313975f $X=-0.045 $Y=2.425 $X2=1.565
+ $Y2=2.955
cc_111 N_VDD_c_69_p N_Y_c_443_n 0.0149397f $X=2.355 $Y=4.287 $X2=1.565 $Y2=2.955
cc_112 N_VDD_c_70_p N_Y_c_443_n 0.00958198f $X=2.38 $Y=4.25 $X2=1.565 $Y2=2.955
cc_113 N_A_27_115#_M1000_g N_A_c_189_n 0.010446f $X=0.905 $Y=0.835 $X2=0.425
+ $Y2=2.38
cc_114 N_A_27_115#_c_117_n N_A_c_189_n 0.0212638f $X=0.845 $Y=1.745 $X2=0.425
+ $Y2=2.38
cc_115 N_A_27_115#_c_123_n N_A_c_189_n 0.0250234f $X=0.26 $Y=2.955 $X2=0.425
+ $Y2=2.38
cc_116 N_A_27_115#_c_124_n N_A_c_189_n 0.0200248f $X=1.72 $Y=1.745 $X2=0.425
+ $Y2=2.38
cc_117 N_A_27_115#_c_123_n N_A_c_207_n 0.00550627f $X=0.26 $Y=2.955 $X2=0.475
+ $Y2=2.53
cc_118 N_A_27_115#_c_124_n N_A_c_190_n 8.37626e-19 $X=1.72 $Y=1.745 $X2=0.71
+ $Y2=2.455
cc_119 N_A_27_115#_c_119_n N_A_c_195_n 0.00428847f $X=1.805 $Y=2.285 $X2=1.94
+ $Y2=1.605
cc_120 N_A_27_115#_c_124_n N_A_c_195_n 0.00407778f $X=1.72 $Y=1.745 $X2=1.94
+ $Y2=1.605
cc_121 N_A_27_115#_M1000_g N_A_c_196_n 0.0206211f $X=0.905 $Y=0.835 $X2=0.45
+ $Y2=1.17
cc_122 N_A_27_115#_c_120_n N_A_c_196_n 0.00564955f $X=0.26 $Y=0.755 $X2=0.45
+ $Y2=1.17
cc_123 N_A_27_115#_c_120_n N_A_c_200_n 0.0202283f $X=0.26 $Y=0.755 $X2=0.45
+ $Y2=1.295
cc_124 N_A_27_115#_c_124_n N_A_c_200_n 0.00168707f $X=1.72 $Y=1.745 $X2=0.45
+ $Y2=1.295
cc_125 N_A_27_115#_c_117_n N_A_c_202_n 0.0184982f $X=0.845 $Y=1.745 $X2=0.845
+ $Y2=2.285
cc_126 N_A_27_115#_c_124_n N_A_c_202_n 9.97344e-19 $X=1.72 $Y=1.745 $X2=0.845
+ $Y2=2.285
cc_127 N_A_27_115#_c_124_n N_A_c_203_n 0.0010613f $X=1.72 $Y=1.745 $X2=2.235
+ $Y2=1.605
cc_128 N_A_27_115#_c_125_n N_A_c_203_n 4.73221e-19 $X=1.805 $Y=2.285 $X2=2.235
+ $Y2=1.605
cc_129 N_A_27_115#_c_123_n N_A_c_218_n 0.0118732f $X=0.26 $Y=2.955 $X2=0.845
+ $Y2=2.765
cc_130 N_A_27_115#_c_119_n N_A_c_204_n 0.00657692f $X=1.805 $Y=2.285 $X2=2.145
+ $Y2=2.85
cc_131 N_A_27_115#_c_124_n N_A_c_204_n 4.20036e-19 $X=1.72 $Y=1.745 $X2=2.145
+ $Y2=2.85
cc_132 N_A_27_115#_c_125_n N_A_c_204_n 0.0441291f $X=1.805 $Y=2.285 $X2=2.145
+ $Y2=2.85
cc_133 N_A_27_115#_c_117_n N_A_c_205_n 9.48646e-19 $X=0.845 $Y=1.745 $X2=0.845
+ $Y2=2.285
cc_134 N_A_27_115#_c_123_n N_A_c_205_n 0.00840379f $X=0.26 $Y=2.955 $X2=0.845
+ $Y2=2.285
cc_135 N_A_27_115#_c_124_n N_A_c_205_n 0.0130076f $X=1.72 $Y=1.745 $X2=0.845
+ $Y2=2.285
cc_136 N_A_27_115#_c_124_n N_A_c_206_n 0.0140397f $X=1.72 $Y=1.745 $X2=2.235
+ $Y2=1.74
cc_137 N_A_27_115#_M1003_g N_A_c_247_n 0.0126423f $X=1.865 $Y=3.235 $X2=2
+ $Y2=2.85
cc_138 N_A_27_115#_c_125_n N_A_c_247_n 0.00625535f $X=1.805 $Y=2.285 $X2=2
+ $Y2=2.85
cc_139 N_A_27_115#_c_123_n N_A_c_249_n 0.00186628f $X=0.26 $Y=2.955 $X2=1.23
+ $Y2=2.85
cc_140 N_A_27_115#_M1003_g N_A_c_250_n 9.56269e-19 $X=1.865 $Y=3.235 $X2=2.145
+ $Y2=2.85
cc_141 N_A_27_115#_M1003_g N_A_238_89#_M1007_g 0.0306522f $X=1.865 $Y=3.235
+ $X2=1.265 $Y2=3.235
cc_142 N_A_27_115#_c_119_n N_A_238_89#_M1007_g 0.0104023f $X=1.805 $Y=2.285
+ $X2=1.265 $Y2=3.235
cc_143 N_A_27_115#_c_124_n N_A_238_89#_M1007_g 0.0147853f $X=1.72 $Y=1.745
+ $X2=1.265 $Y2=3.235
cc_144 N_A_27_115#_c_125_n N_A_238_89#_M1007_g 0.00467915f $X=1.805 $Y=2.285
+ $X2=1.265 $Y2=3.235
cc_145 N_A_27_115#_c_117_n N_A_238_89#_c_312_n 0.0459061f $X=0.845 $Y=1.745
+ $X2=1.325 $Y2=1.37
cc_146 N_A_27_115#_c_124_n N_A_238_89#_c_312_n 0.00220335f $X=1.72 $Y=1.745
+ $X2=1.325 $Y2=1.37
cc_147 N_A_27_115#_M1000_g N_A_238_89#_c_313_n 0.0459061f $X=0.905 $Y=0.835
+ $X2=1.325 $Y2=1.205
cc_148 N_A_27_115#_M1000_g N_A_238_89#_c_316_n 0.00444529f $X=0.905 $Y=0.835
+ $X2=2.785 $Y2=1.37
cc_149 N_A_27_115#_c_119_n N_A_238_89#_c_316_n 5.57661e-19 $X=1.805 $Y=2.285
+ $X2=2.785 $Y2=1.37
cc_150 N_A_27_115#_c_124_n N_A_238_89#_c_316_n 0.0449127f $X=1.72 $Y=1.745
+ $X2=2.785 $Y2=1.37
cc_151 N_A_27_115#_M1003_g N_B_c_390_n 0.0491054f $X=1.865 $Y=3.235 $X2=2.225
+ $Y2=2.53
cc_152 N_A_27_115#_c_119_n N_B_c_386_n 0.0541601f $X=1.805 $Y=2.285 $X2=2.655
+ $Y2=2.325
cc_153 N_A_27_115#_M1003_g N_Y_c_433_n 0.00249536f $X=1.865 $Y=3.235 $X2=1.425
+ $Y2=2.11
cc_154 N_A_27_115#_c_119_n N_Y_c_433_n 0.00232323f $X=1.805 $Y=2.285 $X2=1.425
+ $Y2=2.11
cc_155 N_A_27_115#_c_124_n N_Y_c_433_n 0.0106304f $X=1.72 $Y=1.745 $X2=1.425
+ $Y2=2.11
cc_156 N_A_27_115#_c_125_n N_Y_c_433_n 0.0239314f $X=1.805 $Y=2.285 $X2=1.425
+ $Y2=2.11
cc_157 N_A_27_115#_M1003_g N_Y_c_450_n 0.00742342f $X=1.865 $Y=3.235 $X2=1.537
+ $Y2=2.895
cc_158 N_A_27_115#_c_119_n N_Y_c_450_n 0.00211862f $X=1.805 $Y=2.285 $X2=1.537
+ $Y2=2.895
cc_159 N_A_27_115#_c_125_n N_Y_c_450_n 6.46587e-19 $X=1.805 $Y=2.285 $X2=1.537
+ $Y2=2.895
cc_160 N_A_27_115#_M1000_g Y 0.00162478f $X=0.905 $Y=0.835 $X2=1.425 $Y2=1.95
cc_161 N_A_27_115#_c_124_n Y 0.0149378f $X=1.72 $Y=1.745 $X2=1.425 $Y2=1.95
cc_162 N_A_27_115#_c_125_n Y 0.00729051f $X=1.805 $Y=2.285 $X2=1.425 $Y2=1.95
cc_163 N_A_27_115#_c_119_n N_Y_c_438_n 0.00177801f $X=1.805 $Y=2.285 $X2=1.425
+ $Y2=2.11
cc_164 N_A_27_115#_c_124_n N_Y_c_438_n 0.00529564f $X=1.72 $Y=1.745 $X2=1.425
+ $Y2=2.11
cc_165 N_A_27_115#_c_125_n N_Y_c_438_n 0.00741445f $X=1.805 $Y=2.285 $X2=1.425
+ $Y2=2.11
cc_166 N_A_27_115#_M1000_g N_Y_c_439_n 0.00127075f $X=0.905 $Y=0.835 $X2=1.425
+ $Y2=1
cc_167 N_A_c_189_n N_A_238_89#_M1007_g 0.00462097f $X=0.425 $Y=2.38 $X2=1.265
+ $Y2=3.235
cc_168 N_A_c_195_n N_A_238_89#_M1007_g 0.00424093f $X=1.94 $Y=1.605 $X2=1.265
+ $Y2=3.235
cc_169 N_A_c_202_n N_A_238_89#_M1007_g 0.114385f $X=0.845 $Y=2.285 $X2=1.265
+ $Y2=3.235
cc_170 N_A_c_218_n N_A_238_89#_M1007_g 0.00122231f $X=0.845 $Y=2.765 $X2=1.265
+ $Y2=3.235
cc_171 N_A_c_205_n N_A_238_89#_M1007_g 0.00120277f $X=0.845 $Y=2.285 $X2=1.265
+ $Y2=3.235
cc_172 N_A_c_221_n N_A_238_89#_M1007_g 7.7948e-19 $X=1.085 $Y=2.85 $X2=1.265
+ $Y2=3.235
cc_173 N_A_c_247_n N_A_238_89#_M1007_g 0.00913315f $X=2 $Y=2.85 $X2=1.265
+ $Y2=3.235
cc_174 N_A_c_249_n N_A_238_89#_M1007_g 0.00504822f $X=1.23 $Y=2.85 $X2=1.265
+ $Y2=3.235
cc_175 N_A_M1008_g N_A_238_89#_c_312_n 0.0126897f $X=1.865 $Y=0.835 $X2=1.325
+ $Y2=1.37
cc_176 N_A_M1008_g N_A_238_89#_c_313_n 0.0172863f $X=1.865 $Y=0.835 $X2=1.325
+ $Y2=1.205
cc_177 N_A_M1008_g N_A_238_89#_c_316_n 0.0169961f $X=1.865 $Y=0.835 $X2=2.785
+ $Y2=1.37
cc_178 N_A_c_194_n N_A_238_89#_c_316_n 0.00822635f $X=2.1 $Y=1.605 $X2=2.785
+ $Y2=1.37
cc_179 N_A_c_206_n N_A_238_89#_c_316_n 0.0216132f $X=2.235 $Y=1.74 $X2=2.785
+ $Y2=1.37
cc_180 N_A_c_204_n N_A_238_89#_c_320_n 0.0129458f $X=2.145 $Y=2.85 $X2=2.87
+ $Y2=2.955
cc_181 N_A_c_206_n N_A_238_89#_c_320_n 0.00757462f $X=2.235 $Y=1.74 $X2=2.87
+ $Y2=2.955
cc_182 N_A_c_250_n N_A_238_89#_c_320_n 0.00547471f $X=2.145 $Y=2.85 $X2=2.87
+ $Y2=2.955
cc_183 N_A_M1008_g N_B_c_375_n 0.0545838f $X=1.865 $Y=0.835 $X2=2.225 $Y2=1.17
cc_184 N_A_c_204_n N_B_c_390_n 0.0110965f $X=2.145 $Y=2.85 $X2=2.225 $Y2=2.53
cc_185 N_A_c_250_n N_B_c_390_n 0.0108195f $X=2.145 $Y=2.85 $X2=2.225 $Y2=2.53
cc_186 N_A_c_203_n N_B_c_381_n 0.0137512f $X=2.235 $Y=1.605 $X2=2.3 $Y2=1.245
cc_187 N_A_M1008_g N_B_c_385_n 0.00230834f $X=1.865 $Y=0.835 $X2=2.655 $Y2=2.12
cc_188 N_A_c_203_n N_B_c_385_n 0.0234824f $X=2.235 $Y=1.605 $X2=2.655 $Y2=2.12
cc_189 N_A_c_204_n N_B_c_385_n 0.00252389f $X=2.145 $Y=2.85 $X2=2.655 $Y2=2.12
cc_190 N_A_c_206_n N_B_c_385_n 0.00130506f $X=2.235 $Y=1.74 $X2=2.655 $Y2=2.12
cc_191 N_A_c_204_n N_B_c_394_n 0.00146094f $X=2.145 $Y=2.85 $X2=2.655 $Y2=2.53
cc_192 N_A_c_250_n N_B_c_394_n 0.00122438f $X=2.145 $Y=2.85 $X2=2.655 $Y2=2.53
cc_193 N_A_c_203_n N_B_c_386_n 0.0057573f $X=2.235 $Y=1.605 $X2=2.655 $Y2=2.325
cc_194 N_A_c_204_n N_B_c_386_n 0.00757946f $X=2.145 $Y=2.85 $X2=2.655 $Y2=2.325
cc_195 N_A_c_206_n N_B_c_386_n 0.0016552f $X=2.235 $Y=1.74 $X2=2.655 $Y2=2.325
cc_196 N_A_c_204_n N_B_c_388_n 0.0237616f $X=2.145 $Y=2.85 $X2=2.53 $Y2=2.285
cc_197 N_A_c_203_n B 5.32411e-19 $X=2.235 $Y=1.605 $X2=2.53 $Y2=2.48
cc_198 N_A_c_204_n B 0.00707785f $X=2.145 $Y=2.85 $X2=2.53 $Y2=2.48
cc_199 N_A_c_206_n B 0.00327406f $X=2.235 $Y=1.74 $X2=2.53 $Y2=2.48
cc_200 N_A_c_250_n B 0.00136805f $X=2.145 $Y=2.85 $X2=2.53 $Y2=2.48
cc_201 N_A_c_221_n A_196_521# 0.00327132f $X=1.085 $Y=2.85 $X2=0.98 $Y2=2.605
cc_202 N_A_c_249_n A_196_521# 0.0158919f $X=1.23 $Y=2.85 $X2=0.98 $Y2=2.605
cc_203 N_A_c_247_n N_Y_M1007_d 0.00470028f $X=2 $Y=2.85 $X2=1.34 $Y2=2.605
cc_204 N_A_c_218_n N_Y_c_433_n 0.0110423f $X=0.845 $Y=2.765 $X2=1.425 $Y2=2.11
cc_205 N_A_c_204_n N_Y_c_433_n 0.00873529f $X=2.145 $Y=2.85 $X2=1.425 $Y2=2.11
cc_206 N_A_c_205_n N_Y_c_433_n 0.00811087f $X=0.845 $Y=2.285 $X2=1.425 $Y2=2.11
cc_207 N_A_c_221_n N_Y_c_443_n 0.00106197f $X=1.085 $Y=2.85 $X2=1.565 $Y2=2.955
cc_208 N_A_c_247_n N_Y_c_443_n 0.020967f $X=2 $Y=2.85 $X2=1.565 $Y2=2.955
cc_209 N_A_c_249_n N_Y_c_443_n 0.00145646f $X=1.23 $Y=2.85 $X2=1.565 $Y2=2.955
cc_210 N_A_c_250_n N_Y_c_443_n 0.00142425f $X=2.145 $Y=2.85 $X2=1.565 $Y2=2.955
cc_211 N_A_c_204_n N_Y_c_450_n 0.00530707f $X=2.145 $Y=2.85 $X2=1.537 $Y2=2.895
cc_212 N_A_c_221_n N_Y_c_450_n 0.00470321f $X=1.085 $Y=2.85 $X2=1.537 $Y2=2.895
cc_213 N_A_c_247_n N_Y_c_450_n 0.0217901f $X=2 $Y=2.85 $X2=1.537 $Y2=2.895
cc_214 N_A_c_249_n N_Y_c_450_n 9.55407e-19 $X=1.23 $Y=2.85 $X2=1.537 $Y2=2.895
cc_215 N_A_c_250_n N_Y_c_450_n 8.57579e-19 $X=2.145 $Y=2.85 $X2=1.537 $Y2=2.895
cc_216 N_A_M1008_g N_Y_c_434_n 0.00296624f $X=1.865 $Y=0.835 $X2=1.565 $Y2=0.755
cc_217 N_A_M1008_g Y 0.00504329f $X=1.865 $Y=0.835 $X2=1.425 $Y2=1.95
cc_218 N_A_c_204_n Y 2.67392e-19 $X=2.145 $Y=2.85 $X2=1.425 $Y2=1.95
cc_219 N_A_c_206_n Y 7.53753e-19 $X=2.235 $Y=1.74 $X2=1.425 $Y2=1.95
cc_220 N_A_c_202_n N_Y_c_438_n 3.98944e-19 $X=0.845 $Y=2.285 $X2=1.425 $Y2=2.11
cc_221 N_A_c_205_n N_Y_c_438_n 6.11977e-19 $X=0.845 $Y=2.285 $X2=1.425 $Y2=2.11
cc_222 N_A_c_247_n N_Y_c_438_n 0.0126696f $X=2 $Y=2.85 $X2=1.425 $Y2=2.11
cc_223 N_A_M1008_g N_Y_c_439_n 0.00334017f $X=1.865 $Y=0.835 $X2=1.425 $Y2=1
cc_224 N_A_c_204_n A_388_521# 0.003952f $X=2.145 $Y=2.85 $X2=1.94 $Y2=2.605
cc_225 N_A_c_247_n A_388_521# 0.00457146f $X=2 $Y=2.85 $X2=1.94 $Y2=2.605
cc_226 N_A_c_250_n A_388_521# 0.00897914f $X=2.145 $Y=2.85 $X2=1.94 $Y2=2.605
cc_227 N_A_238_89#_c_316_n N_B_c_379_n 0.0123371f $X=2.785 $Y=1.37 $X2=2.58
+ $Y2=1.245
cc_228 N_A_238_89#_c_316_n N_B_c_381_n 0.00821444f $X=2.785 $Y=1.37 $X2=2.3
+ $Y2=1.245
cc_229 N_A_238_89#_c_318_n N_B_c_382_n 0.0108893f $X=2.87 $Y=0.755 $X2=2.655
+ $Y2=1.17
cc_230 N_A_238_89#_c_316_n N_B_c_385_n 0.0113699f $X=2.785 $Y=1.37 $X2=2.655
+ $Y2=2.12
cc_231 N_A_238_89#_c_320_n N_B_c_385_n 0.0371046f $X=2.87 $Y=2.955 $X2=2.655
+ $Y2=2.12
cc_232 N_A_238_89#_c_316_n N_B_c_386_n 0.00171569f $X=2.785 $Y=1.37 $X2=2.655
+ $Y2=2.325
cc_233 N_A_238_89#_c_316_n N_B_c_387_n 0.00775577f $X=2.785 $Y=1.37 $X2=2.655
+ $Y2=1.245
cc_234 N_A_238_89#_c_316_n N_B_c_388_n 0.00443258f $X=2.785 $Y=1.37 $X2=2.53
+ $Y2=2.285
cc_235 N_A_238_89#_c_320_n N_B_c_388_n 0.0299635f $X=2.87 $Y=2.955 $X2=2.53
+ $Y2=2.285
cc_236 N_A_238_89#_c_320_n B 0.00657877f $X=2.87 $Y=2.955 $X2=2.53 $Y2=2.48
cc_237 N_A_238_89#_M1007_g N_Y_c_433_n 0.0124336f $X=1.265 $Y=3.235 $X2=1.425
+ $Y2=2.11
cc_238 N_A_238_89#_M1007_g N_Y_c_443_n 0.00614636f $X=1.265 $Y=3.235 $X2=1.565
+ $Y2=2.955
cc_239 N_A_238_89#_c_312_n N_Y_c_434_n 9.91436e-19 $X=1.325 $Y=1.37 $X2=1.565
+ $Y2=0.755
cc_240 N_A_238_89#_c_313_n N_Y_c_434_n 0.00514837f $X=1.325 $Y=1.205 $X2=1.565
+ $Y2=0.755
cc_241 N_A_238_89#_c_316_n N_Y_c_434_n 0.0150435f $X=2.785 $Y=1.37 $X2=1.565
+ $Y2=0.755
cc_242 N_A_238_89#_M1007_g Y 0.00604691f $X=1.265 $Y=3.235 $X2=1.425 $Y2=1.95
cc_243 N_A_238_89#_c_312_n Y 0.00612713f $X=1.325 $Y=1.37 $X2=1.425 $Y2=1.95
cc_244 N_A_238_89#_c_316_n Y 0.0165787f $X=2.785 $Y=1.37 $X2=1.425 $Y2=1.95
cc_245 N_A_238_89#_M1007_g N_Y_c_438_n 0.00966885f $X=1.265 $Y=3.235 $X2=1.425
+ $Y2=2.11
cc_246 N_A_238_89#_c_313_n N_Y_c_439_n 0.0053972f $X=1.325 $Y=1.205 $X2=1.425
+ $Y2=1
cc_247 N_A_238_89#_c_316_n N_Y_c_439_n 0.00572048f $X=2.785 $Y=1.37 $X2=1.425
+ $Y2=1
