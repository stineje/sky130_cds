* File: sky130_osu_sc_18T_ls__dffr_l.pxi.spice
* Created: Thu Oct 29 17:35:38 2020
* 
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%GND N_GND_M1017_s N_GND_M1014_s N_GND_M1001_d
+ N_GND_M1003_s N_GND_M1022_d N_GND_M1018_d N_GND_M1007_s N_GND_M1008_d
+ N_GND_M1012_d N_GND_M1017_b N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_12_p
+ N_GND_c_34_p N_GND_c_35_p N_GND_c_63_p N_GND_c_36_p N_GND_c_103_p N_GND_c_37_p
+ N_GND_c_79_p N_GND_c_38_p N_GND_c_17_p N_GND_c_18_p N_GND_c_166_p
+ N_GND_c_167_p GND N_GND_c_5_p PM_SKY130_OSU_SC_18T_LS__DFFR_L%GND
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%VDD N_VDD_M1013_s N_VDD_M1000_d N_VDD_M1021_s
+ N_VDD_M1028_d N_VDD_M1009_d N_VDD_M1026_d N_VDD_M1025_d N_VDD_M1013_b
+ N_VDD_c_223_p N_VDD_c_224_p N_VDD_c_243_p N_VDD_c_244_p N_VDD_c_252_p
+ N_VDD_c_279_p N_VDD_c_264_p N_VDD_c_268_p N_VDD_c_235_p N_VDD_c_236_p
+ N_VDD_c_308_p N_VDD_c_309_p VDD N_VDD_c_225_p N_VDD_c_328_p
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%VDD
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%RN N_RN_M1017_g N_RN_c_345_n N_RN_M1013_g
+ N_RN_c_347_n N_RN_c_348_n RN PM_SKY130_OSU_SC_18T_LS__DFFR_L%RN
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_110_115# N_A_110_115#_M1017_d
+ N_A_110_115#_M1013_d N_A_110_115#_c_378_n N_A_110_115#_M1014_g
+ N_A_110_115#_M1029_g N_A_110_115#_M1026_g N_A_110_115#_c_384_n
+ N_A_110_115#_M1008_g N_A_110_115#_c_388_n N_A_110_115#_c_392_n
+ N_A_110_115#_c_393_n N_A_110_115#_c_394_n N_A_110_115#_c_396_n
+ N_A_110_115#_c_397_n N_A_110_115#_c_398_n N_A_110_115#_c_407_n
+ N_A_110_115#_c_409_n N_A_110_115#_c_411_n N_A_110_115#_c_413_n
+ N_A_110_115#_c_415_n N_A_110_115#_c_417_n
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_110_115#
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_342_518# N_A_342_518#_M1027_d
+ N_A_342_518#_M1023_d N_A_342_518#_M1000_g N_A_342_518#_M1001_g
+ N_A_342_518#_c_556_n N_A_342_518#_c_572_n N_A_342_518#_c_557_n
+ N_A_342_518#_c_559_n N_A_342_518#_c_573_n N_A_342_518#_c_576_n
+ N_A_342_518#_c_561_n N_A_342_518#_c_562_n N_A_342_518#_c_577_n
+ N_A_342_518#_c_565_n N_A_342_518#_c_566_n N_A_342_518#_c_590_n
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_342_518#
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%D N_D_M1003_g N_D_M1021_g D N_D_c_643_n
+ N_D_c_644_n PM_SKY130_OSU_SC_18T_LS__DFFR_L%D
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%CK N_CK_M1023_g N_CK_M1020_g N_CK_M1015_g
+ N_CK_M1011_g N_CK_M1005_g N_CK_c_678_n N_CK_M1031_g N_CK_c_679_n N_CK_c_680_n
+ N_CK_c_685_n N_CK_c_686_n N_CK_c_687_n N_CK_c_688_n N_CK_c_689_n N_CK_c_690_n
+ N_CK_c_691_n N_CK_c_692_n N_CK_c_693_n N_CK_c_694_n N_CK_c_695_n N_CK_c_696_n
+ N_CK_c_697_n N_CK_c_698_n CK N_CK_c_700_n N_CK_c_701_n N_CK_c_702_n
+ N_CK_c_705_n N_CK_c_708_n PM_SKY130_OSU_SC_18T_LS__DFFR_L%CK
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_217_817# N_A_217_817#_M1014_d
+ N_A_217_817#_M1029_s N_A_217_817#_M1022_g N_A_217_817#_M1028_g
+ N_A_217_817#_M1019_g N_A_217_817#_M1006_g N_A_217_817#_c_905_n
+ N_A_217_817#_c_906_n N_A_217_817#_c_907_n N_A_217_817#_c_909_n
+ N_A_217_817#_c_910_n N_A_217_817#_c_911_n N_A_217_817#_c_912_n
+ N_A_217_817#_c_913_n N_A_217_817#_c_914_n N_A_217_817#_c_915_n
+ N_A_217_817#_c_960_n N_A_217_817#_c_916_n N_A_217_817#_c_918_n
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_217_817#
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_618_89# N_A_618_89#_M1005_d
+ N_A_618_89#_M1031_d N_A_618_89#_c_1037_n N_A_618_89#_M1027_g
+ N_A_618_89#_c_1040_n N_A_618_89#_c_1041_n N_A_618_89#_c_1042_n
+ N_A_618_89#_M1030_g N_A_618_89#_c_1044_n N_A_618_89#_M1010_g
+ N_A_618_89#_c_1046_n N_A_618_89#_c_1047_n N_A_618_89#_M1016_g
+ N_A_618_89#_c_1048_n N_A_618_89#_c_1049_n N_A_618_89#_c_1050_n
+ N_A_618_89#_c_1051_n N_A_618_89#_c_1053_n N_A_618_89#_c_1054_n
+ N_A_618_89#_c_1059_n N_A_618_89#_c_1072_n N_A_618_89#_c_1060_n
+ N_A_618_89#_c_1061_n N_A_618_89#_c_1062_n N_A_618_89#_c_1076_n
+ N_A_618_89#_c_1063_n PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_618_89#
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_1160_89# N_A_1160_89#_M1007_d
+ N_A_1160_89#_M1024_s N_A_1160_89#_M1018_g N_A_1160_89#_M1009_g
+ N_A_1160_89#_M1012_g N_A_1160_89#_M1025_g N_A_1160_89#_c_1234_n
+ N_A_1160_89#_c_1235_n N_A_1160_89#_c_1236_n N_A_1160_89#_c_1260_n
+ N_A_1160_89#_c_1263_n N_A_1160_89#_c_1264_n N_A_1160_89#_c_1237_n
+ N_A_1160_89#_c_1240_n N_A_1160_89#_c_1241_n N_A_1160_89#_c_1242_n
+ N_A_1160_89#_c_1243_n N_A_1160_89#_c_1244_n N_A_1160_89#_c_1245_n
+ N_A_1160_89#_c_1246_n N_A_1160_89#_c_1247_n N_A_1160_89#_c_1248_n
+ N_A_1160_89#_c_1249_n PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_1160_89#
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_998_115# N_A_998_115#_M1015_d
+ N_A_998_115#_M1010_d N_A_998_115#_M1007_g N_A_998_115#_c_1390_n
+ N_A_998_115#_M1024_g N_A_998_115#_c_1416_n N_A_998_115#_c_1417_n
+ N_A_998_115#_c_1429_n N_A_998_115#_c_1454_n N_A_998_115#_c_1393_n
+ N_A_998_115#_c_1406_n N_A_998_115#_c_1396_n N_A_998_115#_c_1398_n
+ N_A_998_115#_c_1399_n N_A_998_115#_c_1400_n N_A_998_115#_c_1401_n
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%A_998_115#
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%QN N_QN_M1012_s N_QN_M1025_s N_QN_M1004_g
+ N_QN_M1002_g N_QN_c_1521_n N_QN_c_1525_n N_QN_c_1526_n N_QN_c_1527_n
+ N_QN_c_1528_n N_QN_c_1529_n N_QN_c_1530_n N_QN_c_1531_n QN
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%QN
x_PM_SKY130_OSU_SC_18T_LS__DFFR_L%Q N_Q_M1004_d N_Q_M1002_d N_Q_c_1603_n
+ N_Q_c_1607_n N_Q_c_1605_n N_Q_c_1606_n Q N_Q_c_1612_n
+ PM_SKY130_OSU_SC_18T_LS__DFFR_L%Q
cc_1 N_GND_M1017_b N_RN_M1017_g 0.0613491f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_RN_M1017_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_RN_M1017_g 0.00606474f $X=1.125 $Y=0.152 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_RN_M1017_g 0.00394336f $X=1.21 $Y=0.825 $X2=0.475 $Y2=1.075
cc_5 N_GND_c_5_p N_RN_M1017_g 0.00468827f $X=9.175 $Y=0.17 $X2=0.475 $Y2=1.075
cc_6 N_GND_M1017_b N_RN_c_345_n 0.0376519f $X=-0.05 $Y=0 $X2=0.475 $Y2=2.47
cc_7 N_GND_M1017_b N_RN_M1013_g 0.0288885f $X=-0.05 $Y=0 $X2=0.475 $Y2=4.585
cc_8 N_GND_M1017_b N_RN_c_347_n 0.020318f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.305
cc_9 N_GND_M1017_b N_RN_c_348_n 0.0149094f $X=-0.05 $Y=0 $X2=0.32 $Y2=3.33
cc_10 N_GND_M1017_b N_A_110_115#_c_378_n 0.0183053f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=1.425
cc_11 N_GND_c_4_p N_A_110_115#_c_378_n 0.00713292f $X=1.21 $Y=0.825 $X2=1.425
+ $Y2=1.425
cc_12 N_GND_c_12_p N_A_110_115#_c_378_n 0.00606474f $X=1.985 $Y=0.152 $X2=1.425
+ $Y2=1.425
cc_13 N_GND_c_5_p N_A_110_115#_c_378_n 0.00468827f $X=9.175 $Y=0.17 $X2=1.425
+ $Y2=1.425
cc_14 N_GND_M1017_b N_A_110_115#_M1029_g 0.0665091f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=5.085
cc_15 N_GND_M1017_b N_A_110_115#_M1026_g 0.0711177f $X=-0.05 $Y=0 $X2=7.615
+ $Y2=5.085
cc_16 N_GND_M1017_b N_A_110_115#_c_384_n 0.018156f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.425
cc_17 N_GND_c_17_p N_A_110_115#_c_384_n 0.00606474f $X=7.815 $Y=0.152 $X2=7.685
+ $Y2=1.425
cc_18 N_GND_c_18_p N_A_110_115#_c_384_n 0.00713292f $X=7.9 $Y=0.825 $X2=7.685
+ $Y2=1.425
cc_19 N_GND_c_5_p N_A_110_115#_c_384_n 0.00468827f $X=9.175 $Y=0.17 $X2=7.685
+ $Y2=1.425
cc_20 N_GND_M1017_b N_A_110_115#_c_388_n 0.00156053f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=0.825
cc_21 N_GND_c_3_p N_A_110_115#_c_388_n 0.00757793f $X=1.125 $Y=0.152 $X2=0.69
+ $Y2=0.825
cc_22 N_GND_c_4_p N_A_110_115#_c_388_n 0.0213592f $X=1.21 $Y=0.825 $X2=0.69
+ $Y2=0.825
cc_23 N_GND_c_5_p N_A_110_115#_c_388_n 0.00476261f $X=9.175 $Y=0.17 $X2=0.69
+ $Y2=0.825
cc_24 N_GND_M1017_b N_A_110_115#_c_392_n 0.0021895f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=3.455
cc_25 N_GND_M1017_b N_A_110_115#_c_393_n 0.0216652f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.655
cc_26 N_GND_M1017_b N_A_110_115#_c_394_n 0.0093348f $X=-0.05 $Y=0 $X2=1.145
+ $Y2=1.59
cc_27 N_GND_c_4_p N_A_110_115#_c_394_n 4.24107e-19 $X=1.21 $Y=0.825 $X2=1.145
+ $Y2=1.59
cc_28 N_GND_M1017_b N_A_110_115#_c_396_n 0.0125851f $X=-0.05 $Y=0 $X2=0.955
+ $Y2=1.59
cc_29 N_GND_M1017_b N_A_110_115#_c_397_n 0.0162344f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.74
cc_30 N_GND_M1003_s N_A_110_115#_c_398_n 0.00506021f $X=2.465 $Y=0.575 $X2=7.665
+ $Y2=1.48
cc_31 N_GND_M1022_d N_A_110_115#_c_398_n 0.0109039f $X=4.2 $Y=0.575 $X2=7.665
+ $Y2=1.48
cc_32 N_GND_M1018_d N_A_110_115#_c_398_n 0.00557645f $X=5.95 $Y=0.575 $X2=7.665
+ $Y2=1.48
cc_33 N_GND_M1017_b N_A_110_115#_c_398_n 0.0468573f $X=-0.05 $Y=0 $X2=7.665
+ $Y2=1.48
cc_34 N_GND_c_34_p N_A_110_115#_c_398_n 0.00550371f $X=2.07 $Y=0.825 $X2=7.665
+ $Y2=1.48
cc_35 N_GND_c_35_p N_A_110_115#_c_398_n 0.0120854f $X=2.59 $Y=0.825 $X2=7.665
+ $Y2=1.48
cc_36 N_GND_c_36_p N_A_110_115#_c_398_n 0.00558854f $X=4.34 $Y=0.825 $X2=7.665
+ $Y2=1.48
cc_37 N_GND_c_37_p N_A_110_115#_c_398_n 0.0119903f $X=6.09 $Y=0.825 $X2=7.665
+ $Y2=1.48
cc_38 N_GND_c_38_p N_A_110_115#_c_398_n 0.00640729f $X=7.04 $Y=0.825 $X2=7.665
+ $Y2=1.48
cc_39 N_GND_M1017_b N_A_110_115#_c_407_n 0.00628827f $X=-0.05 $Y=0 $X2=1.375
+ $Y2=1.48
cc_40 N_GND_c_4_p N_A_110_115#_c_407_n 0.00462957f $X=1.21 $Y=0.825 $X2=1.375
+ $Y2=1.48
cc_41 N_GND_M1017_b N_A_110_115#_c_409_n 0.00303307f $X=-0.05 $Y=0 $X2=1.23
+ $Y2=1.48
cc_42 N_GND_c_4_p N_A_110_115#_c_409_n 0.00557352f $X=1.21 $Y=0.825 $X2=1.23
+ $Y2=1.48
cc_43 N_GND_M1017_b N_A_110_115#_c_411_n 0.00560955f $X=-0.05 $Y=0 $X2=7.81
+ $Y2=1.48
cc_44 N_GND_c_18_p N_A_110_115#_c_411_n 0.00509889f $X=7.9 $Y=0.825 $X2=7.81
+ $Y2=1.48
cc_45 N_GND_M1017_b N_A_110_115#_c_413_n 0.00317569f $X=-0.05 $Y=0 $X2=7.81
+ $Y2=1.48
cc_46 N_GND_c_18_p N_A_110_115#_c_413_n 0.00292873f $X=7.9 $Y=0.825 $X2=7.81
+ $Y2=1.48
cc_47 N_GND_M1017_b N_A_110_115#_c_415_n 0.042671f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=1.59
cc_48 N_GND_c_4_p N_A_110_115#_c_415_n 0.00134799f $X=1.21 $Y=0.825 $X2=1.425
+ $Y2=1.59
cc_49 N_GND_M1017_b N_A_110_115#_c_417_n 0.0413355f $X=-0.05 $Y=0 $X2=7.81
+ $Y2=1.59
cc_50 N_GND_c_18_p N_A_110_115#_c_417_n 0.00210433f $X=7.9 $Y=0.825 $X2=7.81
+ $Y2=1.59
cc_51 N_GND_M1017_b N_A_342_518#_M1001_g 0.088777f $X=-0.05 $Y=0 $X2=1.855
+ $Y2=0.945
cc_52 N_GND_c_12_p N_A_342_518#_M1001_g 0.00606474f $X=1.985 $Y=0.152 $X2=1.855
+ $Y2=0.945
cc_53 N_GND_c_34_p N_A_342_518#_M1001_g 0.00713292f $X=2.07 $Y=0.825 $X2=1.855
+ $Y2=0.945
cc_54 N_GND_c_35_p N_A_342_518#_M1001_g 0.00874269f $X=2.59 $Y=0.825 $X2=1.855
+ $Y2=0.945
cc_55 N_GND_c_5_p N_A_342_518#_M1001_g 0.00468827f $X=9.175 $Y=0.17 $X2=1.855
+ $Y2=0.945
cc_56 N_GND_M1017_b N_A_342_518#_c_556_n 0.0188271f $X=-0.05 $Y=0 $X2=2.11
+ $Y2=2.59
cc_57 N_GND_M1017_b N_A_342_518#_c_557_n 0.0219314f $X=-0.05 $Y=0 $X2=3.28
+ $Y2=1.765
cc_58 N_GND_c_35_p N_A_342_518#_c_557_n 0.00673409f $X=2.59 $Y=0.825 $X2=3.28
+ $Y2=1.765
cc_59 N_GND_M1017_b N_A_342_518#_c_559_n 0.00414603f $X=-0.05 $Y=0 $X2=2.195
+ $Y2=1.765
cc_60 N_GND_c_34_p N_A_342_518#_c_559_n 0.00187963f $X=2.07 $Y=0.825 $X2=2.195
+ $Y2=1.765
cc_61 N_GND_M1017_b N_A_342_518#_c_561_n 0.00198494f $X=-0.05 $Y=0 $X2=3.365
+ $Y2=1.68
cc_62 N_GND_M1017_b N_A_342_518#_c_562_n 0.00313975f $X=-0.05 $Y=0 $X2=3.465
+ $Y2=0.825
cc_63 N_GND_c_63_p N_A_342_518#_c_562_n 0.0151129f $X=4.255 $Y=0.152 $X2=3.465
+ $Y2=0.825
cc_64 N_GND_c_5_p N_A_342_518#_c_562_n 0.00958198f $X=9.175 $Y=0.17 $X2=3.465
+ $Y2=0.825
cc_65 N_GND_M1017_b N_A_342_518#_c_565_n 0.0338764f $X=-0.05 $Y=0 $X2=1.94
+ $Y2=2.755
cc_66 N_GND_M1017_b N_A_342_518#_c_566_n 0.00486423f $X=-0.05 $Y=0 $X2=2.11
+ $Y2=2.755
cc_67 N_GND_M1017_b N_D_M1003_g 0.0418804f $X=-0.05 $Y=0 $X2=2.805 $Y2=1.075
cc_68 N_GND_c_35_p N_D_M1003_g 0.0071489f $X=2.59 $Y=0.825 $X2=2.805 $Y2=1.075
cc_69 N_GND_c_63_p N_D_M1003_g 0.00606474f $X=4.255 $Y=0.152 $X2=2.805 $Y2=1.075
cc_70 N_GND_c_5_p N_D_M1003_g 0.00468827f $X=9.175 $Y=0.17 $X2=2.805 $Y2=1.075
cc_71 N_GND_M1017_b N_D_M1021_g 0.0360004f $X=-0.05 $Y=0 $X2=2.805 $Y2=4.585
cc_72 N_GND_M1017_b D 0.00973922f $X=-0.05 $Y=0 $X2=2.865 $Y2=2.22
cc_73 N_GND_M1017_b N_D_c_643_n 0.00311208f $X=-0.05 $Y=0 $X2=2.865 $Y2=2.22
cc_74 N_GND_M1017_b N_D_c_644_n 0.0324288f $X=-0.05 $Y=0 $X2=2.865 $Y2=2.22
cc_75 N_GND_M1017_b N_CK_c_678_n 0.0311248f $X=-0.05 $Y=0 $X2=6.305 $Y2=2.93
cc_76 N_GND_M1017_b N_CK_c_679_n 0.0442038f $X=-0.05 $Y=0 $X2=6.36 $Y2=2.6
cc_77 N_GND_M1017_b N_CK_c_680_n 0.0183851f $X=-0.05 $Y=0 $X2=6.332 $Y2=1.685
cc_78 N_GND_c_37_p N_CK_c_680_n 0.00356864f $X=6.09 $Y=0.825 $X2=6.332 $Y2=1.685
cc_79 N_GND_c_79_p N_CK_c_680_n 0.00606474f $X=6.955 $Y=0.152 $X2=6.332
+ $Y2=1.685
cc_80 N_GND_c_38_p N_CK_c_680_n 0.00394336f $X=7.04 $Y=0.825 $X2=6.332 $Y2=1.685
cc_81 N_GND_c_5_p N_CK_c_680_n 0.00468827f $X=9.175 $Y=0.17 $X2=6.332 $Y2=1.685
cc_82 N_GND_M1017_b N_CK_c_685_n 0.0131012f $X=-0.05 $Y=0 $X2=6.332 $Y2=1.835
cc_83 N_GND_M1017_b N_CK_c_686_n 0.00609317f $X=-0.05 $Y=0 $X2=3.62 $Y2=2.59
cc_84 N_GND_M1017_b N_CK_c_687_n 0.00921066f $X=-0.05 $Y=0 $X2=3.705 $Y2=1.85
cc_85 N_GND_M1017_b N_CK_c_688_n 0.0254608f $X=-0.05 $Y=0 $X2=3.705 $Y2=1.85
cc_86 N_GND_M1017_b N_CK_c_689_n 0.00838835f $X=-0.05 $Y=0 $X2=4.975 $Y2=1.85
cc_87 N_GND_M1017_b N_CK_c_690_n 0.0252285f $X=-0.05 $Y=0 $X2=4.975 $Y2=1.85
cc_88 N_GND_M1017_b N_CK_c_691_n 0.00543853f $X=-0.05 $Y=0 $X2=5.37 $Y2=2.59
cc_89 N_GND_M1017_b N_CK_c_692_n 5.00459e-19 $X=-0.05 $Y=0 $X2=5.06 $Y2=2.59
cc_90 N_GND_M1017_b N_CK_c_693_n 0.0345662f $X=-0.05 $Y=0 $X2=5.31 $Y2=2.59
cc_91 N_GND_M1017_b N_CK_c_694_n 0.00714094f $X=-0.05 $Y=0 $X2=3.37 $Y2=2.59
cc_92 N_GND_M1017_b N_CK_c_695_n 0.0181831f $X=-0.05 $Y=0 $X2=6.305 $Y2=2.59
cc_93 N_GND_M1017_b N_CK_c_696_n 0.0041728f $X=-0.05 $Y=0 $X2=5.6 $Y2=2.59
cc_94 N_GND_M1017_b N_CK_c_697_n 0.00276905f $X=-0.05 $Y=0 $X2=3.225 $Y2=2.59
cc_95 N_GND_M1017_b N_CK_c_698_n 0.00265612f $X=-0.05 $Y=0 $X2=5.455 $Y2=2.59
cc_96 N_GND_M1017_b CK 0.00239232f $X=-0.05 $Y=0 $X2=6.45 $Y2=2.59
cc_97 N_GND_M1017_b N_CK_c_700_n 7.61111e-19 $X=-0.05 $Y=0 $X2=6.45 $Y2=2.59
cc_98 N_GND_M1017_b N_CK_c_701_n 0.0244095f $X=-0.05 $Y=0 $X2=3.225 $Y2=2.765
cc_99 N_GND_M1017_b N_CK_c_702_n 0.0173906f $X=-0.05 $Y=0 $X2=3.705 $Y2=1.685
cc_100 N_GND_c_63_p N_CK_c_702_n 0.00606474f $X=4.255 $Y=0.152 $X2=3.705
+ $Y2=1.685
cc_101 N_GND_c_5_p N_CK_c_702_n 0.00468827f $X=9.175 $Y=0.17 $X2=3.705 $Y2=1.685
cc_102 N_GND_M1017_b N_CK_c_705_n 0.0175305f $X=-0.05 $Y=0 $X2=4.975 $Y2=1.685
cc_103 N_GND_c_103_p N_CK_c_705_n 0.00606474f $X=6.005 $Y=0.152 $X2=4.975
+ $Y2=1.685
cc_104 N_GND_c_5_p N_CK_c_705_n 0.00468827f $X=9.175 $Y=0.17 $X2=4.975 $Y2=1.685
cc_105 N_GND_M1017_b N_CK_c_708_n 0.0233827f $X=-0.05 $Y=0 $X2=5.455 $Y2=2.765
cc_106 N_GND_M1017_b N_A_217_817#_M1022_g 0.0171814f $X=-0.05 $Y=0 $X2=4.125
+ $Y2=1.075
cc_107 N_GND_c_63_p N_A_217_817#_M1022_g 0.00606474f $X=4.255 $Y=0.152 $X2=4.125
+ $Y2=1.075
cc_108 N_GND_c_36_p N_A_217_817#_M1022_g 0.00354579f $X=4.34 $Y=0.825 $X2=4.125
+ $Y2=1.075
cc_109 N_GND_c_5_p N_A_217_817#_M1022_g 0.00468827f $X=9.175 $Y=0.17 $X2=4.125
+ $Y2=1.075
cc_110 N_GND_M1017_b N_A_217_817#_M1019_g 0.0163216f $X=-0.05 $Y=0 $X2=4.555
+ $Y2=1.075
cc_111 N_GND_c_36_p N_A_217_817#_M1019_g 0.00354579f $X=4.34 $Y=0.825 $X2=4.555
+ $Y2=1.075
cc_112 N_GND_c_103_p N_A_217_817#_M1019_g 0.00606474f $X=6.005 $Y=0.152
+ $X2=4.555 $Y2=1.075
cc_113 N_GND_c_5_p N_A_217_817#_M1019_g 0.00468827f $X=9.175 $Y=0.17 $X2=4.555
+ $Y2=1.075
cc_114 N_GND_M1017_b N_A_217_817#_c_905_n 0.0105855f $X=-0.05 $Y=0 $X2=4.2
+ $Y2=1.85
cc_115 N_GND_M1017_b N_A_217_817#_c_906_n 0.0105265f $X=-0.05 $Y=0 $X2=4.2
+ $Y2=2.765
cc_116 N_GND_M1017_b N_A_217_817#_c_907_n 0.0240953f $X=-0.05 $Y=0 $X2=4.48
+ $Y2=1.85
cc_117 N_GND_c_36_p N_A_217_817#_c_907_n 8.07204e-19 $X=4.34 $Y=0.825 $X2=4.48
+ $Y2=1.85
cc_118 N_GND_M1017_b N_A_217_817#_c_909_n 0.0232417f $X=-0.05 $Y=0 $X2=4.48
+ $Y2=2.765
cc_119 N_GND_M1017_b N_A_217_817#_c_910_n 0.0172857f $X=-0.05 $Y=0 $X2=1.21
+ $Y2=4.475
cc_120 N_GND_M1017_b N_A_217_817#_c_911_n 0.0126209f $X=-0.05 $Y=0 $X2=1.555
+ $Y2=2.02
cc_121 N_GND_M1017_b N_A_217_817#_c_912_n 0.00251117f $X=-0.05 $Y=0 $X2=1.295
+ $Y2=2.02
cc_122 N_GND_M1017_b N_A_217_817#_c_913_n 0.00871176f $X=-0.05 $Y=0 $X2=4.295
+ $Y2=2.765
cc_123 N_GND_M1017_b N_A_217_817#_c_914_n 0.0339774f $X=-0.05 $Y=0 $X2=4.06
+ $Y2=1.85
cc_124 N_GND_M1017_b N_A_217_817#_c_915_n 0.001822f $X=-0.05 $Y=0 $X2=1.785
+ $Y2=1.85
cc_125 N_GND_M1017_b N_A_217_817#_c_916_n 0.00245573f $X=-0.05 $Y=0 $X2=4.205
+ $Y2=1.85
cc_126 N_GND_c_36_p N_A_217_817#_c_916_n 0.00177942f $X=4.34 $Y=0.825 $X2=4.205
+ $Y2=1.85
cc_127 N_GND_M1017_b N_A_217_817#_c_918_n 0.0140372f $X=-0.05 $Y=0 $X2=1.64
+ $Y2=0.825
cc_128 N_GND_c_12_p N_A_217_817#_c_918_n 0.00734006f $X=1.985 $Y=0.152 $X2=1.64
+ $Y2=0.825
cc_129 N_GND_c_5_p N_A_217_817#_c_918_n 0.00475776f $X=9.175 $Y=0.17 $X2=1.64
+ $Y2=0.825
cc_130 N_GND_M1017_b N_A_618_89#_c_1037_n 0.0173059f $X=-0.05 $Y=0 $X2=3.165
+ $Y2=1.685
cc_131 N_GND_c_63_p N_A_618_89#_c_1037_n 0.00606474f $X=4.255 $Y=0.152 $X2=3.165
+ $Y2=1.685
cc_132 N_GND_c_5_p N_A_618_89#_c_1037_n 0.00468827f $X=9.175 $Y=0.17 $X2=3.165
+ $Y2=1.685
cc_133 N_GND_M1017_b N_A_618_89#_c_1040_n 0.0203057f $X=-0.05 $Y=0 $X2=3.285
+ $Y2=2.225
cc_134 N_GND_M1017_b N_A_618_89#_c_1041_n 0.0187566f $X=-0.05 $Y=0 $X2=3.69
+ $Y2=2.3
cc_135 N_GND_M1017_b N_A_618_89#_c_1042_n 0.00755029f $X=-0.05 $Y=0 $X2=3.36
+ $Y2=2.3
cc_136 N_GND_M1017_b N_A_618_89#_M1030_g 0.032457f $X=-0.05 $Y=0 $X2=3.765
+ $Y2=4.585
cc_137 N_GND_M1017_b N_A_618_89#_c_1044_n 0.0559794f $X=-0.05 $Y=0 $X2=4.84
+ $Y2=2.3
cc_138 N_GND_M1017_b N_A_618_89#_M1010_g 0.0319667f $X=-0.05 $Y=0 $X2=4.915
+ $Y2=4.585
cc_139 N_GND_M1017_b N_A_618_89#_c_1046_n 0.0270462f $X=-0.05 $Y=0 $X2=5.32
+ $Y2=2.3
cc_140 N_GND_M1017_b N_A_618_89#_c_1047_n 0.0125754f $X=-0.05 $Y=0 $X2=5.395
+ $Y2=2.225
cc_141 N_GND_M1017_b N_A_618_89#_c_1048_n 0.0141451f $X=-0.05 $Y=0 $X2=3.285
+ $Y2=1.76
cc_142 N_GND_M1017_b N_A_618_89#_c_1049_n 0.00426512f $X=-0.05 $Y=0 $X2=3.765
+ $Y2=2.3
cc_143 N_GND_M1017_b N_A_618_89#_c_1050_n 0.00426512f $X=-0.05 $Y=0 $X2=4.915
+ $Y2=2.3
cc_144 N_GND_M1017_b N_A_618_89#_c_1051_n 0.0116005f $X=-0.05 $Y=0 $X2=6.435
+ $Y2=1.85
cc_145 N_GND_c_37_p N_A_618_89#_c_1051_n 0.00564434f $X=6.09 $Y=0.825 $X2=6.435
+ $Y2=1.85
cc_146 N_GND_M1017_b N_A_618_89#_c_1053_n 0.0256431f $X=-0.05 $Y=0 $X2=5.455
+ $Y2=1.85
cc_147 N_GND_M1017_b N_A_618_89#_c_1054_n 0.00554907f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=0.825
cc_148 N_GND_c_37_p N_A_618_89#_c_1054_n 4.65312e-19 $X=6.09 $Y=0.825 $X2=6.52
+ $Y2=0.825
cc_149 N_GND_c_79_p N_A_618_89#_c_1054_n 0.00736239f $X=6.955 $Y=0.152 $X2=6.52
+ $Y2=0.825
cc_150 N_GND_c_38_p N_A_618_89#_c_1054_n 0.0213592f $X=7.04 $Y=0.825 $X2=6.52
+ $Y2=0.825
cc_151 N_GND_c_5_p N_A_618_89#_c_1054_n 0.00476261f $X=9.175 $Y=0.17 $X2=6.52
+ $Y2=0.825
cc_152 N_GND_M1017_b N_A_618_89#_c_1059_n 0.00330742f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=2.105
cc_153 N_GND_M1017_b N_A_618_89#_c_1060_n 0.0143188f $X=-0.05 $Y=0 $X2=6.795
+ $Y2=3.1
cc_154 N_GND_M1017_b N_A_618_89#_c_1061_n 0.0012444f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=1.85
cc_155 N_GND_M1017_b N_A_618_89#_c_1062_n 0.0102335f $X=-0.05 $Y=0 $X2=6.795
+ $Y2=2.19
cc_156 N_GND_M1017_b N_A_618_89#_c_1063_n 0.01755f $X=-0.05 $Y=0 $X2=5.455
+ $Y2=1.685
cc_157 N_GND_c_103_p N_A_618_89#_c_1063_n 0.00606474f $X=6.005 $Y=0.152
+ $X2=5.455 $Y2=1.685
cc_158 N_GND_c_5_p N_A_618_89#_c_1063_n 0.00468827f $X=9.175 $Y=0.17 $X2=5.455
+ $Y2=1.685
cc_159 N_GND_M1017_b N_A_1160_89#_M1018_g 0.0319752f $X=-0.05 $Y=0 $X2=5.875
+ $Y2=1.075
cc_160 N_GND_c_103_p N_A_1160_89#_M1018_g 0.00606474f $X=6.005 $Y=0.152
+ $X2=5.875 $Y2=1.075
cc_161 N_GND_c_37_p N_A_1160_89#_M1018_g 0.00360474f $X=6.09 $Y=0.825 $X2=5.875
+ $Y2=1.075
cc_162 N_GND_c_5_p N_A_1160_89#_M1018_g 0.00468827f $X=9.175 $Y=0.17 $X2=5.875
+ $Y2=1.075
cc_163 N_GND_M1017_b N_A_1160_89#_M1009_g 0.0330331f $X=-0.05 $Y=0 $X2=5.875
+ $Y2=4.585
cc_164 N_GND_M1017_b N_A_1160_89#_M1012_g 0.0324889f $X=-0.05 $Y=0 $X2=8.635
+ $Y2=0.945
cc_165 N_GND_c_18_p N_A_1160_89#_M1012_g 0.00394336f $X=7.9 $Y=0.825 $X2=8.635
+ $Y2=0.945
cc_166 N_GND_c_166_p N_A_1160_89#_M1012_g 0.00606474f $X=8.765 $Y=0.152
+ $X2=8.635 $Y2=0.945
cc_167 N_GND_c_167_p N_A_1160_89#_M1012_g 0.00354579f $X=8.85 $Y=0.825 $X2=8.635
+ $Y2=0.945
cc_168 N_GND_c_5_p N_A_1160_89#_M1012_g 0.00468827f $X=9.175 $Y=0.17 $X2=8.635
+ $Y2=0.945
cc_169 N_GND_M1017_b N_A_1160_89#_c_1234_n 0.0140996f $X=-0.05 $Y=0 $X2=8.61
+ $Y2=1.8
cc_170 N_GND_M1017_b N_A_1160_89#_c_1235_n 0.0365245f $X=-0.05 $Y=0 $X2=8.61
+ $Y2=2.855
cc_171 N_GND_M1017_b N_A_1160_89#_c_1236_n 0.00495925f $X=-0.05 $Y=0 $X2=8.61
+ $Y2=3.005
cc_172 N_GND_M1017_b N_A_1160_89#_c_1237_n 0.0086066f $X=-0.05 $Y=0 $X2=7.47
+ $Y2=0.825
cc_173 N_GND_c_17_p N_A_1160_89#_c_1237_n 0.0075556f $X=7.815 $Y=0.152 $X2=7.47
+ $Y2=0.825
cc_174 N_GND_c_5_p N_A_1160_89#_c_1237_n 0.00475776f $X=9.175 $Y=0.17 $X2=7.47
+ $Y2=0.825
cc_175 N_GND_M1017_b N_A_1160_89#_c_1240_n 0.00534479f $X=-0.05 $Y=0 $X2=7.47
+ $Y2=3.695
cc_176 N_GND_M1017_b N_A_1160_89#_c_1241_n 0.00133335f $X=-0.05 $Y=0 $X2=7.47
+ $Y2=2.19
cc_177 N_GND_M1017_b N_A_1160_89#_c_1242_n 0.0641658f $X=-0.05 $Y=0 $X2=8.375
+ $Y2=2.19
cc_178 N_GND_M1017_b N_A_1160_89#_c_1243_n 0.00189525f $X=-0.05 $Y=0 $X2=6.08
+ $Y2=2.19
cc_179 N_GND_M1017_b N_A_1160_89#_c_1244_n 0.0039674f $X=-0.05 $Y=0 $X2=5.935
+ $Y2=2.19
cc_180 N_GND_M1017_b N_A_1160_89#_c_1245_n 0.0029877f $X=-0.05 $Y=0 $X2=8.52
+ $Y2=2.19
cc_181 N_GND_M1017_b N_A_1160_89#_c_1246_n 0.0195866f $X=-0.05 $Y=0 $X2=8.52
+ $Y2=2.19
cc_182 N_GND_M1017_b N_A_1160_89#_c_1247_n 0.0263478f $X=-0.05 $Y=0 $X2=5.935
+ $Y2=2.19
cc_183 N_GND_M1017_b N_A_1160_89#_c_1248_n 0.0296433f $X=-0.05 $Y=0 $X2=8.52
+ $Y2=2.19
cc_184 N_GND_M1017_b N_A_1160_89#_c_1249_n 0.0154776f $X=-0.05 $Y=0 $X2=8.522
+ $Y2=2.025
cc_185 N_GND_M1017_b N_A_998_115#_M1007_g 0.0337662f $X=-0.05 $Y=0 $X2=7.255
+ $Y2=0.945
cc_186 N_GND_c_38_p N_A_998_115#_M1007_g 0.00713292f $X=7.04 $Y=0.825 $X2=7.255
+ $Y2=0.945
cc_187 N_GND_c_17_p N_A_998_115#_M1007_g 0.00606474f $X=7.815 $Y=0.152 $X2=7.255
+ $Y2=0.945
cc_188 N_GND_c_5_p N_A_998_115#_M1007_g 0.00468827f $X=9.175 $Y=0.17 $X2=7.255
+ $Y2=0.945
cc_189 N_GND_M1017_b N_A_998_115#_c_1390_n 0.037144f $X=-0.05 $Y=0 $X2=7.255
+ $Y2=2.015
cc_190 N_GND_c_38_p N_A_998_115#_c_1390_n 0.00202046f $X=7.04 $Y=0.825 $X2=7.255
+ $Y2=2.015
cc_191 N_GND_M1017_b N_A_998_115#_M1024_g 0.0524105f $X=-0.05 $Y=0 $X2=7.255
+ $Y2=5.085
cc_192 N_GND_M1017_b N_A_998_115#_c_1393_n 0.00313975f $X=-0.05 $Y=0 $X2=5.215
+ $Y2=0.825
cc_193 N_GND_c_103_p N_A_998_115#_c_1393_n 0.0149205f $X=6.005 $Y=0.152
+ $X2=5.215 $Y2=0.825
cc_194 N_GND_c_5_p N_A_998_115#_c_1393_n 0.00958198f $X=9.175 $Y=0.17 $X2=5.215
+ $Y2=0.825
cc_195 N_GND_M1017_b N_A_998_115#_c_1396_n 0.0223568f $X=-0.05 $Y=0 $X2=6.985
+ $Y2=1.85
cc_196 N_GND_c_37_p N_A_998_115#_c_1396_n 5.03331e-19 $X=6.09 $Y=0.825 $X2=6.985
+ $Y2=1.85
cc_197 N_GND_M1017_b N_A_998_115#_c_1398_n 0.00120467f $X=-0.05 $Y=0 $X2=4.78
+ $Y2=1.85
cc_198 N_GND_M1017_b N_A_998_115#_c_1399_n 0.0112983f $X=-0.05 $Y=0 $X2=4.635
+ $Y2=1.85
cc_199 N_GND_M1017_b N_A_998_115#_c_1400_n 7.27503e-19 $X=-0.05 $Y=0 $X2=7.13
+ $Y2=1.85
cc_200 N_GND_M1017_b N_A_998_115#_c_1401_n 0.00230483f $X=-0.05 $Y=0 $X2=7.13
+ $Y2=1.85
cc_201 N_GND_c_38_p N_A_998_115#_c_1401_n 9.46397e-19 $X=7.04 $Y=0.825 $X2=7.13
+ $Y2=1.85
cc_202 N_GND_M1017_b N_QN_M1004_g 0.0707753f $X=-0.05 $Y=0 $X2=9.065 $Y2=0.945
cc_203 N_GND_c_167_p N_QN_M1004_g 0.00354579f $X=8.85 $Y=0.825 $X2=9.065
+ $Y2=0.945
cc_204 N_GND_c_5_p N_QN_M1004_g 0.00468827f $X=9.175 $Y=0.17 $X2=9.065 $Y2=0.945
cc_205 N_GND_M1017_b N_QN_M1002_g 0.0186095f $X=-0.05 $Y=0 $X2=9.065 $Y2=5.085
cc_206 N_GND_M1017_b N_QN_c_1521_n 0.0114763f $X=-0.05 $Y=0 $X2=8.42 $Y2=0.825
cc_207 N_GND_c_18_p N_QN_c_1521_n 0.0213592f $X=7.9 $Y=0.825 $X2=8.42 $Y2=0.825
cc_208 N_GND_c_166_p N_QN_c_1521_n 0.00736239f $X=8.765 $Y=0.152 $X2=8.42
+ $Y2=0.825
cc_209 N_GND_c_5_p N_QN_c_1521_n 0.00476261f $X=9.175 $Y=0.17 $X2=8.42 $Y2=0.825
cc_210 N_GND_M1017_b N_QN_c_1525_n 0.0171269f $X=-0.05 $Y=0 $X2=8.92 $Y2=1.85
cc_211 N_GND_M1017_b N_QN_c_1526_n 0.00387782f $X=-0.05 $Y=0 $X2=8.505 $Y2=1.85
cc_212 N_GND_M1017_b N_QN_c_1527_n 0.0176115f $X=-0.05 $Y=0 $X2=8.92 $Y2=2.765
cc_213 N_GND_M1017_b N_QN_c_1528_n 0.00442737f $X=-0.05 $Y=0 $X2=8.505 $Y2=2.765
cc_214 N_GND_M1017_b N_QN_c_1529_n 0.0034889f $X=-0.05 $Y=0 $X2=9.005 $Y2=2.395
cc_215 N_GND_M1017_b N_QN_c_1530_n 0.0291912f $X=-0.05 $Y=0 $X2=9.005 $Y2=2.395
cc_216 N_GND_M1017_b N_QN_c_1531_n 0.00138285f $X=-0.05 $Y=0 $X2=8.42 $Y2=2.96
cc_217 N_GND_M1017_b QN 0.00299158f $X=-0.05 $Y=0 $X2=8.425 $Y2=2.96
cc_218 N_GND_M1017_b N_Q_c_1603_n 0.0151031f $X=-0.05 $Y=0 $X2=9.28 $Y2=0.825
cc_219 N_GND_c_5_p N_Q_c_1603_n 0.00476261f $X=9.175 $Y=0.17 $X2=9.28 $Y2=0.825
cc_220 N_GND_M1017_b N_Q_c_1605_n 0.0625704f $X=-0.05 $Y=0 $X2=9.395 $Y2=3.16
cc_221 N_GND_M1017_b N_Q_c_1606_n 0.0184431f $X=-0.05 $Y=0 $X2=9.395 $Y2=1.515
cc_222 N_VDD_M1013_b N_RN_M1013_g 0.0266406f $X=-0.05 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_223 N_VDD_c_223_p N_RN_M1013_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_224 N_VDD_c_224_p N_RN_M1013_g 0.00606474f $X=1.915 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_225 N_VDD_c_225_p N_RN_M1013_g 0.00468827f $X=9.175 $Y=6.49 $X2=0.475
+ $Y2=4.585
cc_226 N_VDD_M1013_s N_RN_c_348_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32
+ $Y2=3.33
cc_227 N_VDD_M1013_b N_RN_c_348_n 0.00618364f $X=-0.05 $Y=2.905 $X2=0.32
+ $Y2=3.33
cc_228 N_VDD_c_223_p N_RN_c_348_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_229 N_VDD_M1013_s RN 0.0162774f $X=0.135 $Y=3.085 $X2=0.325 $Y2=3.33
cc_230 N_VDD_c_223_p RN 0.00522047f $X=0.26 $Y=4.135 $X2=0.325 $Y2=3.33
cc_231 N_VDD_M1013_b N_A_110_115#_M1029_g 0.0773537f $X=-0.05 $Y=2.905 $X2=1.425
+ $Y2=5.085
cc_232 N_VDD_c_224_p N_A_110_115#_M1029_g 0.00606474f $X=1.915 $Y=6.507
+ $X2=1.425 $Y2=5.085
cc_233 N_VDD_c_225_p N_A_110_115#_M1029_g 0.00468827f $X=9.175 $Y=6.49 $X2=1.425
+ $Y2=5.085
cc_234 N_VDD_M1013_b N_A_110_115#_M1026_g 0.0795907f $X=-0.05 $Y=2.905 $X2=7.615
+ $Y2=5.085
cc_235 N_VDD_c_235_p N_A_110_115#_M1026_g 0.00606474f $X=7.745 $Y=6.507
+ $X2=7.615 $Y2=5.085
cc_236 N_VDD_c_236_p N_A_110_115#_M1026_g 0.00713292f $X=7.83 $Y=4.475 $X2=7.615
+ $Y2=5.085
cc_237 N_VDD_c_225_p N_A_110_115#_M1026_g 0.00468827f $X=9.175 $Y=6.49 $X2=7.615
+ $Y2=5.085
cc_238 N_VDD_M1013_b N_A_110_115#_c_392_n 0.00549797f $X=-0.05 $Y=2.905 $X2=0.69
+ $Y2=3.455
cc_239 N_VDD_c_224_p N_A_110_115#_c_392_n 0.00757793f $X=1.915 $Y=6.507 $X2=0.69
+ $Y2=3.455
cc_240 N_VDD_c_225_p N_A_110_115#_c_392_n 0.00476261f $X=9.175 $Y=6.49 $X2=0.69
+ $Y2=3.455
cc_241 N_VDD_M1013_b N_A_342_518#_M1000_g 0.085824f $X=-0.05 $Y=2.905 $X2=1.785
+ $Y2=5.085
cc_242 N_VDD_c_224_p N_A_342_518#_M1000_g 0.00606474f $X=1.915 $Y=6.507
+ $X2=1.785 $Y2=5.085
cc_243 N_VDD_c_243_p N_A_342_518#_M1000_g 0.00713292f $X=2 $Y=4.475 $X2=1.785
+ $Y2=5.085
cc_244 N_VDD_c_244_p N_A_342_518#_M1000_g 0.0185359f $X=2.59 $Y=3.795 $X2=1.785
+ $Y2=5.085
cc_245 N_VDD_c_225_p N_A_342_518#_M1000_g 0.00468827f $X=9.175 $Y=6.49 $X2=1.785
+ $Y2=5.085
cc_246 N_VDD_M1013_b N_A_342_518#_c_572_n 0.00442125f $X=-0.05 $Y=2.905 $X2=2.11
+ $Y2=3.1
cc_247 N_VDD_M1021_s N_A_342_518#_c_573_n 0.0125004f $X=2.465 $Y=3.085 $X2=3.295
+ $Y2=3.185
cc_248 N_VDD_M1013_b N_A_342_518#_c_573_n 0.0201537f $X=-0.05 $Y=2.905 $X2=3.295
+ $Y2=3.185
cc_249 N_VDD_c_244_p N_A_342_518#_c_573_n 0.00952036f $X=2.59 $Y=3.795 $X2=3.295
+ $Y2=3.185
cc_250 N_VDD_M1013_b N_A_342_518#_c_576_n 0.00930634f $X=-0.05 $Y=2.905
+ $X2=2.195 $Y2=3.185
cc_251 N_VDD_M1013_b N_A_342_518#_c_577_n 0.00313975f $X=-0.05 $Y=2.905
+ $X2=3.465 $Y2=3.455
cc_252 N_VDD_c_252_p N_A_342_518#_c_577_n 0.0151129f $X=4.255 $Y=6.507 $X2=3.465
+ $Y2=3.455
cc_253 N_VDD_c_225_p N_A_342_518#_c_577_n 0.00958198f $X=9.175 $Y=6.49 $X2=3.465
+ $Y2=3.455
cc_254 N_VDD_M1013_b N_A_342_518#_c_565_n 0.0113251f $X=-0.05 $Y=2.905 $X2=1.94
+ $Y2=2.755
cc_255 N_VDD_M1013_b N_A_342_518#_c_566_n 5.41491e-19 $X=-0.05 $Y=2.905 $X2=2.11
+ $Y2=2.755
cc_256 N_VDD_M1013_b N_D_M1021_g 0.0218296f $X=-0.05 $Y=2.905 $X2=2.805
+ $Y2=4.585
cc_257 N_VDD_c_244_p N_D_M1021_g 0.00713292f $X=2.59 $Y=3.795 $X2=2.805
+ $Y2=4.585
cc_258 N_VDD_c_252_p N_D_M1021_g 0.00606474f $X=4.255 $Y=6.507 $X2=2.805
+ $Y2=4.585
cc_259 N_VDD_c_225_p N_D_M1021_g 0.00468827f $X=9.175 $Y=6.49 $X2=2.805
+ $Y2=4.585
cc_260 N_VDD_M1013_b N_CK_M1023_g 0.020128f $X=-0.05 $Y=2.905 $X2=3.165
+ $Y2=4.585
cc_261 N_VDD_c_252_p N_CK_M1023_g 0.00606474f $X=4.255 $Y=6.507 $X2=3.165
+ $Y2=4.585
cc_262 N_VDD_c_225_p N_CK_M1023_g 0.00468827f $X=9.175 $Y=6.49 $X2=3.165
+ $Y2=4.585
cc_263 N_VDD_M1013_b N_CK_M1011_g 0.020128f $X=-0.05 $Y=2.905 $X2=5.515
+ $Y2=4.585
cc_264 N_VDD_c_264_p N_CK_M1011_g 0.00606474f $X=6.005 $Y=6.507 $X2=5.515
+ $Y2=4.585
cc_265 N_VDD_c_225_p N_CK_M1011_g 0.00468827f $X=9.175 $Y=6.49 $X2=5.515
+ $Y2=4.585
cc_266 N_VDD_M1013_b N_CK_c_678_n 0.00774555f $X=-0.05 $Y=2.905 $X2=6.305
+ $Y2=2.93
cc_267 N_VDD_M1013_b N_CK_M1031_g 0.0237243f $X=-0.05 $Y=2.905 $X2=6.305
+ $Y2=4.585
cc_268 N_VDD_c_268_p N_CK_M1031_g 0.00354579f $X=6.09 $Y=3.455 $X2=6.305
+ $Y2=4.585
cc_269 N_VDD_c_235_p N_CK_M1031_g 0.00606474f $X=7.745 $Y=6.507 $X2=6.305
+ $Y2=4.585
cc_270 N_VDD_c_225_p N_CK_M1031_g 0.00468827f $X=9.175 $Y=6.49 $X2=6.305
+ $Y2=4.585
cc_271 N_VDD_c_268_p N_CK_c_695_n 0.00634153f $X=6.09 $Y=3.455 $X2=6.305
+ $Y2=2.59
cc_272 N_VDD_M1013_b N_CK_c_697_n 6.42499e-19 $X=-0.05 $Y=2.905 $X2=3.225
+ $Y2=2.59
cc_273 N_VDD_M1013_b N_CK_c_698_n 0.0022456f $X=-0.05 $Y=2.905 $X2=5.455
+ $Y2=2.59
cc_274 N_VDD_M1013_b N_CK_c_700_n 0.00302835f $X=-0.05 $Y=2.905 $X2=6.45
+ $Y2=2.59
cc_275 N_VDD_M1013_b N_CK_c_701_n 0.00487135f $X=-0.05 $Y=2.905 $X2=3.225
+ $Y2=2.765
cc_276 N_VDD_M1013_b N_CK_c_708_n 0.00487051f $X=-0.05 $Y=2.905 $X2=5.455
+ $Y2=2.765
cc_277 N_VDD_M1013_b N_A_217_817#_M1028_g 0.0192219f $X=-0.05 $Y=2.905 $X2=4.125
+ $Y2=4.585
cc_278 N_VDD_c_252_p N_A_217_817#_M1028_g 0.00606474f $X=4.255 $Y=6.507
+ $X2=4.125 $Y2=4.585
cc_279 N_VDD_c_279_p N_A_217_817#_M1028_g 0.00354579f $X=4.34 $Y=3.795 $X2=4.125
+ $Y2=4.585
cc_280 N_VDD_c_225_p N_A_217_817#_M1028_g 0.00468827f $X=9.175 $Y=6.49 $X2=4.125
+ $Y2=4.585
cc_281 N_VDD_M1013_b N_A_217_817#_M1006_g 0.0181098f $X=-0.05 $Y=2.905 $X2=4.555
+ $Y2=4.585
cc_282 N_VDD_c_279_p N_A_217_817#_M1006_g 0.00354579f $X=4.34 $Y=3.795 $X2=4.555
+ $Y2=4.585
cc_283 N_VDD_c_264_p N_A_217_817#_M1006_g 0.00606474f $X=6.005 $Y=6.507
+ $X2=4.555 $Y2=4.585
cc_284 N_VDD_c_225_p N_A_217_817#_M1006_g 0.00468827f $X=9.175 $Y=6.49 $X2=4.555
+ $Y2=4.585
cc_285 N_VDD_c_279_p N_A_217_817#_c_909_n 8.24975e-19 $X=4.34 $Y=3.795 $X2=4.48
+ $Y2=2.765
cc_286 N_VDD_M1013_b N_A_217_817#_c_910_n 0.0307874f $X=-0.05 $Y=2.905 $X2=1.21
+ $Y2=4.475
cc_287 N_VDD_c_224_p N_A_217_817#_c_910_n 0.00745733f $X=1.915 $Y=6.507 $X2=1.21
+ $Y2=4.475
cc_288 N_VDD_c_225_p N_A_217_817#_c_910_n 0.00476261f $X=9.175 $Y=6.49 $X2=1.21
+ $Y2=4.475
cc_289 N_VDD_M1013_b N_A_217_817#_c_913_n 0.00424346f $X=-0.05 $Y=2.905
+ $X2=4.295 $Y2=2.765
cc_290 N_VDD_c_279_p N_A_217_817#_c_913_n 0.004428f $X=4.34 $Y=3.795 $X2=4.295
+ $Y2=2.765
cc_291 N_VDD_M1013_b N_A_618_89#_M1030_g 0.0215131f $X=-0.05 $Y=2.905 $X2=3.765
+ $Y2=4.585
cc_292 N_VDD_c_252_p N_A_618_89#_M1030_g 0.00606474f $X=4.255 $Y=6.507 $X2=3.765
+ $Y2=4.585
cc_293 N_VDD_c_225_p N_A_618_89#_M1030_g 0.00468827f $X=9.175 $Y=6.49 $X2=3.765
+ $Y2=4.585
cc_294 N_VDD_M1013_b N_A_618_89#_M1010_g 0.0214821f $X=-0.05 $Y=2.905 $X2=4.915
+ $Y2=4.585
cc_295 N_VDD_c_264_p N_A_618_89#_M1010_g 0.00606474f $X=6.005 $Y=6.507 $X2=4.915
+ $Y2=4.585
cc_296 N_VDD_c_225_p N_A_618_89#_M1010_g 0.00468827f $X=9.175 $Y=6.49 $X2=4.915
+ $Y2=4.585
cc_297 N_VDD_M1013_b N_A_618_89#_c_1072_n 0.00156053f $X=-0.05 $Y=2.905 $X2=6.52
+ $Y2=3.455
cc_298 N_VDD_c_235_p N_A_618_89#_c_1072_n 0.00736239f $X=7.745 $Y=6.507 $X2=6.52
+ $Y2=3.455
cc_299 N_VDD_c_225_p N_A_618_89#_c_1072_n 0.00476261f $X=9.175 $Y=6.49 $X2=6.52
+ $Y2=3.455
cc_300 N_VDD_M1013_b N_A_618_89#_c_1060_n 0.00560125f $X=-0.05 $Y=2.905
+ $X2=6.795 $Y2=3.1
cc_301 N_VDD_M1013_b N_A_618_89#_c_1076_n 0.0139078f $X=-0.05 $Y=2.905 $X2=6.795
+ $Y2=3.185
cc_302 N_VDD_M1013_b N_A_1160_89#_M1009_g 0.0197647f $X=-0.05 $Y=2.905 $X2=5.875
+ $Y2=4.585
cc_303 N_VDD_c_264_p N_A_1160_89#_M1009_g 0.00606474f $X=6.005 $Y=6.507
+ $X2=5.875 $Y2=4.585
cc_304 N_VDD_c_268_p N_A_1160_89#_M1009_g 0.00354579f $X=6.09 $Y=3.455 $X2=5.875
+ $Y2=4.585
cc_305 N_VDD_c_225_p N_A_1160_89#_M1009_g 0.00468827f $X=9.175 $Y=6.49 $X2=5.875
+ $Y2=4.585
cc_306 N_VDD_M1013_b N_A_1160_89#_M1025_g 0.0740454f $X=-0.05 $Y=2.905 $X2=8.635
+ $Y2=5.085
cc_307 N_VDD_c_236_p N_A_1160_89#_M1025_g 0.0067289f $X=7.83 $Y=4.475 $X2=8.635
+ $Y2=5.085
cc_308 N_VDD_c_308_p N_A_1160_89#_M1025_g 0.00606474f $X=8.765 $Y=6.507
+ $X2=8.635 $Y2=5.085
cc_309 N_VDD_c_309_p N_A_1160_89#_M1025_g 0.00354579f $X=8.85 $Y=4.475 $X2=8.635
+ $Y2=5.085
cc_310 N_VDD_c_225_p N_A_1160_89#_M1025_g 0.00468827f $X=9.175 $Y=6.49 $X2=8.635
+ $Y2=5.085
cc_311 N_VDD_M1013_b N_A_1160_89#_c_1236_n 0.00913729f $X=-0.05 $Y=2.905
+ $X2=8.61 $Y2=3.005
cc_312 N_VDD_M1013_b N_A_1160_89#_c_1260_n 0.00618977f $X=-0.05 $Y=2.905
+ $X2=7.04 $Y2=4.475
cc_313 N_VDD_c_235_p N_A_1160_89#_c_1260_n 0.00736239f $X=7.745 $Y=6.507
+ $X2=7.04 $Y2=4.475
cc_314 N_VDD_c_225_p N_A_1160_89#_c_1260_n 0.00476261f $X=9.175 $Y=6.49 $X2=7.04
+ $Y2=4.475
cc_315 N_VDD_M1013_b N_A_1160_89#_c_1263_n 0.0136924f $X=-0.05 $Y=2.905
+ $X2=7.385 $Y2=3.78
cc_316 N_VDD_M1013_b N_A_1160_89#_c_1264_n 0.00887894f $X=-0.05 $Y=2.905
+ $X2=7.125 $Y2=3.78
cc_317 N_VDD_M1013_b N_A_1160_89#_c_1240_n 0.00694317f $X=-0.05 $Y=2.905
+ $X2=7.47 $Y2=3.695
cc_318 N_VDD_M1013_b N_A_998_115#_M1024_g 0.0821041f $X=-0.05 $Y=2.905 $X2=7.255
+ $Y2=5.085
cc_319 N_VDD_c_235_p N_A_998_115#_M1024_g 0.00606474f $X=7.745 $Y=6.507
+ $X2=7.255 $Y2=5.085
cc_320 N_VDD_c_225_p N_A_998_115#_M1024_g 0.00468827f $X=9.175 $Y=6.49 $X2=7.255
+ $Y2=5.085
cc_321 N_VDD_M1013_b N_A_998_115#_c_1406_n 0.00313975f $X=-0.05 $Y=2.905
+ $X2=5.215 $Y2=3.795
cc_322 N_VDD_c_264_p N_A_998_115#_c_1406_n 0.0149205f $X=6.005 $Y=6.507
+ $X2=5.215 $Y2=3.795
cc_323 N_VDD_c_225_p N_A_998_115#_c_1406_n 0.00958198f $X=9.175 $Y=6.49
+ $X2=5.215 $Y2=3.795
cc_324 N_VDD_M1013_b N_A_998_115#_c_1399_n 0.00168314f $X=-0.05 $Y=2.905
+ $X2=4.635 $Y2=1.85
cc_325 N_VDD_M1013_b N_QN_M1002_g 0.0840918f $X=-0.05 $Y=2.905 $X2=9.065
+ $Y2=5.085
cc_326 N_VDD_c_309_p N_QN_M1002_g 0.00354579f $X=8.85 $Y=4.475 $X2=9.065
+ $Y2=5.085
cc_327 N_VDD_c_225_p N_QN_M1002_g 0.00468827f $X=9.175 $Y=6.49 $X2=9.065
+ $Y2=5.085
cc_328 N_VDD_c_328_p N_QN_M1002_g 0.00606474f $X=9.175 $Y=6.44 $X2=9.065
+ $Y2=5.085
cc_329 N_VDD_M1013_b N_QN_c_1531_n 0.0354838f $X=-0.05 $Y=2.905 $X2=8.42
+ $Y2=2.96
cc_330 N_VDD_c_236_p N_QN_c_1531_n 0.0693851f $X=7.83 $Y=4.475 $X2=8.42 $Y2=2.96
cc_331 N_VDD_c_308_p N_QN_c_1531_n 0.00736239f $X=8.765 $Y=6.507 $X2=8.42
+ $Y2=2.96
cc_332 N_VDD_c_225_p N_QN_c_1531_n 0.00476261f $X=9.175 $Y=6.49 $X2=8.42
+ $Y2=2.96
cc_333 N_VDD_M1013_b QN 0.0110801f $X=-0.05 $Y=2.905 $X2=8.425 $Y2=2.96
cc_334 N_VDD_M1013_b N_Q_c_1607_n 0.0342497f $X=-0.05 $Y=2.905 $X2=9.28
+ $Y2=4.475
cc_335 N_VDD_c_225_p N_Q_c_1607_n 0.00476261f $X=9.175 $Y=6.49 $X2=9.28
+ $Y2=4.475
cc_336 N_VDD_c_328_p N_Q_c_1607_n 0.00736239f $X=9.175 $Y=6.44 $X2=9.28
+ $Y2=4.475
cc_337 N_VDD_M1013_b N_Q_c_1605_n 0.0127419f $X=-0.05 $Y=2.905 $X2=9.395
+ $Y2=3.16
cc_338 N_VDD_M1013_b Q 0.0106945f $X=-0.05 $Y=2.905 $X2=9.275 $Y2=3.33
cc_339 N_VDD_M1013_b N_Q_c_1612_n 0.0207082f $X=-0.05 $Y=2.905 $X2=9.275
+ $Y2=3.33
cc_340 RN N_A_110_115#_M1013_d 0.00414531f $X=0.325 $Y=3.33 $X2=0.55 $Y2=3.085
cc_341 N_RN_c_345_n N_A_110_115#_M1029_g 0.00293469f $X=0.475 $Y=2.47 $X2=1.425
+ $Y2=5.085
cc_342 N_RN_M1013_g N_A_110_115#_c_392_n 0.0104129f $X=0.475 $Y=4.585 $X2=0.69
+ $Y2=3.455
cc_343 N_RN_c_348_n N_A_110_115#_c_392_n 0.0282684f $X=0.32 $Y=3.33 $X2=0.69
+ $Y2=3.455
cc_344 RN N_A_110_115#_c_392_n 0.00974028f $X=0.325 $Y=3.33 $X2=0.69 $Y2=3.455
cc_345 N_RN_M1017_g N_A_110_115#_c_393_n 0.0139885f $X=0.475 $Y=1.075 $X2=0.87
+ $Y2=2.655
cc_346 N_RN_c_345_n N_A_110_115#_c_393_n 0.00370757f $X=0.475 $Y=2.47 $X2=0.87
+ $Y2=2.655
cc_347 N_RN_M1013_g N_A_110_115#_c_393_n 0.00363549f $X=0.475 $Y=4.585 $X2=0.87
+ $Y2=2.655
cc_348 N_RN_c_347_n N_A_110_115#_c_393_n 0.0248372f $X=0.32 $Y=2.305 $X2=0.87
+ $Y2=2.655
cc_349 N_RN_c_348_n N_A_110_115#_c_393_n 0.0072511f $X=0.32 $Y=3.33 $X2=0.87
+ $Y2=2.655
cc_350 N_RN_M1017_g N_A_110_115#_c_396_n 0.00375199f $X=0.475 $Y=1.075 $X2=0.955
+ $Y2=1.59
cc_351 N_RN_c_345_n N_A_110_115#_c_396_n 0.00143285f $X=0.475 $Y=2.47 $X2=0.955
+ $Y2=1.59
cc_352 N_RN_c_347_n N_A_110_115#_c_396_n 3.54179e-19 $X=0.32 $Y=2.305 $X2=0.955
+ $Y2=1.59
cc_353 N_RN_c_345_n N_A_110_115#_c_397_n 0.00191737f $X=0.475 $Y=2.47 $X2=0.87
+ $Y2=2.74
cc_354 N_RN_M1013_g N_A_110_115#_c_397_n 0.00385986f $X=0.475 $Y=4.585 $X2=0.87
+ $Y2=2.74
cc_355 N_RN_c_347_n N_A_110_115#_c_397_n 7.08415e-19 $X=0.32 $Y=2.305 $X2=0.87
+ $Y2=2.74
cc_356 N_RN_c_348_n N_A_110_115#_c_397_n 0.0113366f $X=0.32 $Y=3.33 $X2=0.87
+ $Y2=2.74
cc_357 N_RN_M1017_g N_A_110_115#_c_415_n 0.00503705f $X=0.475 $Y=1.075 $X2=1.425
+ $Y2=1.59
cc_358 N_RN_M1013_g N_A_217_817#_c_910_n 0.007087f $X=0.475 $Y=4.585 $X2=1.21
+ $Y2=4.475
cc_359 RN N_A_217_817#_c_910_n 9.10636e-19 $X=0.325 $Y=3.33 $X2=1.21 $Y2=4.475
cc_360 N_A_110_115#_c_398_n N_A_342_518#_M1027_d 0.00558831f $X=7.665 $Y=1.48
+ $X2=3.24 $Y2=0.575
cc_361 N_A_110_115#_c_378_n N_A_342_518#_M1001_g 0.0731012f $X=1.425 $Y=1.425
+ $X2=1.855 $Y2=0.945
cc_362 N_A_110_115#_c_398_n N_A_342_518#_M1001_g 0.0124017f $X=7.665 $Y=1.48
+ $X2=1.855 $Y2=0.945
cc_363 N_A_110_115#_c_398_n N_A_342_518#_c_557_n 0.025935f $X=7.665 $Y=1.48
+ $X2=3.28 $Y2=1.765
cc_364 N_A_110_115#_c_398_n N_A_342_518#_c_559_n 0.00359329f $X=7.665 $Y=1.48
+ $X2=2.195 $Y2=1.765
cc_365 N_A_110_115#_c_398_n N_A_342_518#_c_561_n 0.0151351f $X=7.665 $Y=1.48
+ $X2=3.365 $Y2=1.68
cc_366 N_A_110_115#_M1029_g N_A_342_518#_c_565_n 0.21674f $X=1.425 $Y=5.085
+ $X2=1.94 $Y2=2.755
cc_367 N_A_110_115#_M1029_g N_A_342_518#_c_566_n 9.03256e-19 $X=1.425 $Y=5.085
+ $X2=2.11 $Y2=2.755
cc_368 N_A_110_115#_c_398_n N_A_342_518#_c_590_n 0.0254135f $X=7.665 $Y=1.48
+ $X2=3.457 $Y2=1.415
cc_369 N_A_110_115#_c_398_n N_D_M1003_g 0.0116357f $X=7.665 $Y=1.48 $X2=2.805
+ $Y2=1.075
cc_370 N_A_110_115#_c_398_n N_CK_c_680_n 0.01159f $X=7.665 $Y=1.48 $X2=6.332
+ $Y2=1.685
cc_371 N_A_110_115#_c_398_n N_CK_c_685_n 0.00107886f $X=7.665 $Y=1.48 $X2=6.332
+ $Y2=1.835
cc_372 N_A_110_115#_c_398_n N_CK_c_687_n 0.00496158f $X=7.665 $Y=1.48 $X2=3.705
+ $Y2=1.85
cc_373 N_A_110_115#_c_398_n N_CK_c_688_n 8.06574e-19 $X=7.665 $Y=1.48 $X2=3.705
+ $Y2=1.85
cc_374 N_A_110_115#_c_398_n N_CK_c_689_n 0.00118606f $X=7.665 $Y=1.48 $X2=4.975
+ $Y2=1.85
cc_375 N_A_110_115#_c_398_n N_CK_c_690_n 8.06574e-19 $X=7.665 $Y=1.48 $X2=4.975
+ $Y2=1.85
cc_376 N_A_110_115#_c_398_n N_CK_c_702_n 0.0106495f $X=7.665 $Y=1.48 $X2=3.705
+ $Y2=1.685
cc_377 N_A_110_115#_c_398_n N_CK_c_705_n 0.00177838f $X=7.665 $Y=1.48 $X2=4.975
+ $Y2=1.685
cc_378 N_A_110_115#_c_398_n N_A_217_817#_M1022_g 0.0104272f $X=7.665 $Y=1.48
+ $X2=4.125 $Y2=1.075
cc_379 N_A_110_115#_c_398_n N_A_217_817#_M1019_g 0.00491871f $X=7.665 $Y=1.48
+ $X2=4.555 $Y2=1.075
cc_380 N_A_110_115#_c_398_n N_A_217_817#_c_907_n 2.42482e-19 $X=7.665 $Y=1.48
+ $X2=4.48 $Y2=1.85
cc_381 N_A_110_115#_M1029_g N_A_217_817#_c_910_n 0.0742296f $X=1.425 $Y=5.085
+ $X2=1.21 $Y2=4.475
cc_382 N_A_110_115#_c_392_n N_A_217_817#_c_910_n 0.140442f $X=0.69 $Y=3.455
+ $X2=1.21 $Y2=4.475
cc_383 N_A_110_115#_c_393_n N_A_217_817#_c_910_n 0.0413763f $X=0.87 $Y=2.655
+ $X2=1.21 $Y2=4.475
cc_384 N_A_110_115#_c_397_n N_A_217_817#_c_910_n 0.0134441f $X=0.87 $Y=2.74
+ $X2=1.21 $Y2=4.475
cc_385 N_A_110_115#_M1029_g N_A_217_817#_c_911_n 0.0166119f $X=1.425 $Y=5.085
+ $X2=1.555 $Y2=2.02
cc_386 N_A_110_115#_c_398_n N_A_217_817#_c_911_n 0.00400792f $X=7.665 $Y=1.48
+ $X2=1.555 $Y2=2.02
cc_387 N_A_110_115#_c_407_n N_A_217_817#_c_911_n 0.0022406f $X=1.375 $Y=1.48
+ $X2=1.555 $Y2=2.02
cc_388 N_A_110_115#_c_409_n N_A_217_817#_c_911_n 0.00125872f $X=1.23 $Y=1.48
+ $X2=1.555 $Y2=2.02
cc_389 N_A_110_115#_c_415_n N_A_217_817#_c_911_n 0.00146789f $X=1.425 $Y=1.59
+ $X2=1.555 $Y2=2.02
cc_390 N_A_110_115#_c_393_n N_A_217_817#_c_912_n 0.0141418f $X=0.87 $Y=2.655
+ $X2=1.295 $Y2=2.02
cc_391 N_A_110_115#_c_394_n N_A_217_817#_c_912_n 0.0010034f $X=1.145 $Y=1.59
+ $X2=1.295 $Y2=2.02
cc_392 N_A_110_115#_c_407_n N_A_217_817#_c_912_n 0.00102018f $X=1.375 $Y=1.48
+ $X2=1.295 $Y2=2.02
cc_393 N_A_110_115#_c_409_n N_A_217_817#_c_912_n 0.0112658f $X=1.23 $Y=1.48
+ $X2=1.295 $Y2=2.02
cc_394 N_A_110_115#_c_415_n N_A_217_817#_c_912_n 0.00170324f $X=1.425 $Y=1.59
+ $X2=1.295 $Y2=2.02
cc_395 N_A_110_115#_c_398_n N_A_217_817#_c_914_n 0.183791f $X=7.665 $Y=1.48
+ $X2=4.06 $Y2=1.85
cc_396 N_A_110_115#_M1029_g N_A_217_817#_c_915_n 0.00354431f $X=1.425 $Y=5.085
+ $X2=1.785 $Y2=1.85
cc_397 N_A_110_115#_c_393_n N_A_217_817#_c_915_n 0.00409794f $X=0.87 $Y=2.655
+ $X2=1.785 $Y2=1.85
cc_398 N_A_110_115#_c_398_n N_A_217_817#_c_915_n 0.0254191f $X=7.665 $Y=1.48
+ $X2=1.785 $Y2=1.85
cc_399 N_A_110_115#_c_409_n N_A_217_817#_c_915_n 4.96965e-19 $X=1.23 $Y=1.48
+ $X2=1.785 $Y2=1.85
cc_400 N_A_110_115#_c_415_n N_A_217_817#_c_915_n 3.4709e-19 $X=1.425 $Y=1.59
+ $X2=1.785 $Y2=1.85
cc_401 N_A_110_115#_c_398_n N_A_217_817#_c_960_n 0.0259207f $X=7.665 $Y=1.48
+ $X2=4.205 $Y2=1.85
cc_402 N_A_110_115#_c_398_n N_A_217_817#_c_916_n 0.00546464f $X=7.665 $Y=1.48
+ $X2=4.205 $Y2=1.85
cc_403 N_A_110_115#_c_378_n N_A_217_817#_c_918_n 0.00816167f $X=1.425 $Y=1.425
+ $X2=1.64 $Y2=0.825
cc_404 N_A_110_115#_c_393_n N_A_217_817#_c_918_n 0.00308284f $X=0.87 $Y=2.655
+ $X2=1.64 $Y2=0.825
cc_405 N_A_110_115#_c_398_n N_A_217_817#_c_918_n 0.0227937f $X=7.665 $Y=1.48
+ $X2=1.64 $Y2=0.825
cc_406 N_A_110_115#_c_407_n N_A_217_817#_c_918_n 0.00209779f $X=1.375 $Y=1.48
+ $X2=1.64 $Y2=0.825
cc_407 N_A_110_115#_c_409_n N_A_217_817#_c_918_n 0.0180047f $X=1.23 $Y=1.48
+ $X2=1.64 $Y2=0.825
cc_408 N_A_110_115#_c_398_n N_A_618_89#_M1005_d 0.00421798f $X=7.665 $Y=1.48
+ $X2=6.38 $Y2=0.575
cc_409 N_A_110_115#_c_398_n N_A_618_89#_c_1037_n 0.0102209f $X=7.665 $Y=1.48
+ $X2=3.165 $Y2=1.685
cc_410 N_A_110_115#_c_398_n N_A_618_89#_c_1051_n 0.0115848f $X=7.665 $Y=1.48
+ $X2=6.435 $Y2=1.85
cc_411 N_A_110_115#_c_398_n N_A_618_89#_c_1053_n 0.00232964f $X=7.665 $Y=1.48
+ $X2=5.455 $Y2=1.85
cc_412 N_A_110_115#_c_398_n N_A_618_89#_c_1054_n 0.025543f $X=7.665 $Y=1.48
+ $X2=6.52 $Y2=0.825
cc_413 N_A_110_115#_c_398_n N_A_618_89#_c_1062_n 5.01657e-19 $X=7.665 $Y=1.48
+ $X2=6.795 $Y2=2.19
cc_414 N_A_110_115#_c_398_n N_A_618_89#_c_1063_n 0.0103799f $X=7.665 $Y=1.48
+ $X2=5.455 $Y2=1.685
cc_415 N_A_110_115#_c_398_n N_A_1160_89#_M1018_g 0.0100216f $X=7.665 $Y=1.48
+ $X2=5.875 $Y2=1.075
cc_416 N_A_110_115#_c_417_n N_A_1160_89#_M1012_g 0.00315793f $X=7.81 $Y=1.59
+ $X2=8.635 $Y2=0.945
cc_417 N_A_110_115#_c_417_n N_A_1160_89#_c_1234_n 0.00151565f $X=7.81 $Y=1.59
+ $X2=8.61 $Y2=1.8
cc_418 N_A_110_115#_M1026_g N_A_1160_89#_c_1263_n 0.0100206f $X=7.615 $Y=5.085
+ $X2=7.385 $Y2=3.78
cc_419 N_A_110_115#_M1026_g N_A_1160_89#_c_1237_n 0.0157637f $X=7.615 $Y=5.085
+ $X2=7.47 $Y2=0.825
cc_420 N_A_110_115#_c_384_n N_A_1160_89#_c_1237_n 0.00353845f $X=7.685 $Y=1.425
+ $X2=7.47 $Y2=0.825
cc_421 N_A_110_115#_c_398_n N_A_1160_89#_c_1237_n 0.0244886f $X=7.665 $Y=1.48
+ $X2=7.47 $Y2=0.825
cc_422 N_A_110_115#_c_411_n N_A_1160_89#_c_1237_n 0.00222483f $X=7.81 $Y=1.48
+ $X2=7.47 $Y2=0.825
cc_423 N_A_110_115#_c_413_n N_A_1160_89#_c_1237_n 0.0236844f $X=7.81 $Y=1.48
+ $X2=7.47 $Y2=0.825
cc_424 N_A_110_115#_c_417_n N_A_1160_89#_c_1237_n 0.00632512f $X=7.81 $Y=1.59
+ $X2=7.47 $Y2=0.825
cc_425 N_A_110_115#_M1026_g N_A_1160_89#_c_1240_n 0.0612926f $X=7.615 $Y=5.085
+ $X2=7.47 $Y2=3.695
cc_426 N_A_110_115#_M1026_g N_A_1160_89#_c_1241_n 0.00121075f $X=7.615 $Y=5.085
+ $X2=7.47 $Y2=2.19
cc_427 N_A_110_115#_M1026_g N_A_1160_89#_c_1242_n 0.00787213f $X=7.615 $Y=5.085
+ $X2=8.375 $Y2=2.19
cc_428 N_A_110_115#_c_398_n N_A_1160_89#_c_1242_n 0.0171303f $X=7.665 $Y=1.48
+ $X2=8.375 $Y2=2.19
cc_429 N_A_110_115#_c_411_n N_A_1160_89#_c_1242_n 0.0141753f $X=7.81 $Y=1.48
+ $X2=8.375 $Y2=2.19
cc_430 N_A_110_115#_c_413_n N_A_1160_89#_c_1242_n 0.00159971f $X=7.81 $Y=1.48
+ $X2=8.375 $Y2=2.19
cc_431 N_A_110_115#_c_417_n N_A_1160_89#_c_1242_n 0.00144106f $X=7.81 $Y=1.59
+ $X2=8.375 $Y2=2.19
cc_432 N_A_110_115#_M1026_g N_A_1160_89#_c_1246_n 0.0120256f $X=7.615 $Y=5.085
+ $X2=8.52 $Y2=2.19
cc_433 N_A_110_115#_c_398_n N_A_1160_89#_c_1246_n 0.00118947f $X=7.665 $Y=1.48
+ $X2=8.52 $Y2=2.19
cc_434 N_A_110_115#_c_411_n N_A_1160_89#_c_1246_n 0.00102994f $X=7.81 $Y=1.48
+ $X2=8.52 $Y2=2.19
cc_435 N_A_110_115#_c_413_n N_A_1160_89#_c_1246_n 0.00521974f $X=7.81 $Y=1.48
+ $X2=8.52 $Y2=2.19
cc_436 N_A_110_115#_c_417_n N_A_1160_89#_c_1246_n 0.00329212f $X=7.81 $Y=1.59
+ $X2=8.52 $Y2=2.19
cc_437 N_A_110_115#_M1026_g N_A_1160_89#_c_1248_n 0.0050953f $X=7.615 $Y=5.085
+ $X2=8.52 $Y2=2.19
cc_438 N_A_110_115#_c_398_n N_A_998_115#_M1015_d 0.0051762f $X=7.665 $Y=1.48
+ $X2=4.99 $Y2=0.575
cc_439 N_A_110_115#_c_384_n N_A_998_115#_M1007_g 0.0219629f $X=7.685 $Y=1.425
+ $X2=7.255 $Y2=0.945
cc_440 N_A_110_115#_c_398_n N_A_998_115#_M1007_g 0.0123745f $X=7.665 $Y=1.48
+ $X2=7.255 $Y2=0.945
cc_441 N_A_110_115#_c_417_n N_A_998_115#_M1007_g 0.142765f $X=7.81 $Y=1.59
+ $X2=7.255 $Y2=0.945
cc_442 N_A_110_115#_M1026_g N_A_998_115#_c_1390_n 0.142765f $X=7.615 $Y=5.085
+ $X2=7.255 $Y2=2.015
cc_443 N_A_110_115#_c_398_n N_A_998_115#_c_1390_n 0.00181397f $X=7.665 $Y=1.48
+ $X2=7.255 $Y2=2.015
cc_444 N_A_110_115#_c_398_n N_A_998_115#_c_1416_n 0.0537388f $X=7.665 $Y=1.48
+ $X2=5.045 $Y2=1.43
cc_445 N_A_110_115#_c_398_n N_A_998_115#_c_1417_n 0.0129425f $X=7.665 $Y=1.48
+ $X2=4.72 $Y2=1.43
cc_446 N_A_110_115#_c_398_n N_A_998_115#_c_1396_n 0.183754f $X=7.665 $Y=1.48
+ $X2=6.985 $Y2=1.85
cc_447 N_A_110_115#_c_398_n N_A_998_115#_c_1398_n 0.0252354f $X=7.665 $Y=1.48
+ $X2=4.78 $Y2=1.85
cc_448 N_A_110_115#_c_398_n N_A_998_115#_c_1399_n 0.00616681f $X=7.665 $Y=1.48
+ $X2=4.635 $Y2=1.85
cc_449 N_A_110_115#_c_398_n N_A_998_115#_c_1400_n 0.0259677f $X=7.665 $Y=1.48
+ $X2=7.13 $Y2=1.85
cc_450 N_A_110_115#_c_398_n N_A_998_115#_c_1401_n 0.00340149f $X=7.665 $Y=1.48
+ $X2=7.13 $Y2=1.85
cc_451 N_A_110_115#_c_417_n N_A_998_115#_c_1401_n 3.53041e-19 $X=7.81 $Y=1.59
+ $X2=7.13 $Y2=1.85
cc_452 N_A_110_115#_c_384_n N_QN_c_1521_n 0.0082109f $X=7.685 $Y=1.425 $X2=8.42
+ $Y2=0.825
cc_453 N_A_110_115#_c_411_n N_QN_c_1521_n 0.00696569f $X=7.81 $Y=1.48 $X2=8.42
+ $Y2=0.825
cc_454 N_A_110_115#_c_413_n N_QN_c_1521_n 0.00993531f $X=7.81 $Y=1.48 $X2=8.42
+ $Y2=0.825
cc_455 N_A_110_115#_c_417_n N_QN_c_1521_n 0.00254684f $X=7.81 $Y=1.59 $X2=8.42
+ $Y2=0.825
cc_456 N_A_110_115#_M1026_g N_QN_c_1526_n 0.00427758f $X=7.615 $Y=5.085
+ $X2=8.505 $Y2=1.85
cc_457 N_A_110_115#_M1026_g N_QN_c_1528_n 0.00423893f $X=7.615 $Y=5.085
+ $X2=8.505 $Y2=2.765
cc_458 N_A_110_115#_M1026_g N_QN_c_1531_n 0.0317573f $X=7.615 $Y=5.085 $X2=8.42
+ $Y2=2.96
cc_459 N_A_110_115#_M1026_g QN 0.00472165f $X=7.615 $Y=5.085 $X2=8.425 $Y2=2.96
cc_460 N_A_110_115#_c_398_n A_576_115# 0.00911585f $X=7.665 $Y=1.48 $X2=2.88
+ $Y2=0.575
cc_461 N_A_110_115#_c_398_n A_768_115# 0.0100396f $X=7.665 $Y=1.48 $X2=3.84
+ $Y2=0.575
cc_462 N_A_110_115#_c_398_n A_926_115# 0.00106636f $X=7.665 $Y=1.48 $X2=4.63
+ $Y2=0.575
cc_463 N_A_110_115#_c_398_n A_1118_115# 0.00917995f $X=7.665 $Y=1.48 $X2=5.59
+ $Y2=0.575
cc_464 N_A_342_518#_c_556_n N_D_M1003_g 0.0129746f $X=2.11 $Y=2.59 $X2=2.805
+ $Y2=1.075
cc_465 N_A_342_518#_c_557_n N_D_M1003_g 0.0122665f $X=3.28 $Y=1.765 $X2=2.805
+ $Y2=1.075
cc_466 N_A_342_518#_c_572_n N_D_M1021_g 0.00419666f $X=2.11 $Y=3.1 $X2=2.805
+ $Y2=4.585
cc_467 N_A_342_518#_c_573_n N_D_M1021_g 0.0211478f $X=3.295 $Y=3.185 $X2=2.805
+ $Y2=4.585
cc_468 N_A_342_518#_c_565_n N_D_M1021_g 0.00397893f $X=1.94 $Y=2.755 $X2=2.805
+ $Y2=4.585
cc_469 N_A_342_518#_c_566_n N_D_M1021_g 0.00576391f $X=2.11 $Y=2.755 $X2=2.805
+ $Y2=4.585
cc_470 N_A_342_518#_c_556_n D 0.0055149f $X=2.11 $Y=2.59 $X2=2.865 $Y2=2.22
cc_471 N_A_342_518#_c_557_n D 0.00200799f $X=3.28 $Y=1.765 $X2=2.865 $Y2=2.22
cc_472 N_A_342_518#_c_556_n N_D_c_643_n 0.00613892f $X=2.11 $Y=2.59 $X2=2.865
+ $Y2=2.22
cc_473 N_A_342_518#_c_557_n N_D_c_643_n 0.0086486f $X=3.28 $Y=1.765 $X2=2.865
+ $Y2=2.22
cc_474 N_A_342_518#_c_557_n N_D_c_644_n 0.00207628f $X=3.28 $Y=1.765 $X2=2.865
+ $Y2=2.22
cc_475 N_A_342_518#_c_573_n N_CK_M1023_g 0.0153421f $X=3.295 $Y=3.185 $X2=3.165
+ $Y2=4.585
cc_476 N_A_342_518#_c_557_n N_CK_c_686_n 0.0019742f $X=3.28 $Y=1.765 $X2=3.62
+ $Y2=2.59
cc_477 N_A_342_518#_c_573_n N_CK_c_686_n 0.00883015f $X=3.295 $Y=3.185 $X2=3.62
+ $Y2=2.59
cc_478 N_A_342_518#_c_557_n N_CK_c_687_n 0.012316f $X=3.28 $Y=1.765 $X2=3.705
+ $Y2=1.85
cc_479 N_A_342_518#_c_590_n N_CK_c_687_n 5.28119e-19 $X=3.457 $Y=1.415 $X2=3.705
+ $Y2=1.85
cc_480 N_A_342_518#_c_557_n N_CK_c_688_n 9.45214e-19 $X=3.28 $Y=1.765 $X2=3.705
+ $Y2=1.85
cc_481 N_A_342_518#_c_590_n N_CK_c_688_n 0.00170561f $X=3.457 $Y=1.415 $X2=3.705
+ $Y2=1.85
cc_482 N_A_342_518#_c_573_n N_CK_c_693_n 0.00601583f $X=3.295 $Y=3.185 $X2=5.31
+ $Y2=2.59
cc_483 N_A_342_518#_c_573_n N_CK_c_694_n 0.00409373f $X=3.295 $Y=3.185 $X2=3.37
+ $Y2=2.59
cc_484 N_A_342_518#_c_557_n N_CK_c_697_n 0.00224444f $X=3.28 $Y=1.765 $X2=3.225
+ $Y2=2.59
cc_485 N_A_342_518#_c_573_n N_CK_c_697_n 0.0101098f $X=3.295 $Y=3.185 $X2=3.225
+ $Y2=2.59
cc_486 N_A_342_518#_c_573_n N_CK_c_701_n 0.00150627f $X=3.295 $Y=3.185 $X2=3.225
+ $Y2=2.765
cc_487 N_A_342_518#_c_561_n N_CK_c_702_n 0.00464203f $X=3.365 $Y=1.68 $X2=3.705
+ $Y2=1.685
cc_488 N_A_342_518#_c_590_n N_CK_c_702_n 0.00545632f $X=3.457 $Y=1.415 $X2=3.705
+ $Y2=1.685
cc_489 N_A_342_518#_c_566_n N_A_217_817#_c_910_n 0.00998126f $X=2.11 $Y=2.755
+ $X2=1.21 $Y2=4.475
cc_490 N_A_342_518#_M1001_g N_A_217_817#_c_911_n 0.00170001f $X=1.855 $Y=0.945
+ $X2=1.555 $Y2=2.02
cc_491 N_A_342_518#_c_556_n N_A_217_817#_c_911_n 0.00898241f $X=2.11 $Y=2.59
+ $X2=1.555 $Y2=2.02
cc_492 N_A_342_518#_c_565_n N_A_217_817#_c_911_n 5.21343e-19 $X=1.94 $Y=2.755
+ $X2=1.555 $Y2=2.02
cc_493 N_A_342_518#_M1001_g N_A_217_817#_c_914_n 0.0109775f $X=1.855 $Y=0.945
+ $X2=4.06 $Y2=1.85
cc_494 N_A_342_518#_c_556_n N_A_217_817#_c_914_n 0.0148809f $X=2.11 $Y=2.59
+ $X2=4.06 $Y2=1.85
cc_495 N_A_342_518#_c_557_n N_A_217_817#_c_914_n 0.0477939f $X=3.28 $Y=1.765
+ $X2=4.06 $Y2=1.85
cc_496 N_A_342_518#_c_559_n N_A_217_817#_c_914_n 0.00452388f $X=2.195 $Y=1.765
+ $X2=4.06 $Y2=1.85
cc_497 N_A_342_518#_c_590_n N_A_217_817#_c_914_n 8.61924e-19 $X=3.457 $Y=1.415
+ $X2=4.06 $Y2=1.85
cc_498 N_A_342_518#_M1001_g N_A_217_817#_c_915_n 0.00225183f $X=1.855 $Y=0.945
+ $X2=1.785 $Y2=1.85
cc_499 N_A_342_518#_c_556_n N_A_217_817#_c_915_n 7.31874e-19 $X=2.11 $Y=2.59
+ $X2=1.785 $Y2=1.85
cc_500 N_A_342_518#_c_559_n N_A_217_817#_c_915_n 7.73026e-19 $X=2.195 $Y=1.765
+ $X2=1.785 $Y2=1.85
cc_501 N_A_342_518#_c_565_n N_A_217_817#_c_915_n 0.00124753f $X=1.94 $Y=2.755
+ $X2=1.785 $Y2=1.85
cc_502 N_A_342_518#_M1001_g N_A_217_817#_c_918_n 0.0115512f $X=1.855 $Y=0.945
+ $X2=1.64 $Y2=0.825
cc_503 N_A_342_518#_c_556_n N_A_217_817#_c_918_n 0.0033876f $X=2.11 $Y=2.59
+ $X2=1.64 $Y2=0.825
cc_504 N_A_342_518#_c_559_n N_A_217_817#_c_918_n 0.00785026f $X=2.195 $Y=1.765
+ $X2=1.64 $Y2=0.825
cc_505 N_A_342_518#_c_557_n N_A_618_89#_c_1037_n 0.0022787f $X=3.28 $Y=1.765
+ $X2=3.165 $Y2=1.685
cc_506 N_A_342_518#_c_590_n N_A_618_89#_c_1037_n 0.0060945f $X=3.457 $Y=1.415
+ $X2=3.165 $Y2=1.685
cc_507 N_A_342_518#_c_557_n N_A_618_89#_c_1040_n 0.00324141f $X=3.28 $Y=1.765
+ $X2=3.285 $Y2=2.225
cc_508 N_A_342_518#_c_557_n N_A_618_89#_c_1048_n 0.00993431f $X=3.28 $Y=1.765
+ $X2=3.285 $Y2=1.76
cc_509 N_A_342_518#_c_573_n A_576_617# 0.00732587f $X=3.295 $Y=3.185 $X2=2.88
+ $Y2=3.085
cc_510 D N_CK_c_687_n 0.00551577f $X=2.865 $Y=2.22 $X2=3.705 $Y2=1.85
cc_511 N_D_c_643_n N_CK_c_687_n 0.00478177f $X=2.865 $Y=2.22 $X2=3.705 $Y2=1.85
cc_512 N_D_c_644_n N_CK_c_687_n 2.89615e-19 $X=2.865 $Y=2.22 $X2=3.705 $Y2=1.85
cc_513 N_D_M1021_g N_CK_c_694_n 0.00515433f $X=2.805 $Y=4.585 $X2=3.37 $Y2=2.59
cc_514 D N_CK_c_694_n 0.00375733f $X=2.865 $Y=2.22 $X2=3.37 $Y2=2.59
cc_515 N_D_M1021_g N_CK_c_697_n 0.00494364f $X=2.805 $Y=4.585 $X2=3.225 $Y2=2.59
cc_516 N_D_M1021_g N_CK_c_701_n 0.21604f $X=2.805 $Y=4.585 $X2=3.225 $Y2=2.765
cc_517 N_D_M1003_g N_A_217_817#_c_914_n 0.0030176f $X=2.805 $Y=1.075 $X2=4.06
+ $Y2=1.85
cc_518 D N_A_217_817#_c_914_n 0.0353362f $X=2.865 $Y=2.22 $X2=4.06 $Y2=1.85
cc_519 N_D_c_643_n N_A_217_817#_c_914_n 0.00111625f $X=2.865 $Y=2.22 $X2=4.06
+ $Y2=1.85
cc_520 N_D_c_644_n N_A_217_817#_c_914_n 7.9412e-19 $X=2.865 $Y=2.22 $X2=4.06
+ $Y2=1.85
cc_521 N_D_M1003_g N_A_618_89#_c_1037_n 0.0846533f $X=2.805 $Y=1.075 $X2=3.165
+ $Y2=1.685
cc_522 N_D_M1003_g N_A_618_89#_c_1040_n 0.00932846f $X=2.805 $Y=1.075 $X2=3.285
+ $Y2=2.225
cc_523 D N_A_618_89#_c_1040_n 0.00342011f $X=2.865 $Y=2.22 $X2=3.285 $Y2=2.225
cc_524 N_D_c_643_n N_A_618_89#_c_1040_n 0.00164409f $X=2.865 $Y=2.22 $X2=3.285
+ $Y2=2.225
cc_525 N_D_c_644_n N_A_618_89#_c_1040_n 0.0210215f $X=2.865 $Y=2.22 $X2=3.285
+ $Y2=2.225
cc_526 D N_A_618_89#_c_1042_n 4.62757e-19 $X=2.865 $Y=2.22 $X2=3.36 $Y2=2.3
cc_527 N_CK_c_687_n N_A_217_817#_M1022_g 0.00109079f $X=3.705 $Y=1.85 $X2=4.125
+ $Y2=1.075
cc_528 N_CK_c_702_n N_A_217_817#_M1022_g 0.0483944f $X=3.705 $Y=1.685 $X2=4.125
+ $Y2=1.075
cc_529 N_CK_c_689_n N_A_217_817#_M1019_g 3.67139e-19 $X=4.975 $Y=1.85 $X2=4.555
+ $Y2=1.075
cc_530 N_CK_c_705_n N_A_217_817#_M1019_g 0.0473482f $X=4.975 $Y=1.685 $X2=4.555
+ $Y2=1.075
cc_531 N_CK_c_688_n N_A_217_817#_c_905_n 0.0483944f $X=3.705 $Y=1.85 $X2=4.2
+ $Y2=1.85
cc_532 N_CK_c_693_n N_A_217_817#_c_906_n 0.00679967f $X=5.31 $Y=2.59 $X2=4.2
+ $Y2=2.765
cc_533 N_CK_c_690_n N_A_217_817#_c_907_n 0.0473482f $X=4.975 $Y=1.85 $X2=4.48
+ $Y2=1.85
cc_534 N_CK_c_693_n N_A_217_817#_c_909_n 0.00772879f $X=5.31 $Y=2.59 $X2=4.48
+ $Y2=2.765
cc_535 N_CK_c_686_n N_A_217_817#_c_913_n 0.00401809f $X=3.62 $Y=2.59 $X2=4.295
+ $Y2=2.765
cc_536 N_CK_c_687_n N_A_217_817#_c_913_n 0.0203851f $X=3.705 $Y=1.85 $X2=4.295
+ $Y2=2.765
cc_537 N_CK_c_688_n N_A_217_817#_c_913_n 7.30049e-19 $X=3.705 $Y=1.85 $X2=4.295
+ $Y2=2.765
cc_538 N_CK_c_693_n N_A_217_817#_c_913_n 0.0206884f $X=5.31 $Y=2.59 $X2=4.295
+ $Y2=2.765
cc_539 N_CK_c_686_n N_A_217_817#_c_914_n 0.00443421f $X=3.62 $Y=2.59 $X2=4.06
+ $Y2=1.85
cc_540 N_CK_c_687_n N_A_217_817#_c_914_n 0.0149977f $X=3.705 $Y=1.85 $X2=4.06
+ $Y2=1.85
cc_541 N_CK_c_688_n N_A_217_817#_c_914_n 0.00383172f $X=3.705 $Y=1.85 $X2=4.06
+ $Y2=1.85
cc_542 N_CK_c_694_n N_A_217_817#_c_914_n 0.0126164f $X=3.37 $Y=2.59 $X2=4.06
+ $Y2=1.85
cc_543 N_CK_c_697_n N_A_217_817#_c_914_n 7.12046e-19 $X=3.225 $Y=2.59 $X2=4.06
+ $Y2=1.85
cc_544 N_CK_c_687_n N_A_217_817#_c_960_n 0.00143592f $X=3.705 $Y=1.85 $X2=4.205
+ $Y2=1.85
cc_545 N_CK_c_688_n N_A_217_817#_c_960_n 3.3031e-19 $X=3.705 $Y=1.85 $X2=4.205
+ $Y2=1.85
cc_546 N_CK_c_693_n N_A_217_817#_c_960_n 0.0129652f $X=5.31 $Y=2.59 $X2=4.205
+ $Y2=1.85
cc_547 N_CK_c_687_n N_A_217_817#_c_916_n 0.00742068f $X=3.705 $Y=1.85 $X2=4.205
+ $Y2=1.85
cc_548 N_CK_c_688_n N_A_217_817#_c_916_n 7.18106e-19 $X=3.705 $Y=1.85 $X2=4.205
+ $Y2=1.85
cc_549 N_CK_c_693_n N_A_217_817#_c_916_n 0.00102309f $X=5.31 $Y=2.59 $X2=4.205
+ $Y2=1.85
cc_550 N_CK_c_702_n N_A_618_89#_c_1037_n 0.0252931f $X=3.705 $Y=1.685 $X2=3.165
+ $Y2=1.685
cc_551 N_CK_c_687_n N_A_618_89#_c_1040_n 0.00613747f $X=3.705 $Y=1.85 $X2=3.285
+ $Y2=2.225
cc_552 N_CK_c_687_n N_A_618_89#_c_1041_n 0.00630484f $X=3.705 $Y=1.85 $X2=3.69
+ $Y2=2.3
cc_553 N_CK_c_688_n N_A_618_89#_c_1041_n 0.0183603f $X=3.705 $Y=1.85 $X2=3.69
+ $Y2=2.3
cc_554 N_CK_c_693_n N_A_618_89#_c_1041_n 0.00613485f $X=5.31 $Y=2.59 $X2=3.69
+ $Y2=2.3
cc_555 N_CK_c_686_n N_A_618_89#_c_1042_n 0.00878348f $X=3.62 $Y=2.59 $X2=3.36
+ $Y2=2.3
cc_556 N_CK_c_694_n N_A_618_89#_c_1042_n 0.00137501f $X=3.37 $Y=2.59 $X2=3.36
+ $Y2=2.3
cc_557 N_CK_c_697_n N_A_618_89#_c_1042_n 0.00109468f $X=3.225 $Y=2.59 $X2=3.36
+ $Y2=2.3
cc_558 N_CK_c_701_n N_A_618_89#_c_1042_n 0.00904036f $X=3.225 $Y=2.765 $X2=3.36
+ $Y2=2.3
cc_559 N_CK_M1023_g N_A_618_89#_M1030_g 0.0612221f $X=3.165 $Y=4.585 $X2=3.765
+ $Y2=4.585
cc_560 N_CK_c_686_n N_A_618_89#_M1030_g 0.0081071f $X=3.62 $Y=2.59 $X2=3.765
+ $Y2=4.585
cc_561 N_CK_c_687_n N_A_618_89#_M1030_g 0.00478024f $X=3.705 $Y=1.85 $X2=3.765
+ $Y2=4.585
cc_562 N_CK_c_693_n N_A_618_89#_M1030_g 0.00938974f $X=5.31 $Y=2.59 $X2=3.765
+ $Y2=4.585
cc_563 N_CK_c_694_n N_A_618_89#_M1030_g 4.2e-19 $X=3.37 $Y=2.59 $X2=3.765
+ $Y2=4.585
cc_564 N_CK_c_697_n N_A_618_89#_M1030_g 0.00184124f $X=3.225 $Y=2.59 $X2=3.765
+ $Y2=4.585
cc_565 N_CK_c_701_n N_A_618_89#_M1030_g 0.0128384f $X=3.225 $Y=2.765 $X2=3.765
+ $Y2=4.585
cc_566 N_CK_c_693_n N_A_618_89#_c_1044_n 0.00607908f $X=5.31 $Y=2.59 $X2=4.84
+ $Y2=2.3
cc_567 N_CK_M1011_g N_A_618_89#_M1010_g 0.0612221f $X=5.515 $Y=4.585 $X2=4.915
+ $Y2=4.585
cc_568 N_CK_c_689_n N_A_618_89#_M1010_g 0.00399495f $X=4.975 $Y=1.85 $X2=4.915
+ $Y2=4.585
cc_569 N_CK_c_692_n N_A_618_89#_M1010_g 0.00654233f $X=5.06 $Y=2.59 $X2=4.915
+ $Y2=4.585
cc_570 N_CK_c_693_n N_A_618_89#_M1010_g 0.00497421f $X=5.31 $Y=2.59 $X2=4.915
+ $Y2=4.585
cc_571 N_CK_c_696_n N_A_618_89#_M1010_g 4.2e-19 $X=5.6 $Y=2.59 $X2=4.915
+ $Y2=4.585
cc_572 N_CK_c_698_n N_A_618_89#_M1010_g 0.00128351f $X=5.455 $Y=2.59 $X2=4.915
+ $Y2=4.585
cc_573 N_CK_c_708_n N_A_618_89#_M1010_g 0.0118393f $X=5.455 $Y=2.765 $X2=4.915
+ $Y2=4.585
cc_574 N_CK_c_689_n N_A_618_89#_c_1046_n 0.00909647f $X=4.975 $Y=1.85 $X2=5.32
+ $Y2=2.3
cc_575 N_CK_c_691_n N_A_618_89#_c_1046_n 0.00924811f $X=5.37 $Y=2.59 $X2=5.32
+ $Y2=2.3
cc_576 N_CK_c_693_n N_A_618_89#_c_1046_n 0.00613485f $X=5.31 $Y=2.59 $X2=5.32
+ $Y2=2.3
cc_577 N_CK_c_696_n N_A_618_89#_c_1046_n 0.00137501f $X=5.6 $Y=2.59 $X2=5.32
+ $Y2=2.3
cc_578 N_CK_c_698_n N_A_618_89#_c_1046_n 0.00102633f $X=5.455 $Y=2.59 $X2=5.32
+ $Y2=2.3
cc_579 N_CK_c_708_n N_A_618_89#_c_1046_n 0.00904036f $X=5.455 $Y=2.765 $X2=5.32
+ $Y2=2.3
cc_580 N_CK_c_689_n N_A_618_89#_c_1047_n 0.00649764f $X=4.975 $Y=1.85 $X2=5.395
+ $Y2=2.225
cc_581 N_CK_c_688_n N_A_618_89#_c_1048_n 0.0216263f $X=3.705 $Y=1.85 $X2=3.285
+ $Y2=1.76
cc_582 N_CK_c_697_n N_A_618_89#_c_1048_n 2.45465e-19 $X=3.225 $Y=2.59 $X2=3.285
+ $Y2=1.76
cc_583 N_CK_c_687_n N_A_618_89#_c_1049_n 0.00568091f $X=3.705 $Y=1.85 $X2=3.765
+ $Y2=2.3
cc_584 N_CK_c_689_n N_A_618_89#_c_1050_n 0.00436024f $X=4.975 $Y=1.85 $X2=4.915
+ $Y2=2.3
cc_585 N_CK_c_690_n N_A_618_89#_c_1050_n 0.0183603f $X=4.975 $Y=1.85 $X2=4.915
+ $Y2=2.3
cc_586 N_CK_c_679_n N_A_618_89#_c_1051_n 0.00592387f $X=6.36 $Y=2.6 $X2=6.435
+ $Y2=1.85
cc_587 N_CK_c_685_n N_A_618_89#_c_1051_n 0.00762848f $X=6.332 $Y=1.835 $X2=6.435
+ $Y2=1.85
cc_588 N_CK_c_689_n N_A_618_89#_c_1051_n 0.00853323f $X=4.975 $Y=1.85 $X2=6.435
+ $Y2=1.85
cc_589 N_CK_c_690_n N_A_618_89#_c_1051_n 8.05876e-19 $X=4.975 $Y=1.85 $X2=6.435
+ $Y2=1.85
cc_590 N_CK_c_691_n N_A_618_89#_c_1051_n 0.00132011f $X=5.37 $Y=2.59 $X2=6.435
+ $Y2=1.85
cc_591 N_CK_c_693_n N_A_618_89#_c_1051_n 3.12599e-19 $X=5.31 $Y=2.59 $X2=6.435
+ $Y2=1.85
cc_592 N_CK_c_695_n N_A_618_89#_c_1051_n 0.00341454f $X=6.305 $Y=2.59 $X2=6.435
+ $Y2=1.85
cc_593 N_CK_c_696_n N_A_618_89#_c_1051_n 0.00221563f $X=5.6 $Y=2.59 $X2=6.435
+ $Y2=1.85
cc_594 N_CK_c_698_n N_A_618_89#_c_1051_n 0.00261697f $X=5.455 $Y=2.59 $X2=6.435
+ $Y2=1.85
cc_595 N_CK_c_700_n N_A_618_89#_c_1051_n 8.24249e-19 $X=6.45 $Y=2.59 $X2=6.435
+ $Y2=1.85
cc_596 N_CK_c_708_n N_A_618_89#_c_1051_n 5.56676e-19 $X=5.455 $Y=2.765 $X2=6.435
+ $Y2=1.85
cc_597 N_CK_c_689_n N_A_618_89#_c_1053_n 0.00131283f $X=4.975 $Y=1.85 $X2=5.455
+ $Y2=1.85
cc_598 N_CK_c_690_n N_A_618_89#_c_1053_n 0.0220721f $X=4.975 $Y=1.85 $X2=5.455
+ $Y2=1.85
cc_599 N_CK_c_696_n N_A_618_89#_c_1053_n 8.78837e-19 $X=5.6 $Y=2.59 $X2=5.455
+ $Y2=1.85
cc_600 N_CK_c_698_n N_A_618_89#_c_1053_n 5.27321e-19 $X=5.455 $Y=2.59 $X2=5.455
+ $Y2=1.85
cc_601 N_CK_c_708_n N_A_618_89#_c_1053_n 0.00227671f $X=5.455 $Y=2.765 $X2=5.455
+ $Y2=1.85
cc_602 N_CK_c_680_n N_A_618_89#_c_1054_n 0.0102351f $X=6.332 $Y=1.685 $X2=6.52
+ $Y2=0.825
cc_603 N_CK_c_685_n N_A_618_89#_c_1054_n 0.00236772f $X=6.332 $Y=1.835 $X2=6.52
+ $Y2=0.825
cc_604 N_CK_c_679_n N_A_618_89#_c_1059_n 0.00603032f $X=6.36 $Y=2.6 $X2=6.52
+ $Y2=2.105
cc_605 N_CK_c_678_n N_A_618_89#_c_1060_n 0.00333903f $X=6.305 $Y=2.93 $X2=6.795
+ $Y2=3.1
cc_606 N_CK_M1031_g N_A_618_89#_c_1060_n 0.00495264f $X=6.305 $Y=4.585 $X2=6.795
+ $Y2=3.1
cc_607 N_CK_c_679_n N_A_618_89#_c_1060_n 0.0075286f $X=6.36 $Y=2.6 $X2=6.795
+ $Y2=3.1
cc_608 CK N_A_618_89#_c_1060_n 0.00852929f $X=6.45 $Y=2.59 $X2=6.795 $Y2=3.1
cc_609 N_CK_c_700_n N_A_618_89#_c_1060_n 0.0289277f $X=6.45 $Y=2.59 $X2=6.795
+ $Y2=3.1
cc_610 N_CK_c_679_n N_A_618_89#_c_1061_n 0.00126138f $X=6.36 $Y=2.6 $X2=6.52
+ $Y2=1.85
cc_611 N_CK_c_685_n N_A_618_89#_c_1061_n 8.88113e-19 $X=6.332 $Y=1.835 $X2=6.52
+ $Y2=1.85
cc_612 N_CK_c_678_n N_A_618_89#_c_1062_n 0.001573f $X=6.305 $Y=2.93 $X2=6.795
+ $Y2=2.19
cc_613 N_CK_c_679_n N_A_618_89#_c_1062_n 0.00437187f $X=6.36 $Y=2.6 $X2=6.795
+ $Y2=2.19
cc_614 CK N_A_618_89#_c_1062_n 8.7939e-19 $X=6.45 $Y=2.59 $X2=6.795 $Y2=2.19
cc_615 N_CK_c_700_n N_A_618_89#_c_1062_n 0.00528683f $X=6.45 $Y=2.59 $X2=6.795
+ $Y2=2.19
cc_616 N_CK_c_678_n N_A_618_89#_c_1076_n 0.00260941f $X=6.305 $Y=2.93 $X2=6.795
+ $Y2=3.185
cc_617 CK N_A_618_89#_c_1076_n 0.00259785f $X=6.45 $Y=2.59 $X2=6.795 $Y2=3.185
cc_618 N_CK_c_700_n N_A_618_89#_c_1076_n 0.00706443f $X=6.45 $Y=2.59 $X2=6.795
+ $Y2=3.185
cc_619 N_CK_c_705_n N_A_618_89#_c_1063_n 0.0268981f $X=4.975 $Y=1.685 $X2=5.455
+ $Y2=1.685
cc_620 N_CK_c_679_n N_A_1160_89#_M1018_g 0.00697006f $X=6.36 $Y=2.6 $X2=5.875
+ $Y2=1.075
cc_621 N_CK_c_680_n N_A_1160_89#_M1018_g 0.0287519f $X=6.332 $Y=1.685 $X2=5.875
+ $Y2=1.075
cc_622 N_CK_c_678_n N_A_1160_89#_M1009_g 0.0287701f $X=6.305 $Y=2.93 $X2=5.875
+ $Y2=4.585
cc_623 N_CK_c_679_n N_A_1160_89#_M1009_g 0.0175925f $X=6.36 $Y=2.6 $X2=5.875
+ $Y2=4.585
cc_624 N_CK_c_695_n N_A_1160_89#_M1009_g 0.0114893f $X=6.305 $Y=2.59 $X2=5.875
+ $Y2=4.585
cc_625 N_CK_c_696_n N_A_1160_89#_M1009_g 0.00113587f $X=5.6 $Y=2.59 $X2=5.875
+ $Y2=4.585
cc_626 N_CK_c_698_n N_A_1160_89#_M1009_g 0.00453616f $X=5.455 $Y=2.59 $X2=5.875
+ $Y2=4.585
cc_627 CK N_A_1160_89#_M1009_g 3.05655e-19 $X=6.45 $Y=2.59 $X2=5.875 $Y2=4.585
cc_628 N_CK_c_700_n N_A_1160_89#_M1009_g 0.0026346f $X=6.45 $Y=2.59 $X2=5.875
+ $Y2=4.585
cc_629 N_CK_c_708_n N_A_1160_89#_M1009_g 0.214863f $X=5.455 $Y=2.765 $X2=5.875
+ $Y2=4.585
cc_630 N_CK_c_678_n N_A_1160_89#_c_1242_n 2.34467e-19 $X=6.305 $Y=2.93 $X2=8.375
+ $Y2=2.19
cc_631 N_CK_c_679_n N_A_1160_89#_c_1242_n 0.0033485f $X=6.36 $Y=2.6 $X2=8.375
+ $Y2=2.19
cc_632 N_CK_c_695_n N_A_1160_89#_c_1242_n 0.0179446f $X=6.305 $Y=2.59 $X2=8.375
+ $Y2=2.19
cc_633 CK N_A_1160_89#_c_1242_n 0.0248956f $X=6.45 $Y=2.59 $X2=8.375 $Y2=2.19
cc_634 N_CK_c_700_n N_A_1160_89#_c_1242_n 8.38639e-19 $X=6.45 $Y=2.59 $X2=8.375
+ $Y2=2.19
cc_635 N_CK_c_679_n N_A_1160_89#_c_1243_n 8.66236e-19 $X=6.36 $Y=2.6 $X2=6.08
+ $Y2=2.19
cc_636 N_CK_c_695_n N_A_1160_89#_c_1243_n 0.0247156f $X=6.305 $Y=2.59 $X2=6.08
+ $Y2=2.19
cc_637 N_CK_c_679_n N_A_1160_89#_c_1244_n 8.95026e-19 $X=6.36 $Y=2.6 $X2=5.935
+ $Y2=2.19
cc_638 N_CK_c_695_n N_A_1160_89#_c_1244_n 0.00488871f $X=6.305 $Y=2.59 $X2=5.935
+ $Y2=2.19
cc_639 N_CK_c_679_n N_A_1160_89#_c_1247_n 0.0213817f $X=6.36 $Y=2.6 $X2=5.935
+ $Y2=2.19
cc_640 N_CK_c_695_n N_A_1160_89#_c_1247_n 0.00185875f $X=6.305 $Y=2.59 $X2=5.935
+ $Y2=2.19
cc_641 N_CK_c_685_n N_A_998_115#_c_1390_n 0.00562911f $X=6.332 $Y=1.835
+ $X2=7.255 $Y2=2.015
cc_642 N_CK_c_678_n N_A_998_115#_M1024_g 0.0044653f $X=6.305 $Y=2.93 $X2=7.255
+ $Y2=5.085
cc_643 N_CK_c_689_n N_A_998_115#_c_1416_n 0.0103267f $X=4.975 $Y=1.85 $X2=5.045
+ $Y2=1.43
cc_644 N_CK_c_690_n N_A_998_115#_c_1416_n 0.00227744f $X=4.975 $Y=1.85 $X2=5.045
+ $Y2=1.43
cc_645 N_CK_c_705_n N_A_998_115#_c_1416_n 0.0149609f $X=4.975 $Y=1.685 $X2=5.045
+ $Y2=1.43
cc_646 N_CK_c_691_n N_A_998_115#_c_1429_n 0.00843004f $X=5.37 $Y=2.59 $X2=5.045
+ $Y2=3.185
cc_647 N_CK_c_692_n N_A_998_115#_c_1429_n 0.00323798f $X=5.06 $Y=2.59 $X2=5.045
+ $Y2=3.185
cc_648 N_CK_c_693_n N_A_998_115#_c_1429_n 0.012754f $X=5.31 $Y=2.59 $X2=5.045
+ $Y2=3.185
cc_649 N_CK_c_696_n N_A_998_115#_c_1429_n 0.00146098f $X=5.6 $Y=2.59 $X2=5.045
+ $Y2=3.185
cc_650 N_CK_c_698_n N_A_998_115#_c_1429_n 0.00103871f $X=5.455 $Y=2.59 $X2=5.045
+ $Y2=3.185
cc_651 N_CK_c_708_n N_A_998_115#_c_1429_n 0.00150627f $X=5.455 $Y=2.765
+ $X2=5.045 $Y2=3.185
cc_652 N_CK_c_679_n N_A_998_115#_c_1396_n 0.00128484f $X=6.36 $Y=2.6 $X2=6.985
+ $Y2=1.85
cc_653 N_CK_c_685_n N_A_998_115#_c_1396_n 0.00179204f $X=6.332 $Y=1.835
+ $X2=6.985 $Y2=1.85
cc_654 N_CK_c_689_n N_A_998_115#_c_1396_n 0.0127028f $X=4.975 $Y=1.85 $X2=6.985
+ $Y2=1.85
cc_655 N_CK_c_690_n N_A_998_115#_c_1396_n 0.00362401f $X=4.975 $Y=1.85 $X2=6.985
+ $Y2=1.85
cc_656 N_CK_c_691_n N_A_998_115#_c_1396_n 0.00451177f $X=5.37 $Y=2.59 $X2=6.985
+ $Y2=1.85
cc_657 N_CK_c_696_n N_A_998_115#_c_1396_n 0.0144351f $X=5.6 $Y=2.59 $X2=6.985
+ $Y2=1.85
cc_658 N_CK_c_698_n N_A_998_115#_c_1396_n 6.39375e-19 $X=5.455 $Y=2.59 $X2=6.985
+ $Y2=1.85
cc_659 N_CK_c_689_n N_A_998_115#_c_1398_n 0.00180575f $X=4.975 $Y=1.85 $X2=4.78
+ $Y2=1.85
cc_660 N_CK_c_690_n N_A_998_115#_c_1398_n 9.79344e-19 $X=4.975 $Y=1.85 $X2=4.78
+ $Y2=1.85
cc_661 N_CK_c_693_n N_A_998_115#_c_1398_n 0.0128239f $X=5.31 $Y=2.59 $X2=4.78
+ $Y2=1.85
cc_662 N_CK_c_689_n N_A_998_115#_c_1399_n 0.057541f $X=4.975 $Y=1.85 $X2=4.635
+ $Y2=1.85
cc_663 N_CK_c_692_n N_A_998_115#_c_1399_n 0.0116326f $X=5.06 $Y=2.59 $X2=4.635
+ $Y2=1.85
cc_664 N_CK_c_693_n N_A_998_115#_c_1399_n 0.020361f $X=5.31 $Y=2.59 $X2=4.635
+ $Y2=1.85
cc_665 N_CK_c_696_n N_A_998_115#_c_1399_n 6.61118e-19 $X=5.6 $Y=2.59 $X2=4.635
+ $Y2=1.85
cc_666 N_CK_c_698_n N_A_998_115#_c_1399_n 0.00613815f $X=5.455 $Y=2.59 $X2=4.635
+ $Y2=1.85
cc_667 N_CK_c_705_n N_A_998_115#_c_1399_n 0.00554221f $X=4.975 $Y=1.685
+ $X2=4.635 $Y2=1.85
cc_668 N_CK_c_685_n N_A_998_115#_c_1401_n 2.33995e-19 $X=6.332 $Y=1.835 $X2=7.13
+ $Y2=1.85
cc_669 N_A_217_817#_c_914_n N_A_618_89#_c_1040_n 0.00253253f $X=4.06 $Y=1.85
+ $X2=3.285 $Y2=2.225
cc_670 N_A_217_817#_c_914_n N_A_618_89#_c_1041_n 0.00296105f $X=4.06 $Y=1.85
+ $X2=3.69 $Y2=2.3
cc_671 N_A_217_817#_c_906_n N_A_618_89#_M1030_g 0.215335f $X=4.2 $Y=2.765
+ $X2=3.765 $Y2=4.585
cc_672 N_A_217_817#_c_913_n N_A_618_89#_M1030_g 0.00486364f $X=4.295 $Y=2.765
+ $X2=3.765 $Y2=4.585
cc_673 N_A_217_817#_c_905_n N_A_618_89#_c_1044_n 0.0342351f $X=4.2 $Y=1.85
+ $X2=4.84 $Y2=2.3
cc_674 N_A_217_817#_c_906_n N_A_618_89#_c_1044_n 0.0307748f $X=4.2 $Y=2.765
+ $X2=4.84 $Y2=2.3
cc_675 N_A_217_817#_c_913_n N_A_618_89#_c_1044_n 0.0113171f $X=4.295 $Y=2.765
+ $X2=4.84 $Y2=2.3
cc_676 N_A_217_817#_c_914_n N_A_618_89#_c_1044_n 0.00486036f $X=4.06 $Y=1.85
+ $X2=4.84 $Y2=2.3
cc_677 N_A_217_817#_c_960_n N_A_618_89#_c_1044_n 4.12801e-19 $X=4.205 $Y=1.85
+ $X2=4.84 $Y2=2.3
cc_678 N_A_217_817#_c_916_n N_A_618_89#_c_1044_n 8.69982e-19 $X=4.205 $Y=1.85
+ $X2=4.84 $Y2=2.3
cc_679 N_A_217_817#_c_909_n N_A_618_89#_M1010_g 0.211921f $X=4.48 $Y=2.765
+ $X2=4.915 $Y2=4.585
cc_680 N_A_217_817#_M1022_g N_A_998_115#_c_1417_n 0.00136315f $X=4.125 $Y=1.075
+ $X2=4.72 $Y2=1.43
cc_681 N_A_217_817#_M1019_g N_A_998_115#_c_1417_n 0.0099627f $X=4.555 $Y=1.075
+ $X2=4.72 $Y2=1.43
cc_682 N_A_217_817#_M1028_g N_A_998_115#_c_1454_n 9.13132e-19 $X=4.125 $Y=4.585
+ $X2=4.72 $Y2=3.185
cc_683 N_A_217_817#_M1006_g N_A_998_115#_c_1454_n 0.0096885f $X=4.555 $Y=4.585
+ $X2=4.72 $Y2=3.185
cc_684 N_A_217_817#_c_907_n N_A_998_115#_c_1398_n 0.00229064f $X=4.48 $Y=1.85
+ $X2=4.78 $Y2=1.85
cc_685 N_A_217_817#_c_960_n N_A_998_115#_c_1398_n 0.0241863f $X=4.205 $Y=1.85
+ $X2=4.78 $Y2=1.85
cc_686 N_A_217_817#_c_916_n N_A_998_115#_c_1398_n 0.0012094f $X=4.205 $Y=1.85
+ $X2=4.78 $Y2=1.85
cc_687 N_A_217_817#_M1022_g N_A_998_115#_c_1399_n 0.001069f $X=4.125 $Y=1.075
+ $X2=4.635 $Y2=1.85
cc_688 N_A_217_817#_M1028_g N_A_998_115#_c_1399_n 9.36754e-19 $X=4.125 $Y=4.585
+ $X2=4.635 $Y2=1.85
cc_689 N_A_217_817#_M1019_g N_A_998_115#_c_1399_n 0.00502021f $X=4.555 $Y=1.075
+ $X2=4.635 $Y2=1.85
cc_690 N_A_217_817#_M1006_g N_A_998_115#_c_1399_n 0.00479454f $X=4.555 $Y=4.585
+ $X2=4.635 $Y2=1.85
cc_691 N_A_217_817#_c_907_n N_A_998_115#_c_1399_n 0.0061959f $X=4.48 $Y=1.85
+ $X2=4.635 $Y2=1.85
cc_692 N_A_217_817#_c_909_n N_A_998_115#_c_1399_n 0.00738718f $X=4.48 $Y=2.765
+ $X2=4.635 $Y2=1.85
cc_693 N_A_217_817#_c_913_n N_A_998_115#_c_1399_n 0.0702347f $X=4.295 $Y=2.765
+ $X2=4.635 $Y2=1.85
cc_694 N_A_217_817#_c_960_n N_A_998_115#_c_1399_n 4.18442e-19 $X=4.205 $Y=1.85
+ $X2=4.635 $Y2=1.85
cc_695 N_A_217_817#_c_916_n N_A_998_115#_c_1399_n 0.0157315f $X=4.205 $Y=1.85
+ $X2=4.635 $Y2=1.85
cc_696 N_A_618_89#_c_1047_n N_A_1160_89#_M1018_g 0.0073696f $X=5.395 $Y=2.225
+ $X2=5.875 $Y2=1.075
cc_697 N_A_618_89#_c_1051_n N_A_1160_89#_M1018_g 0.0107575f $X=6.435 $Y=1.85
+ $X2=5.875 $Y2=1.075
cc_698 N_A_618_89#_c_1063_n N_A_1160_89#_M1018_g 0.0974852f $X=5.455 $Y=1.685
+ $X2=5.875 $Y2=1.075
cc_699 N_A_618_89#_c_1072_n N_A_1160_89#_c_1260_n 0.0951397f $X=6.52 $Y=3.455
+ $X2=7.04 $Y2=4.475
cc_700 N_A_618_89#_c_1072_n N_A_1160_89#_c_1264_n 0.00835159f $X=6.52 $Y=3.455
+ $X2=7.125 $Y2=3.78
cc_701 N_A_618_89#_c_1060_n N_A_1160_89#_c_1240_n 0.0293498f $X=6.795 $Y=3.1
+ $X2=7.47 $Y2=3.695
cc_702 N_A_618_89#_c_1076_n N_A_1160_89#_c_1240_n 0.00644034f $X=6.795 $Y=3.185
+ $X2=7.47 $Y2=3.695
cc_703 N_A_618_89#_c_1062_n N_A_1160_89#_c_1241_n 0.00391844f $X=6.795 $Y=2.19
+ $X2=7.47 $Y2=2.19
cc_704 N_A_618_89#_c_1051_n N_A_1160_89#_c_1242_n 0.00314603f $X=6.435 $Y=1.85
+ $X2=8.375 $Y2=2.19
cc_705 N_A_618_89#_c_1059_n N_A_1160_89#_c_1242_n 6.94255e-19 $X=6.52 $Y=2.105
+ $X2=8.375 $Y2=2.19
cc_706 N_A_618_89#_c_1060_n N_A_1160_89#_c_1242_n 0.00492501f $X=6.795 $Y=3.1
+ $X2=8.375 $Y2=2.19
cc_707 N_A_618_89#_c_1062_n N_A_1160_89#_c_1242_n 0.0228595f $X=6.795 $Y=2.19
+ $X2=8.375 $Y2=2.19
cc_708 N_A_618_89#_c_1047_n N_A_1160_89#_c_1243_n 9.14174e-19 $X=5.395 $Y=2.225
+ $X2=6.08 $Y2=2.19
cc_709 N_A_618_89#_c_1051_n N_A_1160_89#_c_1243_n 0.0010261f $X=6.435 $Y=1.85
+ $X2=6.08 $Y2=2.19
cc_710 N_A_618_89#_c_1059_n N_A_1160_89#_c_1243_n 0.00122156f $X=6.52 $Y=2.105
+ $X2=6.08 $Y2=2.19
cc_711 N_A_618_89#_c_1047_n N_A_1160_89#_c_1244_n 0.0035305f $X=5.395 $Y=2.225
+ $X2=5.935 $Y2=2.19
cc_712 N_A_618_89#_c_1051_n N_A_1160_89#_c_1244_n 0.0219931f $X=6.435 $Y=1.85
+ $X2=5.935 $Y2=2.19
cc_713 N_A_618_89#_c_1062_n N_A_1160_89#_c_1244_n 0.00559578f $X=6.795 $Y=2.19
+ $X2=5.935 $Y2=2.19
cc_714 N_A_618_89#_c_1046_n N_A_1160_89#_c_1247_n 0.0073696f $X=5.32 $Y=2.3
+ $X2=5.935 $Y2=2.19
cc_715 N_A_618_89#_c_1051_n N_A_1160_89#_c_1247_n 0.00290516f $X=6.435 $Y=1.85
+ $X2=5.935 $Y2=2.19
cc_716 N_A_618_89#_c_1062_n N_A_1160_89#_c_1247_n 2.97404e-19 $X=6.795 $Y=2.19
+ $X2=5.935 $Y2=2.19
cc_717 N_A_618_89#_c_1054_n N_A_998_115#_M1007_g 0.01304f $X=6.52 $Y=0.825
+ $X2=7.255 $Y2=0.945
cc_718 N_A_618_89#_c_1054_n N_A_998_115#_c_1390_n 7.31267e-19 $X=6.52 $Y=0.825
+ $X2=7.255 $Y2=2.015
cc_719 N_A_618_89#_c_1059_n N_A_998_115#_c_1390_n 6.06312e-19 $X=6.52 $Y=2.105
+ $X2=7.255 $Y2=2.015
cc_720 N_A_618_89#_c_1061_n N_A_998_115#_c_1390_n 9.90959e-19 $X=6.52 $Y=1.85
+ $X2=7.255 $Y2=2.015
cc_721 N_A_618_89#_c_1059_n N_A_998_115#_M1024_g 0.00201047f $X=6.52 $Y=2.105
+ $X2=7.255 $Y2=5.085
cc_722 N_A_618_89#_c_1072_n N_A_998_115#_M1024_g 0.0148031f $X=6.52 $Y=3.455
+ $X2=7.255 $Y2=5.085
cc_723 N_A_618_89#_c_1060_n N_A_998_115#_M1024_g 0.0127431f $X=6.795 $Y=3.1
+ $X2=7.255 $Y2=5.085
cc_724 N_A_618_89#_c_1062_n N_A_998_115#_M1024_g 0.00243213f $X=6.795 $Y=2.19
+ $X2=7.255 $Y2=5.085
cc_725 N_A_618_89#_c_1076_n N_A_998_115#_M1024_g 0.00343288f $X=6.795 $Y=3.185
+ $X2=7.255 $Y2=5.085
cc_726 N_A_618_89#_c_1051_n N_A_998_115#_c_1416_n 0.00436807f $X=6.435 $Y=1.85
+ $X2=5.045 $Y2=1.43
cc_727 N_A_618_89#_c_1053_n N_A_998_115#_c_1416_n 0.00174784f $X=5.455 $Y=1.85
+ $X2=5.045 $Y2=1.43
cc_728 N_A_618_89#_c_1063_n N_A_998_115#_c_1416_n 0.00205316f $X=5.455 $Y=1.685
+ $X2=5.045 $Y2=1.43
cc_729 N_A_618_89#_M1010_g N_A_998_115#_c_1429_n 0.0162544f $X=4.915 $Y=4.585
+ $X2=5.045 $Y2=3.185
cc_730 N_A_618_89#_c_1044_n N_A_998_115#_c_1396_n 0.00156696f $X=4.84 $Y=2.3
+ $X2=6.985 $Y2=1.85
cc_731 N_A_618_89#_c_1046_n N_A_998_115#_c_1396_n 0.00244106f $X=5.32 $Y=2.3
+ $X2=6.985 $Y2=1.85
cc_732 N_A_618_89#_c_1050_n N_A_998_115#_c_1396_n 5.19983e-19 $X=4.915 $Y=2.3
+ $X2=6.985 $Y2=1.85
cc_733 N_A_618_89#_c_1051_n N_A_998_115#_c_1396_n 0.0492477f $X=6.435 $Y=1.85
+ $X2=6.985 $Y2=1.85
cc_734 N_A_618_89#_c_1053_n N_A_998_115#_c_1396_n 0.00455939f $X=5.455 $Y=1.85
+ $X2=6.985 $Y2=1.85
cc_735 N_A_618_89#_c_1061_n N_A_998_115#_c_1396_n 0.011616f $X=6.52 $Y=1.85
+ $X2=6.985 $Y2=1.85
cc_736 N_A_618_89#_c_1062_n N_A_998_115#_c_1396_n 0.00227434f $X=6.795 $Y=2.19
+ $X2=6.985 $Y2=1.85
cc_737 N_A_618_89#_c_1044_n N_A_998_115#_c_1398_n 0.00120486f $X=4.84 $Y=2.3
+ $X2=4.78 $Y2=1.85
cc_738 N_A_618_89#_c_1044_n N_A_998_115#_c_1399_n 0.0124213f $X=4.84 $Y=2.3
+ $X2=4.635 $Y2=1.85
cc_739 N_A_618_89#_M1010_g N_A_998_115#_c_1399_n 0.0111407f $X=4.915 $Y=4.585
+ $X2=4.635 $Y2=1.85
cc_740 N_A_618_89#_c_1054_n N_A_998_115#_c_1400_n 7.64938e-19 $X=6.52 $Y=0.825
+ $X2=7.13 $Y2=1.85
cc_741 N_A_618_89#_c_1059_n N_A_998_115#_c_1400_n 7.64938e-19 $X=6.52 $Y=2.105
+ $X2=7.13 $Y2=1.85
cc_742 N_A_618_89#_c_1054_n N_A_998_115#_c_1401_n 0.00237811f $X=6.52 $Y=0.825
+ $X2=7.13 $Y2=1.85
cc_743 N_A_618_89#_c_1059_n N_A_998_115#_c_1401_n 0.00237811f $X=6.52 $Y=2.105
+ $X2=7.13 $Y2=1.85
cc_744 N_A_618_89#_c_1061_n N_A_998_115#_c_1401_n 0.00399834f $X=6.52 $Y=1.85
+ $X2=7.13 $Y2=1.85
cc_745 N_A_1160_89#_c_1237_n N_A_998_115#_M1007_g 0.0136957f $X=7.47 $Y=0.825
+ $X2=7.255 $Y2=0.945
cc_746 N_A_1160_89#_c_1242_n N_A_998_115#_c_1390_n 7.97313e-19 $X=8.375 $Y=2.19
+ $X2=7.255 $Y2=2.015
cc_747 N_A_1160_89#_c_1260_n N_A_998_115#_M1024_g 0.013288f $X=7.04 $Y=4.475
+ $X2=7.255 $Y2=5.085
cc_748 N_A_1160_89#_c_1263_n N_A_998_115#_M1024_g 0.0203145f $X=7.385 $Y=3.78
+ $X2=7.255 $Y2=5.085
cc_749 N_A_1160_89#_c_1240_n N_A_998_115#_M1024_g 0.0199913f $X=7.47 $Y=3.695
+ $X2=7.255 $Y2=5.085
cc_750 N_A_1160_89#_c_1241_n N_A_998_115#_M1024_g 0.00172166f $X=7.47 $Y=2.19
+ $X2=7.255 $Y2=5.085
cc_751 N_A_1160_89#_c_1242_n N_A_998_115#_M1024_g 0.0122381f $X=8.375 $Y=2.19
+ $X2=7.255 $Y2=5.085
cc_752 N_A_1160_89#_M1018_g N_A_998_115#_c_1396_n 0.00231271f $X=5.875 $Y=1.075
+ $X2=6.985 $Y2=1.85
cc_753 N_A_1160_89#_c_1242_n N_A_998_115#_c_1396_n 0.0809321f $X=8.375 $Y=2.19
+ $X2=6.985 $Y2=1.85
cc_754 N_A_1160_89#_c_1243_n N_A_998_115#_c_1396_n 0.0289631f $X=6.08 $Y=2.19
+ $X2=6.985 $Y2=1.85
cc_755 N_A_1160_89#_c_1244_n N_A_998_115#_c_1396_n 0.00166223f $X=5.935 $Y=2.19
+ $X2=6.985 $Y2=1.85
cc_756 N_A_1160_89#_c_1247_n N_A_998_115#_c_1396_n 0.00187603f $X=5.935 $Y=2.19
+ $X2=6.985 $Y2=1.85
cc_757 N_A_1160_89#_c_1237_n N_A_998_115#_c_1400_n 0.00695031f $X=7.47 $Y=0.825
+ $X2=7.13 $Y2=1.85
cc_758 N_A_1160_89#_c_1242_n N_A_998_115#_c_1400_n 0.028322f $X=8.375 $Y=2.19
+ $X2=7.13 $Y2=1.85
cc_759 N_A_1160_89#_c_1237_n N_A_998_115#_c_1401_n 0.0214571f $X=7.47 $Y=0.825
+ $X2=7.13 $Y2=1.85
cc_760 N_A_1160_89#_c_1242_n N_A_998_115#_c_1401_n 0.0046086f $X=8.375 $Y=2.19
+ $X2=7.13 $Y2=1.85
cc_761 N_A_1160_89#_M1012_g N_QN_M1004_g 0.0391431f $X=8.635 $Y=0.945 $X2=9.065
+ $Y2=0.945
cc_762 N_A_1160_89#_c_1246_n N_QN_M1004_g 4.79563e-19 $X=8.52 $Y=2.19 $X2=9.065
+ $Y2=0.945
cc_763 N_A_1160_89#_c_1249_n N_QN_M1004_g 0.0153129f $X=8.522 $Y=2.025 $X2=9.065
+ $Y2=0.945
cc_764 N_A_1160_89#_c_1235_n N_QN_M1002_g 0.0102953f $X=8.61 $Y=2.855 $X2=9.065
+ $Y2=5.085
cc_765 N_A_1160_89#_c_1236_n N_QN_M1002_g 0.0662174f $X=8.61 $Y=3.005 $X2=9.065
+ $Y2=5.085
cc_766 N_A_1160_89#_M1012_g N_QN_c_1521_n 0.0171793f $X=8.635 $Y=0.945 $X2=8.42
+ $Y2=0.825
cc_767 N_A_1160_89#_c_1234_n N_QN_c_1521_n 0.00351772f $X=8.61 $Y=1.8 $X2=8.42
+ $Y2=0.825
cc_768 N_A_1160_89#_c_1234_n N_QN_c_1525_n 0.011031f $X=8.61 $Y=1.8 $X2=8.92
+ $Y2=1.85
cc_769 N_A_1160_89#_c_1245_n N_QN_c_1525_n 0.00387586f $X=8.52 $Y=2.19 $X2=8.92
+ $Y2=1.85
cc_770 N_A_1160_89#_c_1246_n N_QN_c_1525_n 0.0110498f $X=8.52 $Y=2.19 $X2=8.92
+ $Y2=1.85
cc_771 N_A_1160_89#_c_1249_n N_QN_c_1525_n 0.00799433f $X=8.522 $Y=2.025
+ $X2=8.92 $Y2=1.85
cc_772 N_A_1160_89#_c_1242_n N_QN_c_1526_n 0.0010572f $X=8.375 $Y=2.19 $X2=8.505
+ $Y2=1.85
cc_773 N_A_1160_89#_c_1245_n N_QN_c_1526_n 0.00336135f $X=8.52 $Y=2.19 $X2=8.505
+ $Y2=1.85
cc_774 N_A_1160_89#_c_1246_n N_QN_c_1526_n 0.0120703f $X=8.52 $Y=2.19 $X2=8.505
+ $Y2=1.85
cc_775 N_A_1160_89#_c_1248_n N_QN_c_1526_n 0.00308111f $X=8.52 $Y=2.19 $X2=8.505
+ $Y2=1.85
cc_776 N_A_1160_89#_c_1235_n N_QN_c_1527_n 0.016126f $X=8.61 $Y=2.855 $X2=8.92
+ $Y2=2.765
cc_777 N_A_1160_89#_c_1236_n N_QN_c_1527_n 0.00248624f $X=8.61 $Y=3.005 $X2=8.92
+ $Y2=2.765
cc_778 N_A_1160_89#_c_1245_n N_QN_c_1527_n 0.00253233f $X=8.52 $Y=2.19 $X2=8.92
+ $Y2=2.765
cc_779 N_A_1160_89#_c_1246_n N_QN_c_1527_n 0.00426371f $X=8.52 $Y=2.19 $X2=8.92
+ $Y2=2.765
cc_780 N_A_1160_89#_c_1242_n N_QN_c_1528_n 9.40773e-19 $X=8.375 $Y=2.19
+ $X2=8.505 $Y2=2.765
cc_781 N_A_1160_89#_c_1245_n N_QN_c_1528_n 0.00140341f $X=8.52 $Y=2.19 $X2=8.505
+ $Y2=2.765
cc_782 N_A_1160_89#_c_1246_n N_QN_c_1528_n 0.00471962f $X=8.52 $Y=2.19 $X2=8.505
+ $Y2=2.765
cc_783 N_A_1160_89#_c_1248_n N_QN_c_1528_n 0.00265611f $X=8.52 $Y=2.19 $X2=8.505
+ $Y2=2.765
cc_784 N_A_1160_89#_c_1235_n N_QN_c_1529_n 0.00226435f $X=8.61 $Y=2.855
+ $X2=9.005 $Y2=2.395
cc_785 N_A_1160_89#_c_1245_n N_QN_c_1529_n 0.00377439f $X=8.52 $Y=2.19 $X2=9.005
+ $Y2=2.395
cc_786 N_A_1160_89#_c_1246_n N_QN_c_1529_n 0.00987106f $X=8.52 $Y=2.19 $X2=9.005
+ $Y2=2.395
cc_787 N_A_1160_89#_c_1248_n N_QN_c_1529_n 0.00216137f $X=8.52 $Y=2.19 $X2=9.005
+ $Y2=2.395
cc_788 N_A_1160_89#_c_1249_n N_QN_c_1529_n 0.00323473f $X=8.522 $Y=2.025
+ $X2=9.005 $Y2=2.395
cc_789 N_A_1160_89#_c_1245_n N_QN_c_1530_n 4.60229e-19 $X=8.52 $Y=2.19 $X2=9.005
+ $Y2=2.395
cc_790 N_A_1160_89#_c_1246_n N_QN_c_1530_n 3.0115e-19 $X=8.52 $Y=2.19 $X2=9.005
+ $Y2=2.395
cc_791 N_A_1160_89#_c_1248_n N_QN_c_1530_n 0.021196f $X=8.52 $Y=2.19 $X2=9.005
+ $Y2=2.395
cc_792 N_A_1160_89#_M1025_g N_QN_c_1531_n 0.0462756f $X=8.635 $Y=5.085 $X2=8.42
+ $Y2=2.96
cc_793 N_A_1160_89#_c_1235_n N_QN_c_1531_n 0.00567875f $X=8.61 $Y=2.855 $X2=8.42
+ $Y2=2.96
cc_794 N_A_1160_89#_M1025_g QN 0.00233857f $X=8.635 $Y=5.085 $X2=8.425 $Y2=2.96
cc_795 N_A_1160_89#_c_1236_n QN 0.00508004f $X=8.61 $Y=3.005 $X2=8.425 $Y2=2.96
cc_796 N_A_1160_89#_c_1240_n QN 0.00513409f $X=7.47 $Y=3.695 $X2=8.425 $Y2=2.96
cc_797 N_A_1160_89#_c_1245_n QN 0.00842298f $X=8.52 $Y=2.19 $X2=8.425 $Y2=2.96
cc_798 N_A_1160_89#_c_1246_n QN 0.00359685f $X=8.52 $Y=2.19 $X2=8.425 $Y2=2.96
cc_799 N_A_1160_89#_M1025_g Q 0.0011399f $X=8.635 $Y=5.085 $X2=9.275 $Y2=3.33
cc_800 N_A_998_115#_c_1429_n A_926_617# 0.00342591f $X=5.045 $Y=3.185 $X2=4.63
+ $Y2=3.085
cc_801 N_A_998_115#_c_1454_n A_926_617# 0.00144354f $X=4.72 $Y=3.185 $X2=4.63
+ $Y2=3.085
cc_802 N_A_998_115#_c_1416_n A_926_115# 0.00337089f $X=5.045 $Y=1.43 $X2=4.63
+ $Y2=0.575
cc_803 N_A_998_115#_c_1417_n A_926_115# 0.00148865f $X=4.72 $Y=1.43 $X2=4.63
+ $Y2=0.575
cc_804 N_A_998_115#_c_1399_n A_926_115# 9.4749e-19 $X=4.635 $Y=1.85 $X2=4.63
+ $Y2=0.575
cc_805 N_QN_M1004_g N_Q_c_1603_n 0.011148f $X=9.065 $Y=0.945 $X2=9.28 $Y2=0.825
cc_806 N_QN_M1002_g N_Q_c_1607_n 0.0305875f $X=9.065 $Y=5.085 $X2=9.28 $Y2=4.475
cc_807 N_QN_M1004_g N_Q_c_1605_n 0.0383548f $X=9.065 $Y=0.945 $X2=9.395 $Y2=3.16
cc_808 N_QN_c_1525_n N_Q_c_1605_n 0.0111776f $X=8.92 $Y=1.85 $X2=9.395 $Y2=3.16
cc_809 N_QN_c_1527_n N_Q_c_1605_n 0.0111776f $X=8.92 $Y=2.765 $X2=9.395 $Y2=3.16
cc_810 N_QN_c_1529_n N_Q_c_1605_n 0.0438362f $X=9.005 $Y=2.395 $X2=9.395
+ $Y2=3.16
cc_811 N_QN_M1004_g N_Q_c_1606_n 0.00695117f $X=9.065 $Y=0.945 $X2=9.395
+ $Y2=1.515
cc_812 N_QN_M1002_g Q 0.0145232f $X=9.065 $Y=5.085 $X2=9.275 $Y2=3.33
cc_813 N_QN_c_1527_n Q 0.00245821f $X=8.92 $Y=2.765 $X2=9.275 $Y2=3.33
cc_814 N_QN_c_1531_n Q 0.00553023f $X=8.42 $Y=2.96 $X2=9.275 $Y2=3.33
cc_815 N_QN_M1002_g N_Q_c_1612_n 0.00911548f $X=9.065 $Y=5.085 $X2=9.275
+ $Y2=3.33
