* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_12T_hs__dffs_l
** N=27 EP=0 IP=0 FDC=36
M0 17 SN 7 gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=400 $Y=575 $D=19
M1 gnd 4 17 gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=760 $Y=575 $D=19
M2 18 D gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=1780 $Y=575 $D=19
M3 4 8 18 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=2140 $Y=575 $D=19
M4 19 CK 4 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=2740 $Y=575 $D=19
M5 gnd 7 19 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=3100 $Y=575 $D=19
M6 20 7 gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=3530 $Y=575 $D=19
M7 10 CK 20 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=3890 $Y=575 $D=19
M8 21 8 10 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=4490 $Y=575 $D=19
M9 gnd 9 21 gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=4850 $Y=575 $D=19
M10 8 CK gnd gnd nlowvt L=0.15 W=0.55 m=1 r=3.66667 a=0.0825 p=1.4 mult=1 $X=5280 $Y=575 $D=19
M11 22 10 9 gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6230 $Y=575 $D=19
M12 gnd SN 22 gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6590 $Y=575 $D=19
M13 gnd 9 QN gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7610 $Y=575 $D=19
M14 Q QN gnd gnd nlowvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=8040 $Y=575 $D=19
M15 7 SN vdd vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=400 $Y=3025 $D=79
M16 vdd 4 7 vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=830 $Y=3025 $D=79
M17 12 D vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=1780 $Y=2605 $D=79
M18 4 CK 12 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=2140 $Y=2605 $D=79
M19 13 8 4 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=2740 $Y=2605 $D=79
M20 vdd 7 13 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=3100 $Y=2605 $D=79
M21 14 7 vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=3530 $Y=2605 $D=79
M22 10 8 14 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=3890 $Y=2605 $D=79
M23 15 CK 10 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=4490 $Y=2605 $D=79
M24 vdd 9 15 vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=4850 $Y=2605 $D=79
M25 8 CK vdd vdd pshort L=0.15 W=1.26 m=1 r=8.4 a=0.189 p=2.82 mult=1 $X=5280 $Y=2605 $D=79
M26 9 10 vdd vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=6230 $Y=3025 $D=79
M27 vdd SN 9 vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=6660 $Y=3025 $D=79
M28 vdd 9 QN vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=7610 $Y=3025 $D=79
M29 Q QN vdd vdd pshort L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=8040 $Y=3025 $D=79
X30 gnd vdd Dpar a=18.0409 p=21.64 m=1 $[nwdiode] $X=-55 $Y=2815 $D=185
X31 23 SN Probe probetype=1 $[SN] $X=318 $Y=1533 $D=289
X32 24 D Probe probetype=1 $[D] $X=1913 $Y=1738 $D=289
X33 25 CK Probe probetype=1 $[CK] $X=5498 $Y=2108 $D=289
X34 26 QN Probe probetype=1 $[QN] $X=7473 $Y=2478 $D=289
X35 27 Q Probe probetype=1 $[Q] $X=8323 $Y=2848 $D=289
.ENDS
***************************************
