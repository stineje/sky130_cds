* File: sky130_osu_sc_15T_hs__or2_4.pxi.spice
* Created: Fri Nov 12 14:32:48 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__OR2_4%GND N_GND_M1007_s N_GND_M1002_d N_GND_M1009_s
+ N_GND_M1011_s N_GND_M1007_b N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p
+ N_GND_c_24_p N_GND_c_32_p N_GND_c_38_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_15T_HS__OR2_4%GND
x_PM_SKY130_OSU_SC_15T_HS__OR2_4%VDD N_VDD_M1005_d N_VDD_M1001_d N_VDD_M1006_d
+ N_VDD_M1008_b N_VDD_c_75_p N_VDD_c_81_p N_VDD_c_88_p N_VDD_c_94_p
+ N_VDD_c_100_p N_VDD_c_105_p VDD N_VDD_c_76_p
+ PM_SKY130_OSU_SC_15T_HS__OR2_4%VDD
x_PM_SKY130_OSU_SC_15T_HS__OR2_4%B N_B_M1007_g N_B_M1008_g N_B_c_126_n
+ N_B_c_127_n B PM_SKY130_OSU_SC_15T_HS__OR2_4%B
x_PM_SKY130_OSU_SC_15T_HS__OR2_4%A N_A_M1002_g N_A_M1005_g N_A_c_154_n
+ N_A_c_155_n A PM_SKY130_OSU_SC_15T_HS__OR2_4%A
x_PM_SKY130_OSU_SC_15T_HS__OR2_4%A_27_565# N_A_27_565#_M1007_d
+ N_A_27_565#_M1008_s N_A_27_565#_M1004_g N_A_27_565#_c_228_n
+ N_A_27_565#_M1000_g N_A_27_565#_c_197_n N_A_27_565#_c_198_n
+ N_A_27_565#_M1009_g N_A_27_565#_c_233_n N_A_27_565#_M1001_g
+ N_A_27_565#_c_203_n N_A_27_565#_c_205_n N_A_27_565#_c_206_n
+ N_A_27_565#_M1010_g N_A_27_565#_c_240_n N_A_27_565#_M1003_g
+ N_A_27_565#_c_211_n N_A_27_565#_c_212_n N_A_27_565#_M1011_g
+ N_A_27_565#_c_245_n N_A_27_565#_M1006_g N_A_27_565#_c_217_n
+ N_A_27_565#_c_218_n N_A_27_565#_c_219_n N_A_27_565#_c_220_n
+ N_A_27_565#_c_252_n N_A_27_565#_c_256_n N_A_27_565#_c_258_n
+ N_A_27_565#_c_221_n N_A_27_565#_c_222_n N_A_27_565#_c_225_n
+ N_A_27_565#_c_227_n PM_SKY130_OSU_SC_15T_HS__OR2_4%A_27_565#
x_PM_SKY130_OSU_SC_15T_HS__OR2_4%Y N_Y_M1004_d N_Y_M1010_d N_Y_M1000_s
+ N_Y_M1003_s N_Y_c_331_n N_Y_c_335_n N_Y_c_336_n N_Y_c_340_n N_Y_c_341_n
+ N_Y_c_344_n Y N_Y_c_346_n N_Y_c_349_n N_Y_c_350_n N_Y_c_353_n
+ PM_SKY130_OSU_SC_15T_HS__OR2_4%Y
cc_1 N_GND_M1007_b N_B_M1007_g 0.0919998f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_B_M1007_g 0.00866533f $X=0.26 $Y=0.865 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_B_M1007_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.895
cc_4 N_GND_c_4_p N_B_M1007_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=0.895
cc_5 N_GND_M1007_b N_B_M1008_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_6 N_GND_M1007_b N_B_c_126_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.415
cc_7 N_GND_M1007_b N_B_c_127_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.415
cc_8 N_GND_M1007_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.7
cc_9 N_GND_M1007_b N_A_M1002_g 0.0494465f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.895
cc_10 N_GND_c_3_p N_A_M1002_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.895
cc_11 N_GND_c_11_p N_A_M1002_g 0.00388248f $X=1.12 $Y=0.865 $X2=0.905 $Y2=0.895
cc_12 N_GND_c_4_p N_A_M1002_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.905 $Y2=0.895
cc_13 N_GND_M1007_b N_A_M1005_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_14 N_GND_M1007_b N_A_c_154_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.125
cc_15 N_GND_M1007_b N_A_c_155_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.125
cc_16 N_GND_M1007_b N_A_27_565#_M1004_g 0.0255964f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.895
cc_17 N_GND_c_11_p N_A_27_565#_M1004_g 0.00388248f $X=1.12 $Y=0.865 $X2=1.335
+ $Y2=0.895
cc_18 N_GND_c_18_p N_A_27_565#_M1004_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.895
cc_19 N_GND_c_4_p N_A_27_565#_M1004_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.335
+ $Y2=0.895
cc_20 N_GND_M1007_b N_A_27_565#_c_197_n 0.0466273f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.55
cc_21 N_GND_M1007_b N_A_27_565#_c_198_n 0.00954592f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.625
cc_22 N_GND_M1007_b N_A_27_565#_M1009_g 0.0245289f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.895
cc_23 N_GND_c_18_p N_A_27_565#_M1009_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.895
cc_24 N_GND_c_24_p N_A_27_565#_M1009_g 0.00390533f $X=1.98 $Y=0.865 $X2=1.765
+ $Y2=0.895
cc_25 N_GND_c_4_p N_A_27_565#_M1009_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.765
+ $Y2=0.895
cc_26 N_GND_M1007_b N_A_27_565#_c_203_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_27 N_GND_c_24_p N_A_27_565#_c_203_n 0.00256938f $X=1.98 $Y=0.865 $X2=2.12
+ $Y2=1.585
cc_28 N_GND_M1007_b N_A_27_565#_c_205_n 0.0439685f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.585
cc_29 N_GND_M1007_b N_A_27_565#_c_206_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.625
cc_30 N_GND_M1007_b N_A_27_565#_M1010_g 0.0245289f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.895
cc_31 N_GND_c_24_p N_A_27_565#_M1010_g 0.00390533f $X=1.98 $Y=0.865 $X2=2.195
+ $Y2=0.895
cc_32 N_GND_c_32_p N_A_27_565#_M1010_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.895
cc_33 N_GND_c_4_p N_A_27_565#_M1010_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.195
+ $Y2=0.895
cc_34 N_GND_M1007_b N_A_27_565#_c_211_n 0.0369419f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.585
cc_35 N_GND_M1007_b N_A_27_565#_c_212_n 0.0268552f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.625
cc_36 N_GND_M1007_b N_A_27_565#_M1011_g 0.0341369f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.895
cc_37 N_GND_c_32_p N_A_27_565#_M1011_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.895
cc_38 N_GND_c_38_p N_A_27_565#_M1011_g 0.00866533f $X=2.84 $Y=0.865 $X2=2.625
+ $Y2=0.895
cc_39 N_GND_c_4_p N_A_27_565#_M1011_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.625
+ $Y2=0.895
cc_40 N_GND_M1007_b N_A_27_565#_c_217_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.625
cc_41 N_GND_M1007_b N_A_27_565#_c_218_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.625
cc_42 N_GND_M1007_b N_A_27_565#_c_219_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.585
cc_43 N_GND_M1007_b N_A_27_565#_c_220_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.625
cc_44 N_GND_M1007_b N_A_27_565#_c_221_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.285
cc_45 N_GND_M1007_b N_A_27_565#_c_222_n 0.00953944f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.865
cc_46 N_GND_c_3_p N_A_27_565#_c_222_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.865
cc_47 N_GND_c_4_p N_A_27_565#_c_222_n 0.00475776f $X=2.38 $Y=0.19 $X2=0.69
+ $Y2=0.865
cc_48 N_GND_M1007_b N_A_27_565#_c_225_n 0.0190355f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_49 N_GND_c_11_p N_A_27_565#_c_225_n 0.00702738f $X=1.12 $Y=0.865 $X2=1.43
+ $Y2=1.675
cc_50 N_GND_M1007_b N_A_27_565#_c_227_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.675
cc_51 N_GND_M1007_b N_Y_c_331_n 0.00558158f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.865
cc_52 N_GND_c_18_p N_Y_c_331_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.865
cc_53 N_GND_c_24_p N_Y_c_331_n 8.14297e-19 $X=1.98 $Y=0.865 $X2=1.55 $Y2=0.865
cc_54 N_GND_c_4_p N_Y_c_331_n 0.00475776f $X=2.38 $Y=0.19 $X2=1.55 $Y2=0.865
cc_55 N_GND_M1007_b N_Y_c_335_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_56 N_GND_M1007_b N_Y_c_336_n 0.00656459f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.865
cc_57 N_GND_c_24_p N_Y_c_336_n 8.14297e-19 $X=1.98 $Y=0.865 $X2=2.41 $Y2=0.865
cc_58 N_GND_c_32_p N_Y_c_336_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.865
cc_59 N_GND_c_4_p N_Y_c_336_n 0.00475776f $X=2.38 $Y=0.19 $X2=2.41 $Y2=0.865
cc_60 N_GND_M1007_b N_Y_c_340_n 0.0152877f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.33
cc_61 N_GND_M1007_b N_Y_c_341_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.335
cc_62 N_GND_c_11_p N_Y_c_341_n 0.00134236f $X=1.12 $Y=0.865 $X2=1.55 $Y2=1.335
cc_63 N_GND_c_24_p N_Y_c_341_n 7.53951e-19 $X=1.98 $Y=0.865 $X2=1.55 $Y2=1.335
cc_64 N_GND_M1007_b N_Y_c_344_n 0.00463624f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.215
cc_65 N_GND_M1007_b Y 0.0305055f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.96
cc_66 N_GND_M1009_s N_Y_c_346_n 0.00418405f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.22
cc_67 N_GND_M1007_b N_Y_c_346_n 0.00793787f $X=-0.045 $Y=0 $X2=2.265 $Y2=1.22
cc_68 N_GND_c_24_p N_Y_c_346_n 0.0142303f $X=1.98 $Y=0.865 $X2=2.265 $Y2=1.22
cc_69 N_GND_M1007_b N_Y_c_349_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.33
cc_70 N_GND_M1007_b N_Y_c_350_n 0.00409378f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.335
cc_71 N_GND_c_24_p N_Y_c_350_n 7.53951e-19 $X=1.98 $Y=0.865 $X2=2.41 $Y2=1.335
cc_72 N_GND_c_38_p N_Y_c_350_n 0.00134236f $X=2.84 $Y=0.865 $X2=2.41 $Y2=1.335
cc_73 N_GND_M1007_b N_Y_c_353_n 0.06145f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.215
cc_74 N_VDD_M1008_b N_B_M1008_g 0.0264002f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_75 N_VDD_c_75_p N_B_M1008_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475 $Y2=3.825
cc_76 N_VDD_c_76_p N_B_M1008_g 0.00429146f $X=2.38 $Y=5.36 $X2=0.475 $Y2=3.825
cc_77 N_VDD_M1008_b N_B_c_127_n 0.00375034f $X=-0.045 $Y=2.645 $X2=0.27
+ $Y2=2.415
cc_78 N_VDD_M1008_b B 0.0108395f $X=-0.045 $Y=2.645 $X2=0.27 $Y2=2.7
cc_79 N_VDD_M1008_b N_A_M1005_g 0.0199048f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_80 N_VDD_c_75_p N_A_M1005_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905 $Y2=3.825
cc_81 N_VDD_c_81_p N_A_M1005_g 0.00362996f $X=1.12 $Y=3.885 $X2=0.905 $Y2=3.825
cc_82 N_VDD_c_76_p N_A_M1005_g 0.00429146f $X=2.38 $Y=5.36 $X2=0.905 $Y2=3.825
cc_83 N_VDD_M1008_b N_A_c_155_n 0.00153494f $X=-0.045 $Y=2.645 $X2=0.95
+ $Y2=2.125
cc_84 N_VDD_M1005_d A 0.0077995f $X=0.98 $Y=2.825 $X2=0.95 $Y2=3.07
cc_85 N_VDD_c_81_p A 0.00247404f $X=1.12 $Y=3.885 $X2=0.95 $Y2=3.07
cc_86 N_VDD_M1008_b N_A_27_565#_c_228_n 0.0174876f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.7
cc_87 N_VDD_c_81_p N_A_27_565#_c_228_n 0.00362996f $X=1.12 $Y=3.885 $X2=1.335
+ $Y2=2.7
cc_88 N_VDD_c_88_p N_A_27_565#_c_228_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335
+ $Y2=2.7
cc_89 N_VDD_c_76_p N_A_27_565#_c_228_n 0.00429146f $X=2.38 $Y=5.36 $X2=1.335
+ $Y2=2.7
cc_90 N_VDD_M1008_b N_A_27_565#_c_198_n 0.00428234f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_91 N_VDD_M1008_b N_A_27_565#_c_233_n 0.0173909f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.7
cc_92 N_VDD_c_81_p N_A_27_565#_c_233_n 3.67508e-19 $X=1.12 $Y=3.885 $X2=1.765
+ $Y2=2.7
cc_93 N_VDD_c_88_p N_A_27_565#_c_233_n 0.00500229f $X=1.895 $Y=5.397 $X2=1.765
+ $Y2=2.7
cc_94 N_VDD_c_94_p N_A_27_565#_c_233_n 0.00382402f $X=1.98 $Y=3.205 $X2=1.765
+ $Y2=2.7
cc_95 N_VDD_c_76_p N_A_27_565#_c_233_n 0.00430409f $X=2.38 $Y=5.36 $X2=1.765
+ $Y2=2.7
cc_96 N_VDD_M1008_b N_A_27_565#_c_206_n 0.00396043f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.625
cc_97 N_VDD_c_94_p N_A_27_565#_c_206_n 0.00379272f $X=1.98 $Y=3.205 $X2=2.12
+ $Y2=2.625
cc_98 N_VDD_M1008_b N_A_27_565#_c_240_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.7
cc_99 N_VDD_c_94_p N_A_27_565#_c_240_n 0.00362996f $X=1.98 $Y=3.205 $X2=2.195
+ $Y2=2.7
cc_100 N_VDD_c_100_p N_A_27_565#_c_240_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.195
+ $Y2=2.7
cc_101 N_VDD_c_76_p N_A_27_565#_c_240_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.195
+ $Y2=2.7
cc_102 N_VDD_M1008_b N_A_27_565#_c_212_n 0.00840215f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.625
cc_103 N_VDD_M1008_b N_A_27_565#_c_245_n 0.0212947f $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.7
cc_104 N_VDD_c_100_p N_A_27_565#_c_245_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.625
+ $Y2=2.7
cc_105 N_VDD_c_105_p N_A_27_565#_c_245_n 0.00751602f $X=2.84 $Y=3.205 $X2=2.625
+ $Y2=2.7
cc_106 N_VDD_c_76_p N_A_27_565#_c_245_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.625
+ $Y2=2.7
cc_107 N_VDD_M1008_b N_A_27_565#_c_217_n 0.0021704f $X=-0.045 $Y=2.645 $X2=1.352
+ $Y2=2.625
cc_108 N_VDD_M1008_b N_A_27_565#_c_218_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=1.765 $Y2=2.625
cc_109 N_VDD_M1008_b N_A_27_565#_c_220_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.195 $Y2=2.625
cc_110 N_VDD_M1008_b N_A_27_565#_c_252_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.545
cc_111 N_VDD_c_75_p N_A_27_565#_c_252_n 0.00452684f $X=1.035 $Y=5.397 $X2=0.26
+ $Y2=3.545
cc_112 N_VDD_c_76_p N_A_27_565#_c_252_n 0.00435496f $X=2.38 $Y=5.36 $X2=0.26
+ $Y2=3.545
cc_113 N_VDD_M1008_b N_A_27_565#_c_221_n 0.00106577f $X=-0.045 $Y=2.645 $X2=0.61
+ $Y2=3.285
cc_114 N_VDD_M1008_b N_Y_c_335_n 0.00410619f $X=-0.045 $Y=2.645 $X2=1.55
+ $Y2=2.33
cc_115 N_VDD_c_88_p N_Y_c_335_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.33
cc_116 N_VDD_c_76_p N_Y_c_335_n 0.00434939f $X=2.38 $Y=5.36 $X2=1.55 $Y2=2.33
cc_117 N_VDD_M1008_b N_Y_c_340_n 0.0042387f $X=-0.045 $Y=2.645 $X2=2.41 $Y2=2.33
cc_118 N_VDD_c_100_p N_Y_c_340_n 0.0045126f $X=2.755 $Y=5.397 $X2=2.41 $Y2=2.33
cc_119 N_VDD_c_76_p N_Y_c_340_n 0.00434939f $X=2.38 $Y=5.36 $X2=2.41 $Y2=2.33
cc_120 N_VDD_c_94_p N_Y_c_349_n 0.00634153f $X=1.98 $Y=3.205 $X2=2.265 $Y2=2.33
cc_121 N_B_M1007_g N_A_M1002_g 0.0430073f $X=0.475 $Y=0.895 $X2=0.905 $Y2=0.895
cc_122 N_B_c_126_n N_A_M1005_g 0.112923f $X=0.475 $Y=2.415 $X2=0.905 $Y2=3.825
cc_123 N_B_M1007_g N_A_c_154_n 0.0148656f $X=0.475 $Y=0.895 $X2=0.95 $Y2=2.125
cc_124 N_B_M1007_g N_A_c_155_n 0.00121111f $X=0.475 $Y=0.895 $X2=0.95 $Y2=2.125
cc_125 N_B_M1008_g N_A_27_565#_c_256_n 0.0142177f $X=0.475 $Y=3.825 $X2=0.525
+ $Y2=3.37
cc_126 B N_A_27_565#_c_256_n 0.00520961f $X=0.27 $Y=2.7 $X2=0.525 $Y2=3.37
cc_127 N_B_c_127_n N_A_27_565#_c_258_n 0.00369517f $X=0.27 $Y=2.415 $X2=0.345
+ $Y2=3.37
cc_128 B N_A_27_565#_c_258_n 0.00431991f $X=0.27 $Y=2.7 $X2=0.345 $Y2=3.37
cc_129 N_B_M1007_g N_A_27_565#_c_221_n 0.0231435f $X=0.475 $Y=0.895 $X2=0.61
+ $Y2=3.285
cc_130 N_B_M1008_g N_A_27_565#_c_221_n 0.026563f $X=0.475 $Y=3.825 $X2=0.61
+ $Y2=3.285
cc_131 N_B_c_126_n N_A_27_565#_c_221_n 0.00764878f $X=0.475 $Y=2.415 $X2=0.61
+ $Y2=3.285
cc_132 N_B_c_127_n N_A_27_565#_c_221_n 0.0350086f $X=0.27 $Y=2.415 $X2=0.61
+ $Y2=3.285
cc_133 B N_A_27_565#_c_221_n 0.00758489f $X=0.27 $Y=2.7 $X2=0.61 $Y2=3.285
cc_134 N_B_M1007_g N_A_27_565#_c_222_n 0.00996235f $X=0.475 $Y=0.895 $X2=0.69
+ $Y2=0.865
cc_135 N_B_M1007_g N_A_27_565#_c_227_n 0.0113001f $X=0.475 $Y=0.895 $X2=0.65
+ $Y2=1.675
cc_136 N_A_M1002_g N_A_27_565#_M1004_g 0.0337969f $X=0.905 $Y=0.895 $X2=1.335
+ $Y2=0.895
cc_137 A N_A_27_565#_c_228_n 0.00374181f $X=0.95 $Y=3.07 $X2=1.335 $Y2=2.7
cc_138 N_A_M1005_g N_A_27_565#_c_197_n 0.00914307f $X=0.905 $Y=3.825 $X2=1.37
+ $Y2=2.55
cc_139 N_A_c_154_n N_A_27_565#_c_197_n 0.0204279f $X=0.95 $Y=2.125 $X2=1.37
+ $Y2=2.55
cc_140 N_A_c_155_n N_A_27_565#_c_197_n 0.00375034f $X=0.95 $Y=2.125 $X2=1.37
+ $Y2=2.55
cc_141 N_A_M1002_g N_A_27_565#_c_205_n 0.0119161f $X=0.905 $Y=0.895 $X2=1.84
+ $Y2=1.585
cc_142 N_A_M1005_g N_A_27_565#_c_217_n 0.0554147f $X=0.905 $Y=3.825 $X2=1.352
+ $Y2=2.625
cc_143 N_A_c_155_n N_A_27_565#_c_217_n 0.00358357f $X=0.95 $Y=2.125 $X2=1.352
+ $Y2=2.625
cc_144 N_A_M1005_g N_A_27_565#_c_256_n 0.00457566f $X=0.905 $Y=3.825 $X2=0.525
+ $Y2=3.37
cc_145 N_A_M1002_g N_A_27_565#_c_221_n 0.00429604f $X=0.905 $Y=0.895 $X2=0.61
+ $Y2=3.285
cc_146 N_A_M1005_g N_A_27_565#_c_221_n 0.00776428f $X=0.905 $Y=3.825 $X2=0.61
+ $Y2=3.285
cc_147 N_A_c_154_n N_A_27_565#_c_221_n 0.0021255f $X=0.95 $Y=2.125 $X2=0.61
+ $Y2=3.285
cc_148 N_A_c_155_n N_A_27_565#_c_221_n 0.0822139f $X=0.95 $Y=2.125 $X2=0.61
+ $Y2=3.285
cc_149 A N_A_27_565#_c_221_n 0.00866797f $X=0.95 $Y=3.07 $X2=0.61 $Y2=3.285
cc_150 N_A_M1002_g N_A_27_565#_c_222_n 0.00996235f $X=0.905 $Y=0.895 $X2=0.69
+ $Y2=0.865
cc_151 N_A_M1002_g N_A_27_565#_c_225_n 0.0163305f $X=0.905 $Y=0.895 $X2=1.43
+ $Y2=1.675
cc_152 N_A_c_154_n N_A_27_565#_c_225_n 0.00276813f $X=0.95 $Y=2.125 $X2=1.43
+ $Y2=1.675
cc_153 N_A_c_155_n N_A_27_565#_c_225_n 0.0114342f $X=0.95 $Y=2.125 $X2=1.43
+ $Y2=1.675
cc_154 A A_110_565# 0.0123256f $X=0.95 $Y=3.07 $X2=0.55 $Y2=2.825
cc_155 N_A_c_155_n N_Y_c_335_n 0.0206732f $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.33
cc_156 A N_Y_c_335_n 0.00659455f $X=0.95 $Y=3.07 $X2=1.55 $Y2=2.33
cc_157 N_A_M1002_g N_Y_c_341_n 8.23842e-19 $X=0.905 $Y=0.895 $X2=1.55 $Y2=1.335
cc_158 N_A_c_154_n N_Y_c_344_n 3.73261e-19 $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.215
cc_159 N_A_c_155_n N_Y_c_344_n 0.0059581f $X=0.95 $Y=2.125 $X2=1.55 $Y2=2.215
cc_160 N_A_M1002_g Y 6.73508e-19 $X=0.905 $Y=0.895 $X2=1.555 $Y2=1.96
cc_161 N_A_c_155_n Y 0.00825539f $X=0.95 $Y=2.125 $X2=1.555 $Y2=1.96
cc_162 N_A_27_565#_c_256_n A_110_565# 0.00613297f $X=0.525 $Y=3.37 $X2=0.55
+ $Y2=2.825
cc_163 N_A_27_565#_c_221_n A_110_565# 0.00377193f $X=0.61 $Y=3.285 $X2=0.55
+ $Y2=2.825
cc_164 N_A_27_565#_M1004_g N_Y_c_331_n 0.00339663f $X=1.335 $Y=0.895 $X2=1.55
+ $Y2=0.865
cc_165 N_A_27_565#_M1009_g N_Y_c_331_n 0.00339663f $X=1.765 $Y=0.895 $X2=1.55
+ $Y2=0.865
cc_166 N_A_27_565#_c_205_n N_Y_c_331_n 0.00171364f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=0.865
cc_167 N_A_27_565#_c_225_n N_Y_c_331_n 0.00520269f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.865
cc_168 N_A_27_565#_c_228_n N_Y_c_335_n 0.00234922f $X=1.335 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_169 N_A_27_565#_c_197_n N_Y_c_335_n 0.00744772f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_170 N_A_27_565#_c_198_n N_Y_c_335_n 0.0168228f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_171 N_A_27_565#_c_233_n N_Y_c_335_n 0.00401146f $X=1.765 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_172 N_A_27_565#_c_205_n N_Y_c_335_n 0.0013767f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.33
cc_173 N_A_27_565#_c_225_n N_Y_c_335_n 0.00273485f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_174 N_A_27_565#_M1010_g N_Y_c_336_n 0.00339663f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=0.865
cc_175 N_A_27_565#_c_211_n N_Y_c_336_n 0.00280419f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=0.865
cc_176 N_A_27_565#_M1011_g N_Y_c_336_n 0.00339663f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=0.865
cc_177 N_A_27_565#_c_240_n N_Y_c_340_n 0.00401146f $X=2.195 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_178 N_A_27_565#_c_211_n N_Y_c_340_n 0.00250559f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.33
cc_179 N_A_27_565#_c_212_n N_Y_c_340_n 0.0206674f $X=2.55 $Y=2.625 $X2=2.41
+ $Y2=2.33
cc_180 N_A_27_565#_c_245_n N_Y_c_340_n 0.00401146f $X=2.625 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_181 N_A_27_565#_M1004_g N_Y_c_341_n 0.00542903f $X=1.335 $Y=0.895 $X2=1.55
+ $Y2=1.335
cc_182 N_A_27_565#_M1009_g N_Y_c_341_n 0.00259902f $X=1.765 $Y=0.895 $X2=1.55
+ $Y2=1.335
cc_183 N_A_27_565#_c_225_n N_Y_c_341_n 0.00238892f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=1.335
cc_184 N_A_27_565#_c_197_n N_Y_c_344_n 0.00821104f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.215
cc_185 N_A_27_565#_c_198_n N_Y_c_344_n 0.00229755f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.215
cc_186 N_A_27_565#_c_205_n N_Y_c_344_n 0.00174847f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.215
cc_187 N_A_27_565#_c_225_n N_Y_c_344_n 0.00181779f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.215
cc_188 N_A_27_565#_M1004_g Y 0.00251111f $X=1.335 $Y=0.895 $X2=1.555 $Y2=1.96
cc_189 N_A_27_565#_c_197_n Y 0.00892438f $X=1.37 $Y=2.55 $X2=1.555 $Y2=1.96
cc_190 N_A_27_565#_M1009_g Y 0.00251111f $X=1.765 $Y=0.895 $X2=1.555 $Y2=1.96
cc_191 N_A_27_565#_c_205_n Y 0.012793f $X=1.84 $Y=1.585 $X2=1.555 $Y2=1.96
cc_192 N_A_27_565#_c_225_n Y 0.0147088f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_193 N_A_27_565#_M1009_g N_Y_c_346_n 0.0130095f $X=1.765 $Y=0.895 $X2=2.265
+ $Y2=1.22
cc_194 N_A_27_565#_c_203_n N_Y_c_346_n 0.00213861f $X=2.12 $Y=1.585 $X2=2.265
+ $Y2=1.22
cc_195 N_A_27_565#_M1010_g N_Y_c_346_n 0.0130095f $X=2.195 $Y=0.895 $X2=2.265
+ $Y2=1.22
cc_196 N_A_27_565#_c_205_n N_Y_c_349_n 0.0121767f $X=1.84 $Y=1.585 $X2=2.265
+ $Y2=2.33
cc_197 N_A_27_565#_c_218_n N_Y_c_349_n 0.0158479f $X=1.765 $Y=2.625 $X2=2.265
+ $Y2=2.33
cc_198 N_A_27_565#_M1010_g N_Y_c_350_n 0.00259902f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=1.335
cc_199 N_A_27_565#_M1011_g N_Y_c_350_n 0.00939545f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=1.335
cc_200 N_A_27_565#_M1010_g N_Y_c_353_n 0.00251111f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=2.215
cc_201 N_A_27_565#_c_211_n N_Y_c_353_n 0.0184054f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_202 N_A_27_565#_M1011_g N_Y_c_353_n 0.00251111f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=2.215
cc_203 N_A_27_565#_c_219_n N_Y_c_353_n 0.00140336f $X=2.195 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_204 N_A_27_565#_c_220_n N_Y_c_353_n 0.00372651f $X=2.195 $Y=2.625 $X2=2.41
+ $Y2=2.215
