* File: sky130_osu_sc_18T_ms__inv_3.pxi.spice
* Created: Thu Oct 29 17:29:56 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__INV_3%GND N_GND_M1000_d N_GND_M1002_d N_GND_M1000_b
+ N_GND_c_2_p N_GND_c_9_p N_GND_c_3_p N_GND_c_17_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_MS__INV_3%GND
x_PM_SKY130_OSU_SC_18T_MS__INV_3%VDD N_VDD_M1001_d N_VDD_M1003_d N_VDD_M1001_b
+ N_VDD_c_47_p N_VDD_c_52_p N_VDD_c_48_p N_VDD_c_59_p VDD N_VDD_c_49_p
+ PM_SKY130_OSU_SC_18T_MS__INV_3%VDD
x_PM_SKY130_OSU_SC_18T_MS__INV_3%A N_A_c_79_n N_A_M1000_g N_A_c_83_n N_A_c_106_n
+ N_A_M1001_g N_A_c_84_n N_A_c_85_n N_A_c_86_n N_A_M1002_g N_A_c_111_n
+ N_A_M1003_g N_A_c_90_n N_A_c_92_n N_A_c_93_n N_A_M1004_g N_A_c_117_n
+ N_A_M1005_g N_A_c_97_n N_A_c_98_n N_A_c_99_n N_A_c_100_n N_A_c_101_n
+ N_A_c_102_n N_A_c_103_n A N_A_c_104_n N_A_c_105_n
+ PM_SKY130_OSU_SC_18T_MS__INV_3%A
x_PM_SKY130_OSU_SC_18T_MS__INV_3%Y N_Y_M1000_s N_Y_M1004_s N_Y_M1001_s
+ N_Y_M1005_s N_Y_c_175_n N_Y_c_193_n Y N_Y_c_179_n N_Y_c_194_n N_Y_c_181_n
+ N_Y_c_183_n N_Y_c_197_n N_Y_c_184_n N_Y_c_185_n N_Y_c_189_n
+ PM_SKY130_OSU_SC_18T_MS__INV_3%Y
cc_1 N_GND_M1000_b N_A_c_79_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.7
cc_2 N_GND_c_2_p N_A_c_79_n 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.7
cc_3 N_GND_c_3_p N_A_c_79_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.7
cc_4 N_GND_c_4_p N_A_c_79_n 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=1.7
cc_5 N_GND_M1000_b N_A_c_83_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.81
cc_6 N_GND_M1000_b N_A_c_84_n 0.0162043f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.775
cc_7 N_GND_M1000_b N_A_c_85_n 0.0114349f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.885
cc_8 N_GND_M1000_b N_A_c_86_n 0.0166526f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.7
cc_9 N_GND_c_9_p N_A_c_86_n 0.00356864f $X=1.12 $Y=0.825 $X2=0.905 $Y2=1.7
cc_10 N_GND_c_3_p N_A_c_86_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.7
cc_11 N_GND_c_4_p N_A_c_86_n 0.00468827f $X=1.02 $Y=0.17 $X2=0.905 $Y2=1.7
cc_12 N_GND_M1000_b N_A_c_90_n 0.037872f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.775
cc_13 N_GND_c_9_p N_A_c_90_n 0.00283047f $X=1.12 $Y=0.825 $X2=1.26 $Y2=1.775
cc_14 N_GND_M1000_b N_A_c_92_n 0.0305509f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.885
cc_15 N_GND_M1000_b N_A_c_93_n 0.0225344f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.7
cc_16 N_GND_c_9_p N_A_c_93_n 0.00356864f $X=1.12 $Y=0.825 $X2=1.335 $Y2=1.7
cc_17 N_GND_c_17_p N_A_c_93_n 0.00606474f $X=1.12 $Y=0.152 $X2=1.335 $Y2=1.7
cc_18 N_GND_c_4_p N_A_c_93_n 0.00468827f $X=1.02 $Y=0.17 $X2=1.335 $Y2=1.7
cc_19 N_GND_M1000_b N_A_c_97_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.775
cc_20 N_GND_M1000_b N_A_c_98_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.885
cc_21 N_GND_M1000_b N_A_c_99_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.775
cc_22 N_GND_M1000_b N_A_c_100_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.885
cc_23 N_GND_M1000_b N_A_c_101_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.305
cc_24 N_GND_M1000_b N_A_c_102_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_25 N_GND_M1000_b N_A_c_103_n 0.0348407f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_26 N_GND_M1000_b N_A_c_104_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.33
cc_27 N_GND_M1000_b N_A_c_105_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.14
cc_28 N_GND_M1000_b N_Y_c_175_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.595
cc_29 N_GND_c_2_p N_Y_c_175_n 0.00134236f $X=0.26 $Y=0.825 $X2=0.69 $Y2=1.595
cc_30 N_GND_c_9_p N_Y_c_175_n 7.53951e-19 $X=1.12 $Y=0.825 $X2=0.69 $Y2=1.595
cc_31 N_GND_M1000_b Y 0.0456345f $X=-0.045 $Y=0 $X2=0.76 $Y2=2.2
cc_32 N_GND_M1002_d N_Y_c_179_n 0.0127699f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1.48
cc_33 N_GND_c_9_p N_Y_c_179_n 0.0142303f $X=1.12 $Y=0.825 $X2=1.405 $Y2=1.48
cc_34 N_GND_M1000_b N_Y_c_181_n 0.0142042f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.595
cc_35 N_GND_c_9_p N_Y_c_181_n 7.53951e-19 $X=1.12 $Y=0.825 $X2=1.55 $Y2=1.595
cc_36 N_GND_M1000_b N_Y_c_183_n 0.0950169f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.845
cc_37 N_GND_M1000_b N_Y_c_184_n 0.00312976f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.96
cc_38 N_GND_M1000_b N_Y_c_185_n 0.00155118f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_39 N_GND_c_9_p N_Y_c_185_n 8.14297e-19 $X=1.12 $Y=0.825 $X2=0.69 $Y2=0.825
cc_40 N_GND_c_3_p N_Y_c_185_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.825
cc_41 N_GND_c_4_p N_Y_c_185_n 0.00475776f $X=1.02 $Y=0.17 $X2=0.69 $Y2=0.825
cc_42 N_GND_M1000_b N_Y_c_189_n 0.00156053f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_43 N_GND_c_9_p N_Y_c_189_n 8.14297e-19 $X=1.12 $Y=0.825 $X2=1.55 $Y2=0.825
cc_44 N_GND_c_17_p N_Y_c_189_n 0.00757793f $X=1.12 $Y=0.152 $X2=1.55 $Y2=0.825
cc_45 N_GND_c_4_p N_Y_c_189_n 0.00476261f $X=1.02 $Y=0.17 $X2=1.55 $Y2=0.825
cc_46 N_VDD_M1001_b N_A_c_106_n 0.0181616f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=2.96
cc_47 N_VDD_c_47_p N_A_c_106_n 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=2.96
cc_48 N_VDD_c_48_p N_A_c_106_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=2.96
cc_49 N_VDD_c_49_p N_A_c_106_n 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=2.96
cc_50 N_VDD_M1001_b N_A_c_85_n 0.00448664f $X=-0.045 $Y=2.905 $X2=0.83 $Y2=2.885
cc_51 N_VDD_M1001_b N_A_c_111_n 0.0159283f $X=-0.045 $Y=2.905 $X2=0.905 $Y2=2.96
cc_52 N_VDD_c_52_p N_A_c_111_n 0.00354579f $X=1.12 $Y=3.455 $X2=0.905 $Y2=2.96
cc_53 N_VDD_c_48_p N_A_c_111_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=2.96
cc_54 N_VDD_c_49_p N_A_c_111_n 0.00468827f $X=1.02 $Y=6.49 $X2=0.905 $Y2=2.96
cc_55 N_VDD_M1001_b N_A_c_92_n 0.00774816f $X=-0.045 $Y=2.905 $X2=1.26 $Y2=2.885
cc_56 N_VDD_c_52_p N_A_c_92_n 0.00341318f $X=1.12 $Y=3.455 $X2=1.26 $Y2=2.885
cc_57 N_VDD_M1001_b N_A_c_117_n 0.0221472f $X=-0.045 $Y=2.905 $X2=1.335 $Y2=2.96
cc_58 N_VDD_c_52_p N_A_c_117_n 0.00354579f $X=1.12 $Y=3.455 $X2=1.335 $Y2=2.96
cc_59 N_VDD_c_59_p N_A_c_117_n 0.00606474f $X=1.12 $Y=6.507 $X2=1.335 $Y2=2.96
cc_60 N_VDD_c_49_p N_A_c_117_n 0.00468827f $X=1.02 $Y=6.49 $X2=1.335 $Y2=2.96
cc_61 N_VDD_M1001_b N_A_c_98_n 0.00244521f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.885
cc_62 N_VDD_M1001_b N_A_c_100_n 8.75564e-19 $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=2.885
cc_63 N_VDD_M1001_d A 0.0162774f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.325
cc_64 N_VDD_c_47_p A 0.00522047f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.325
cc_65 N_VDD_c_52_p A 9.09141e-19 $X=1.12 $Y=3.455 $X2=0.32 $Y2=3.325
cc_66 N_VDD_M1001_d N_A_c_104_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_67 N_VDD_M1001_b N_A_c_104_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=3.33
cc_68 N_VDD_c_47_p N_A_c_104_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_69 N_VDD_M1001_b N_Y_c_193_n 0.00248543f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=2.845
cc_70 N_VDD_M1001_b N_Y_c_194_n 0.00520877f $X=-0.045 $Y=2.905 $X2=1.405
+ $Y2=2.96
cc_71 N_VDD_c_52_p N_Y_c_194_n 0.0090257f $X=1.12 $Y=3.455 $X2=1.405 $Y2=2.96
cc_72 N_VDD_M1001_b N_Y_c_183_n 0.0111011f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.845
cc_73 N_VDD_M1001_b N_Y_c_197_n 0.00361433f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_74 N_VDD_c_48_p N_Y_c_197_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69 $Y2=2.96
cc_75 N_VDD_c_49_p N_Y_c_197_n 0.00475776f $X=1.02 $Y=6.49 $X2=0.69 $Y2=2.96
cc_76 N_VDD_M1001_b N_Y_c_184_n 0.00745764f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.96
cc_77 N_VDD_c_59_p N_Y_c_184_n 0.00757793f $X=1.12 $Y=6.507 $X2=1.55 $Y2=2.96
cc_78 N_VDD_c_49_p N_Y_c_184_n 0.00476261f $X=1.02 $Y=6.49 $X2=1.55 $Y2=2.96
cc_79 A N_Y_M1001_s 0.00251573f $X=0.32 $Y=3.325 $X2=0.55 $Y2=3.085
cc_80 N_A_c_79_n N_Y_c_175_n 0.00942005f $X=0.475 $Y=1.7 $X2=0.69 $Y2=1.595
cc_81 N_A_c_86_n N_Y_c_175_n 0.00259753f $X=0.905 $Y=1.7 $X2=0.69 $Y2=1.595
cc_82 N_A_c_103_n N_Y_c_175_n 6.32153e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=1.595
cc_83 N_A_c_106_n N_Y_c_193_n 0.00169643f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.845
cc_84 N_A_c_85_n N_Y_c_193_n 0.00259868f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.845
cc_85 N_A_c_111_n N_Y_c_193_n 0.00144225f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.845
cc_86 N_A_c_98_n N_Y_c_193_n 0.00102602f $X=0.475 $Y=2.885 $X2=0.69 $Y2=2.845
cc_87 N_A_c_100_n N_Y_c_193_n 0.00150284f $X=0.905 $Y=2.885 $X2=0.69 $Y2=2.845
cc_88 N_A_c_102_n N_Y_c_193_n 0.00173027f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.845
cc_89 N_A_c_103_n N_Y_c_193_n 2.98633e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.845
cc_90 A N_Y_c_193_n 0.00815006f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.845
cc_91 N_A_c_104_n N_Y_c_193_n 0.0071561f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.845
cc_92 N_A_c_79_n Y 0.00150089f $X=0.475 $Y=1.7 $X2=0.76 $Y2=2.2
cc_93 N_A_c_83_n Y 0.00792324f $X=0.475 $Y=2.81 $X2=0.76 $Y2=2.2
cc_94 N_A_c_84_n Y 0.0163225f $X=0.83 $Y=1.775 $X2=0.76 $Y2=2.2
cc_95 N_A_c_85_n Y 0.0038871f $X=0.83 $Y=2.885 $X2=0.76 $Y2=2.2
cc_96 N_A_c_86_n Y 0.00150089f $X=0.905 $Y=1.7 $X2=0.76 $Y2=2.2
cc_97 N_A_c_102_n Y 0.0178517f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_98 N_A_c_103_n Y 0.00610708f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_99 N_A_c_104_n Y 0.0182346f $X=0.32 $Y=3.33 $X2=0.76 $Y2=2.2
cc_100 N_A_c_105_n Y 0.00675469f $X=0.535 $Y=2.14 $X2=0.76 $Y2=2.2
cc_101 N_A_c_86_n N_Y_c_179_n 0.0130014f $X=0.905 $Y=1.7 $X2=1.405 $Y2=1.48
cc_102 N_A_c_90_n N_Y_c_179_n 0.0022289f $X=1.26 $Y=1.775 $X2=1.405 $Y2=1.48
cc_103 N_A_c_93_n N_Y_c_179_n 0.0129682f $X=1.335 $Y=1.7 $X2=1.405 $Y2=1.48
cc_104 N_A_c_111_n N_Y_c_194_n 0.0069535f $X=0.905 $Y=2.96 $X2=1.405 $Y2=2.96
cc_105 N_A_c_92_n N_Y_c_194_n 0.0176406f $X=1.26 $Y=2.885 $X2=1.405 $Y2=2.96
cc_106 N_A_c_117_n N_Y_c_194_n 0.00693713f $X=1.335 $Y=2.96 $X2=1.405 $Y2=2.96
cc_107 N_A_c_100_n N_Y_c_194_n 0.00560085f $X=0.905 $Y=2.885 $X2=1.405 $Y2=2.96
cc_108 N_A_c_93_n N_Y_c_181_n 0.00401708f $X=1.335 $Y=1.7 $X2=1.55 $Y2=1.595
cc_109 N_A_c_92_n N_Y_c_183_n 0.00397242f $X=1.26 $Y=2.885 $X2=1.55 $Y2=2.845
cc_110 N_A_c_93_n N_Y_c_183_n 0.00700756f $X=1.335 $Y=1.7 $X2=1.55 $Y2=2.845
cc_111 N_A_c_117_n N_Y_c_183_n 0.00214586f $X=1.335 $Y=2.96 $X2=1.55 $Y2=2.845
cc_112 N_A_c_106_n N_Y_c_197_n 0.00199065f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.96
cc_113 N_A_c_85_n N_Y_c_197_n 0.00864247f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.96
cc_114 N_A_c_111_n N_Y_c_197_n 0.0035213f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.96
cc_115 N_A_c_102_n N_Y_c_197_n 0.00165526f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_116 N_A_c_103_n N_Y_c_197_n 2.38128e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_117 A N_Y_c_197_n 0.00938699f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.96
cc_118 N_A_c_104_n N_Y_c_197_n 0.0226156f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_119 N_A_c_92_n N_Y_c_184_n 0.011693f $X=1.26 $Y=2.885 $X2=1.55 $Y2=2.96
cc_120 N_A_c_79_n N_Y_c_185_n 0.00231637f $X=0.475 $Y=1.7 $X2=0.69 $Y2=0.825
cc_121 N_A_c_84_n N_Y_c_185_n 0.00256118f $X=0.83 $Y=1.775 $X2=0.69 $Y2=0.825
cc_122 N_A_c_86_n N_Y_c_185_n 0.00231637f $X=0.905 $Y=1.7 $X2=0.69 $Y2=0.825
cc_123 N_A_c_102_n N_Y_c_185_n 0.00110256f $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_124 N_A_c_93_n N_Y_c_189_n 0.0057847f $X=1.335 $Y=1.7 $X2=1.55 $Y2=0.825
