* File: sky130_osu_sc_15T_ls__nand2_l.pex.spice
* Created: Fri Nov 12 14:58:30 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__NAND2_L%GND 1 17 19 26 33 36
r24 33 36 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r25 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r26 17 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r27 17 24 4.26217 $w=1.7e-07 $l=2.14243e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=1.05 $Y2=0.305
r28 17 19 3.29607 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=1.197 $Y=0.152
+ $X2=0.965 $Y2=0.152
r29 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r30 1 26 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NAND2_L%VDD 1 2 17 21 23 30 35 38
r15 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r16 28 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r17 26 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r18 24 33 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r19 24 26 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r20 23 28 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.245
r21 23 26 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r22 19 33 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r23 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r24 17 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r25 17 33 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r26 2 30 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=3.565 $X2=1.12 $Y2=4.565
r27 1 21 600 $w=1.7e-07 $l=1.06066e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.565
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NAND2_L%A 3 7 10 14 20
r27 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r28 14 17 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.32 $Y=2.425
+ $X2=0.32 $Y2=3.07
r29 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=2.425 $X2=0.32 $Y2=2.425
r30 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.425
+ $X2=0.367 $Y2=2.59
r31 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=2.425
+ $X2=0.367 $Y2=2.26
r32 7 12 822.989 $w=1.5e-07 $l=1.605e-06 $layer=POLY_cond $X=0.475 $Y=4.195
+ $X2=0.475 $Y2=2.59
r33 3 11 730.691 $w=1.5e-07 $l=1.425e-06 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NAND2_L%B 3 7 10 14 19 22
c35 10 0 1.91696e-19 $X=0.915 $Y=1.675
c36 3 0 1.57512e-19 $X=0.835 $Y=0.835
r37 17 19 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.915 $Y=1.675
+ $X2=1.06 $Y2=1.675
r38 14 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.06 $Y=2.7 $X2=1.06
+ $Y2=2.7
r39 12 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.76
+ $X2=1.06 $Y2=1.675
r40 12 14 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.06 $Y=1.76
+ $X2=1.06 $Y2=2.7
r41 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=1.675 $X2=0.915 $Y2=1.675
r42 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=1.51
r43 5 10 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.84
+ $X2=0.905 $Y2=1.675
r44 5 7 1207.56 $w=1.5e-07 $l=2.355e-06 $layer=POLY_cond $X=0.905 $Y=1.84
+ $X2=0.905 $Y2=4.195
r45 3 11 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.835 $Y=0.835
+ $X2=0.835 $Y2=1.51
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__NAND2_L%Y 1 3 10 16 21 22 26 32
c37 22 0 1.57512e-19 $X=0.405 $Y=1.22
c38 16 0 1.91696e-19 $X=0.69 $Y=2.33
r39 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.215
+ $X2=0.69 $Y2=2.33
r40 24 26 0.12036 $w=1.7e-07 $l=1.25e-07 $layer=MET1_cond $X=0.69 $Y=2.215
+ $X2=0.69 $Y2=2.09
r41 23 26 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=0.69 $Y=1.305
+ $X2=0.69 $Y2=2.09
r42 22 29 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=1.22
+ $X2=0.26 $Y2=1.22
r43 21 23 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=1.22
+ $X2=0.69 $Y2=1.305
r44 21 22 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=1.22
+ $X2=0.405 $Y2=1.22
r45 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.33
+ $X2=0.69 $Y2=2.33
r46 16 19 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=0.69 $Y=2.33
+ $X2=0.69 $Y2=4.565
r47 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.22
+ $X2=0.26 $Y2=1.22
r48 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.26 $Y=0.74
+ $X2=0.26 $Y2=1.22
r49 3 19 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.565 $X2=0.69 $Y2=4.565
r50 1 10 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

