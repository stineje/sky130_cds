* File: sky130_osu_sc_12T_ms__and2_1.pex.spice
* Created: Fri Nov 12 15:20:09 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__AND2_1%GND 1 17 19 26 35 38
r36 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r37 24 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.755
r38 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r39 17 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r40 17 19 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r41 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r42 1 26 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.91 $Y=0.575
+ $X2=1.05 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_1%VDD 1 2 17 21 23 30 36 38 41
r29 38 41 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r30 28 36 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r31 28 30 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.295
r32 26 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r33 24 35 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r34 24 26 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r35 23 36 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r36 23 26 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r37 19 35 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r38 19 21 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135 $X2=0.26
+ $Y2=3.635
r39 17 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r40 17 35 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r41 2 30 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.295
r42 1 21 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_1%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=2.85
+ $X2=0.275 $Y2=2.85
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.85
+ $X2=0.27 $Y2=2.85
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.285
+ $X2=0.27 $Y2=2.85
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.285 $X2=0.27 $Y2=2.285
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.285
+ $X2=0.475 $Y2=2.285
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.45
+ $X2=0.475 $Y2=2.285
r38 5 7 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.475 $Y=2.45
+ $X2=0.475 $Y2=3.235
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=2.285
r40 1 3 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_1%B 3 7 10 14 22
r41 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.48
+ $X2=0.955 $Y2=2.48
r42 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.48
+ $X2=0.95 $Y2=2.48
r43 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=1.945
+ $X2=0.95 $Y2=2.48
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.945 $X2=0.95 $Y2=1.945
r45 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=1.945
+ $X2=0.922 $Y2=2.11
r46 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=1.945
+ $X2=0.922 $Y2=1.78
r47 7 12 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.11
r48 3 11 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.835 $Y=0.835
+ $X2=0.835 $Y2=1.78
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_1%A_27_115# 1 3 11 15 16 18 19 24 26 27 32
+ 36 38 39 40
r69 39 40 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.065
+ $X2=0.65 $Y2=3.235
r70 34 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.455
+ $X2=0.61 $Y2=1.455
r71 34 36 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.455
+ $X2=1.43 $Y2=1.455
r72 32 40 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.69 $Y=3.295 $X2=0.69
+ $Y2=3.235
r73 28 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.54 $X2=0.61
+ $Y2=1.455
r74 28 39 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=3.065
r75 26 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.455
+ $X2=0.61 $Y2=1.455
r76 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.455
+ $X2=0.345 $Y2=1.455
r77 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.345 $Y2=1.455
r78 22 24 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r79 21 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.455 $X2=1.43 $Y2=1.455
r80 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.33
+ $X2=1.352 $Y2=2.48
r81 16 21 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.412 $Y2=1.455
r82 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=2.33
r83 15 19 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=3.235
+ $X2=1.335 $Y2=2.48
r84 9 21 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.412 $Y2=1.455
r85 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.835
r86 3 32 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.295
r87 1 24 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__AND2_1%Y 1 3 10 16 26 29 32
r35 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=2.11
r36 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=1.74
r37 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r38 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.74
r39 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r40 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.11
r41 16 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.955
r42 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r43 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r44 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r45 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r46 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41 $Y=0.575
+ $X2=1.55 $Y2=0.755
.ends

