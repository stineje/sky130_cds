magic
tech sky130A
magscale 1 2
timestamp 1612373574
<< nwell >>
rect -9 529 286 1119
<< nmoslvt >>
rect 80 115 110 225
rect 166 115 196 225
<< pmos >>
rect 80 713 110 965
rect 152 713 182 965
<< ndiff >>
rect 27 165 80 225
rect 27 131 35 165
rect 69 131 80 165
rect 27 115 80 131
rect 110 165 166 225
rect 110 131 121 165
rect 155 131 166 165
rect 110 115 166 131
rect 196 165 249 225
rect 196 131 207 165
rect 241 131 249 165
rect 196 115 249 131
<< pdiff >>
rect 27 949 80 965
rect 27 809 35 949
rect 69 809 80 949
rect 27 713 80 809
rect 110 713 152 965
rect 182 949 235 965
rect 182 809 193 949
rect 227 809 235 949
rect 182 713 235 809
<< ndiffc >>
rect 35 131 69 165
rect 121 131 155 165
rect 207 131 241 165
<< pdiffc >>
rect 35 809 69 949
rect 193 809 227 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 152 965 182 991
rect 80 399 110 713
rect 152 532 182 713
rect 152 516 225 532
rect 152 482 181 516
rect 215 482 225 516
rect 152 466 225 482
rect 56 383 110 399
rect 56 349 66 383
rect 100 349 110 383
rect 56 333 110 349
rect 80 225 110 333
rect 166 225 196 466
rect 80 89 110 115
rect 166 89 196 115
<< polycont >>
rect 181 482 215 516
rect 66 349 100 383
<< locali >>
rect 0 1089 286 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 286 1089
rect 35 949 69 965
rect 35 483 69 809
rect 193 949 227 1049
rect 193 793 227 809
rect 113 383 147 523
rect 181 516 215 597
rect 181 466 215 482
rect 50 349 66 383
rect 100 349 147 383
rect 35 165 69 181
rect 35 61 69 131
rect 121 165 155 227
rect 121 115 155 131
rect 207 165 241 181
rect 207 61 241 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 181 597 215 631
rect 35 449 69 483
rect 113 523 147 557
rect 121 227 155 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 286 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 286 1089
rect 0 1049 286 1055
rect 169 631 227 637
rect 148 597 181 631
rect 215 597 227 631
rect 169 591 227 597
rect 101 557 159 563
rect 79 523 113 557
rect 147 523 159 557
rect 101 517 159 523
rect 23 483 81 489
rect 23 449 35 483
rect 69 449 155 483
rect 23 443 81 449
rect 121 267 155 449
rect 109 261 167 267
rect 109 227 121 261
rect 155 227 167 261
rect 109 221 167 227
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 137 341 137 341 1 Y
port 1 n
rlabel viali 198 614 198 614 1 A
port 2 n
rlabel viali 130 540 130 540 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
