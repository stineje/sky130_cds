magic
tech sky130A
magscale 1 2
timestamp 1604007754
<< checkpaint >>
rect -1269 2461 1967 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1967 -1129
<< nwell >>
rect -9 529 707 1119
<< locali >>
rect 0 1049 704 1110
rect 0 0 704 61
<< metal1 >>
rect 0 1049 704 1110
rect 0 0 704 61
<< labels >>
rlabel metal1 363 26 363 26 1 gnd
rlabel metal1 374 1076 374 1076 1 vdd
<< end >>
