* File: sky130_osu_sc_12T_ms__dffr_l.pxi.spice
* Created: Fri Nov 12 15:22:47 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%GND N_GND_M1021_s N_GND_M1018_s N_GND_M1005_d
+ N_GND_M1007_s N_GND_M1027_d N_GND_M1023_d N_GND_M1012_s N_GND_M1013_d
+ N_GND_M1016_d N_GND_M1021_b N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_12_p
+ N_GND_c_47_p N_GND_c_48_p N_GND_c_49_p N_GND_c_50_p N_GND_c_51_p N_GND_c_52_p
+ N_GND_c_53_p N_GND_c_54_p N_GND_c_55_p N_GND_c_19_p N_GND_c_16_p N_GND_c_172_p
+ N_GND_c_173_p GND N_GND_c_5_p PM_SKY130_OSU_SC_12T_MS__DFFR_L%GND
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%VDD N_VDD_M1004_s N_VDD_M1002_d N_VDD_M1028_s
+ N_VDD_M1022_d N_VDD_M1009_d N_VDD_M1030_d N_VDD_M1011_d N_VDD_M1004_b
+ N_VDD_c_247_p N_VDD_c_248_p N_VDD_c_267_p N_VDD_c_273_p N_VDD_c_275_p
+ N_VDD_c_302_p N_VDD_c_288_p N_VDD_c_292_p N_VDD_c_259_p N_VDD_c_260_p
+ N_VDD_c_331_p N_VDD_c_332_p N_VDD_c_356_p VDD N_VDD_c_249_p
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%RN N_RN_M1021_g N_RN_c_380_n N_RN_M1004_g
+ N_RN_c_382_n N_RN_c_383_n RN PM_SKY130_OSU_SC_12T_MS__DFFR_L%RN
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_110_115# N_A_110_115#_M1021_d
+ N_A_110_115#_M1004_d N_A_110_115#_c_413_n N_A_110_115#_M1018_g
+ N_A_110_115#_M1015_g N_A_110_115#_c_418_n N_A_110_115#_M1030_g
+ N_A_110_115#_c_421_n N_A_110_115#_M1013_g N_A_110_115#_c_425_n
+ N_A_110_115#_c_427_n N_A_110_115#_c_431_n N_A_110_115#_c_432_n
+ N_A_110_115#_c_433_n N_A_110_115#_c_435_n N_A_110_115#_c_436_n
+ N_A_110_115#_c_437_n N_A_110_115#_c_439_n N_A_110_115#_c_534_p
+ N_A_110_115#_c_441_n N_A_110_115#_c_461_n N_A_110_115#_c_565_p
+ N_A_110_115#_c_465_n N_A_110_115#_c_466_n
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_110_115#
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_342_442# N_A_342_442#_M1031_d
+ N_A_342_442#_M1024_d N_A_342_442#_M1002_g N_A_342_442#_M1005_g
+ N_A_342_442#_c_614_n N_A_342_442#_c_615_n N_A_342_442#_c_631_n
+ N_A_342_442#_c_616_n N_A_342_442#_c_618_n N_A_342_442#_c_620_n
+ N_A_342_442#_c_634_n N_A_342_442#_c_621_n N_A_342_442#_c_622_n
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_342_442#
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%D N_D_M1007_g N_D_M1028_g N_D_c_698_n
+ N_D_c_699_n D PM_SKY130_OSU_SC_12T_MS__DFFR_L%D
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%CK N_CK_M1024_g N_CK_M1026_g N_CK_M1019_g
+ N_CK_M1000_g N_CK_c_735_n N_CK_M1010_g N_CK_c_740_n N_CK_M1029_g N_CK_c_741_n
+ N_CK_c_742_n N_CK_c_743_n N_CK_c_744_n N_CK_c_747_n N_CK_c_748_n N_CK_c_751_n
+ N_CK_c_752_n N_CK_c_753_n N_CK_c_754_n N_CK_c_755_n N_CK_c_756_n N_CK_c_757_n
+ N_CK_c_758_n N_CK_c_759_n N_CK_c_760_n N_CK_c_761_n N_CK_c_762_n N_CK_c_763_n
+ N_CK_c_764_n CK PM_SKY130_OSU_SC_12T_MS__DFFR_L%CK
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_217_605# N_A_217_605#_M1018_d
+ N_A_217_605#_M1015_s N_A_217_605#_M1027_g N_A_217_605#_M1022_g
+ N_A_217_605#_c_990_n N_A_217_605#_c_992_n N_A_217_605#_c_993_n
+ N_A_217_605#_c_994_n N_A_217_605#_M1025_g N_A_217_605#_M1014_g
+ N_A_217_605#_c_999_n N_A_217_605#_c_1000_n N_A_217_605#_c_1001_n
+ N_A_217_605#_c_1002_n N_A_217_605#_c_1005_n N_A_217_605#_c_1006_n
+ N_A_217_605#_c_1008_n N_A_217_605#_c_1009_n N_A_217_605#_c_1058_n
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_217_605#
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_618_89# N_A_618_89#_M1010_d
+ N_A_618_89#_M1029_d N_A_618_89#_c_1124_n N_A_618_89#_M1031_g
+ N_A_618_89#_c_1127_n N_A_618_89#_c_1128_n N_A_618_89#_c_1129_n
+ N_A_618_89#_M1017_g N_A_618_89#_c_1131_n N_A_618_89#_M1003_g
+ N_A_618_89#_c_1133_n N_A_618_89#_M1020_g N_A_618_89#_c_1137_n
+ N_A_618_89#_c_1138_n N_A_618_89#_c_1139_n N_A_618_89#_c_1140_n
+ N_A_618_89#_c_1141_n N_A_618_89#_c_1142_n N_A_618_89#_c_1157_n
+ N_A_618_89#_c_1147_n N_A_618_89#_c_1148_n N_A_618_89#_c_1161_n
+ N_A_618_89#_c_1149_n N_A_618_89#_c_1241_n N_A_618_89#_c_1150_n
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_618_89#
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_1160_89# N_A_1160_89#_M1012_d
+ N_A_1160_89#_M1006_s N_A_1160_89#_M1023_g N_A_1160_89#_M1009_g
+ N_A_1160_89#_M1016_g N_A_1160_89#_M1011_g N_A_1160_89#_c_1326_n
+ N_A_1160_89#_c_1330_n N_A_1160_89#_c_1331_n N_A_1160_89#_c_1332_n
+ N_A_1160_89#_c_1333_n N_A_1160_89#_c_1335_n N_A_1160_89#_c_1336_n
+ N_A_1160_89#_c_1337_n N_A_1160_89#_c_1338_n N_A_1160_89#_c_1339_n
+ N_A_1160_89#_c_1340_n N_A_1160_89#_c_1341_n N_A_1160_89#_c_1343_n
+ N_A_1160_89#_c_1368_n N_A_1160_89#_c_1371_n N_A_1160_89#_c_1372_n
+ N_A_1160_89#_c_1344_n N_A_1160_89#_c_1347_n N_A_1160_89#_c_1348_n
+ N_A_1160_89#_c_1349_n N_A_1160_89#_c_1350_n N_A_1160_89#_c_1351_n
+ N_A_1160_89#_c_1352_n N_A_1160_89#_c_1353_n N_A_1160_89#_c_1354_n
+ N_A_1160_89#_c_1355_n PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_1160_89#
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_998_115# N_A_998_115#_M1019_d
+ N_A_998_115#_M1003_d N_A_998_115#_M1012_g N_A_998_115#_M1006_g
+ N_A_998_115#_c_1538_n N_A_998_115#_c_1540_n N_A_998_115#_c_1585_n
+ N_A_998_115#_c_1621_n N_A_998_115#_c_1557_n N_A_998_115#_c_1541_n
+ N_A_998_115#_c_1542_n N_A_998_115#_c_1544_n N_A_998_115#_c_1547_n
+ N_A_998_115#_c_1548_n N_A_998_115#_c_1549_n N_A_998_115#_c_1551_n
+ N_A_998_115#_c_1552_n PM_SKY130_OSU_SC_12T_MS__DFFR_L%A_998_115#
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%QN N_QN_M1016_s N_QN_M1011_s N_QN_M1008_g
+ N_QN_M1001_g N_QN_c_1680_n N_QN_c_1681_n N_QN_c_1685_n N_QN_c_1686_n
+ N_QN_c_1688_n N_QN_c_1689_n N_QN_c_1690_n N_QN_c_1691_n QN
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%QN
x_PM_SKY130_OSU_SC_12T_MS__DFFR_L%Q N_Q_M1008_d N_Q_M1001_d N_Q_c_1771_n
+ N_Q_c_1775_n N_Q_c_1773_n N_Q_c_1774_n N_Q_c_1780_n Q
+ PM_SKY130_OSU_SC_12T_MS__DFFR_L%Q
cc_1 N_GND_M1021_b N_RN_M1021_g 0.0616724f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_RN_M1021_g 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_RN_M1021_g 0.00606474f $X=1.125 $Y=0.152 $X2=0.475 $Y2=0.835
cc_4 N_GND_c_4_p N_RN_M1021_g 0.00359543f $X=1.21 $Y=0.74 $X2=0.475 $Y2=0.835
cc_5 N_GND_c_5_p N_RN_M1021_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.475 $Y2=0.835
cc_6 N_GND_M1021_b N_RN_c_380_n 0.0376794f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.99
cc_7 N_GND_M1021_b N_RN_M1004_g 0.0288885f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.235
cc_8 N_GND_M1021_b N_RN_c_382_n 0.0149094f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_9 N_GND_M1021_b N_RN_c_383_n 0.020332f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.825
cc_10 N_GND_M1021_b N_A_110_115#_c_413_n 0.0181101f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=1.045
cc_11 N_GND_c_4_p N_A_110_115#_c_413_n 0.00502587f $X=1.21 $Y=0.74 $X2=1.425
+ $Y2=1.045
cc_12 N_GND_c_12_p N_A_110_115#_c_413_n 0.00606474f $X=1.985 $Y=0.152 $X2=1.425
+ $Y2=1.045
cc_13 N_GND_c_5_p N_A_110_115#_c_413_n 0.00468827f $X=9.175 $Y=0.19 $X2=1.425
+ $Y2=1.045
cc_14 N_GND_M1021_b N_A_110_115#_M1015_g 0.060904f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=3.445
cc_15 N_GND_M1021_b N_A_110_115#_c_418_n 0.0603547f $X=-0.05 $Y=0 $X2=7.615
+ $Y2=1.52
cc_16 N_GND_c_16_p N_A_110_115#_c_418_n 0.00335985f $X=7.9 $Y=0.74 $X2=7.615
+ $Y2=1.52
cc_17 N_GND_M1021_b N_A_110_115#_M1030_g 0.0560425f $X=-0.05 $Y=0 $X2=7.615
+ $Y2=3.445
cc_18 N_GND_M1021_b N_A_110_115#_c_421_n 0.0181101f $X=-0.05 $Y=0 $X2=7.685
+ $Y2=1.045
cc_19 N_GND_c_19_p N_A_110_115#_c_421_n 0.00606474f $X=7.815 $Y=0.152 $X2=7.685
+ $Y2=1.045
cc_20 N_GND_c_16_p N_A_110_115#_c_421_n 0.00502587f $X=7.9 $Y=0.74 $X2=7.685
+ $Y2=1.045
cc_21 N_GND_c_5_p N_A_110_115#_c_421_n 0.00468827f $X=9.175 $Y=0.19 $X2=7.685
+ $Y2=1.045
cc_22 N_GND_M1021_b N_A_110_115#_c_425_n 0.0450929f $X=-0.05 $Y=0 $X2=1.425
+ $Y2=1.21
cc_23 N_GND_c_4_p N_A_110_115#_c_425_n 0.00336f $X=1.21 $Y=0.74 $X2=1.425
+ $Y2=1.21
cc_24 N_GND_M1021_b N_A_110_115#_c_427_n 0.00155788f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=0.755
cc_25 N_GND_c_3_p N_A_110_115#_c_427_n 0.0075272f $X=1.125 $Y=0.152 $X2=0.69
+ $Y2=0.755
cc_26 N_GND_c_4_p N_A_110_115#_c_427_n 0.0140971f $X=1.21 $Y=0.74 $X2=0.69
+ $Y2=0.755
cc_27 N_GND_c_5_p N_A_110_115#_c_427_n 0.00474817f $X=9.175 $Y=0.19 $X2=0.69
+ $Y2=0.755
cc_28 N_GND_M1021_b N_A_110_115#_c_431_n 0.0021895f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=2.95
cc_29 N_GND_M1021_b N_A_110_115#_c_432_n 0.0188948f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.175
cc_30 N_GND_M1021_b N_A_110_115#_c_433_n 0.00886322f $X=-0.05 $Y=0 $X2=1.135
+ $Y2=1.21
cc_31 N_GND_c_4_p N_A_110_115#_c_433_n 4.91534e-19 $X=1.21 $Y=0.74 $X2=1.135
+ $Y2=1.21
cc_32 N_GND_M1021_b N_A_110_115#_c_435_n 0.0159872f $X=-0.05 $Y=0 $X2=0.955
+ $Y2=1.21
cc_33 N_GND_M1021_b N_A_110_115#_c_436_n 0.0162344f $X=-0.05 $Y=0 $X2=0.87
+ $Y2=2.26
cc_34 N_GND_M1021_b N_A_110_115#_c_437_n 0.0015072f $X=-0.05 $Y=0 $X2=1.22
+ $Y2=1.21
cc_35 N_GND_c_4_p N_A_110_115#_c_437_n 0.00797325f $X=1.21 $Y=0.74 $X2=1.22
+ $Y2=1.21
cc_36 N_GND_M1021_b N_A_110_115#_c_439_n 0.00428422f $X=-0.05 $Y=0 $X2=7.89
+ $Y2=1.21
cc_37 N_GND_c_16_p N_A_110_115#_c_439_n 0.00849521f $X=7.9 $Y=0.74 $X2=7.89
+ $Y2=1.21
cc_38 N_GND_M1018_s N_A_110_115#_c_441_n 5.79494e-19 $X=1.085 $Y=0.575 $X2=7.805
+ $Y2=1
cc_39 N_GND_M1005_d N_A_110_115#_c_441_n 0.00254601f $X=1.93 $Y=0.575 $X2=7.805
+ $Y2=1
cc_40 N_GND_M1007_s N_A_110_115#_c_441_n 0.00263312f $X=2.465 $Y=0.575 $X2=7.805
+ $Y2=1
cc_41 N_GND_M1027_d N_A_110_115#_c_441_n 0.00722605f $X=4.2 $Y=0.575 $X2=7.805
+ $Y2=1
cc_42 N_GND_M1023_d N_A_110_115#_c_441_n 0.00364862f $X=5.95 $Y=0.575 $X2=7.805
+ $Y2=1
cc_43 N_GND_M1012_s N_A_110_115#_c_441_n 0.00254601f $X=6.915 $Y=0.575 $X2=7.805
+ $Y2=1
cc_44 N_GND_M1013_d N_A_110_115#_c_441_n 0.00227813f $X=7.76 $Y=0.575 $X2=7.805
+ $Y2=1
cc_45 N_GND_M1021_b N_A_110_115#_c_441_n 0.0190105f $X=-0.05 $Y=0 $X2=7.805
+ $Y2=1
cc_46 N_GND_c_12_p N_A_110_115#_c_441_n 0.00424466f $X=1.985 $Y=0.152 $X2=7.805
+ $Y2=1
cc_47 N_GND_c_47_p N_A_110_115#_c_441_n 0.0070662f $X=2.07 $Y=0.74 $X2=7.805
+ $Y2=1
cc_48 N_GND_c_48_p N_A_110_115#_c_441_n 0.00599718f $X=2.505 $Y=0.152 $X2=7.805
+ $Y2=1
cc_49 N_GND_c_49_p N_A_110_115#_c_441_n 0.012085f $X=2.59 $Y=0.755 $X2=7.805
+ $Y2=1
cc_50 N_GND_c_50_p N_A_110_115#_c_441_n 0.0196453f $X=4.255 $Y=0.152 $X2=7.805
+ $Y2=1
cc_51 N_GND_c_51_p N_A_110_115#_c_441_n 0.00720909f $X=4.34 $Y=0.74 $X2=7.805
+ $Y2=1
cc_52 N_GND_c_52_p N_A_110_115#_c_441_n 0.0196423f $X=6.005 $Y=0.152 $X2=7.805
+ $Y2=1
cc_53 N_GND_c_53_p N_A_110_115#_c_441_n 0.0139942f $X=6.09 $Y=0.755 $X2=7.805
+ $Y2=1
cc_54 N_GND_c_54_p N_A_110_115#_c_441_n 0.0102455f $X=6.955 $Y=0.152 $X2=7.805
+ $Y2=1
cc_55 N_GND_c_55_p N_A_110_115#_c_441_n 0.00848976f $X=7.04 $Y=0.74 $X2=7.805
+ $Y2=1
cc_56 N_GND_c_19_p N_A_110_115#_c_441_n 0.00815276f $X=7.815 $Y=0.152 $X2=7.805
+ $Y2=1
cc_57 N_GND_c_16_p N_A_110_115#_c_441_n 0.00655132f $X=7.9 $Y=0.74 $X2=7.805
+ $Y2=1
cc_58 N_GND_M1018_s N_A_110_115#_c_461_n 0.0017057f $X=1.085 $Y=0.575 $X2=1.305
+ $Y2=1
cc_59 N_GND_M1021_b N_A_110_115#_c_461_n 0.00113133f $X=-0.05 $Y=0 $X2=1.305
+ $Y2=1
cc_60 N_GND_c_4_p N_A_110_115#_c_461_n 0.00660647f $X=1.21 $Y=0.74 $X2=1.305
+ $Y2=1
cc_61 N_GND_c_12_p N_A_110_115#_c_461_n 0.00391005f $X=1.985 $Y=0.152 $X2=1.305
+ $Y2=1
cc_62 N_GND_M1021_b N_A_110_115#_c_465_n 0.00487424f $X=-0.05 $Y=0 $X2=1.22
+ $Y2=1.37
cc_63 N_GND_M1021_b N_A_110_115#_c_466_n 0.00285541f $X=-0.05 $Y=0 $X2=7.89
+ $Y2=1.37
cc_64 N_GND_M1021_b N_A_342_442#_M1005_g 0.087851f $X=-0.05 $Y=0 $X2=1.855
+ $Y2=0.755
cc_65 N_GND_c_12_p N_A_342_442#_M1005_g 0.00606474f $X=1.985 $Y=0.152 $X2=1.855
+ $Y2=0.755
cc_66 N_GND_c_47_p N_A_342_442#_M1005_g 0.00502587f $X=2.07 $Y=0.74 $X2=1.855
+ $Y2=0.755
cc_67 N_GND_c_5_p N_A_342_442#_M1005_g 0.00468827f $X=9.175 $Y=0.19 $X2=1.855
+ $Y2=0.755
cc_68 N_GND_M1021_b N_A_342_442#_c_614_n 0.0245154f $X=-0.05 $Y=0 $X2=1.94
+ $Y2=2.375
cc_69 N_GND_M1021_b N_A_342_442#_c_615_n 0.0182652f $X=-0.05 $Y=0 $X2=2.11
+ $Y2=2.21
cc_70 N_GND_M1021_b N_A_342_442#_c_616_n 0.0217838f $X=-0.05 $Y=0 $X2=3.28
+ $Y2=1.285
cc_71 N_GND_c_49_p N_A_342_442#_c_616_n 0.00673409f $X=2.59 $Y=0.755 $X2=3.28
+ $Y2=1.285
cc_72 N_GND_M1021_b N_A_342_442#_c_618_n 0.00653128f $X=-0.05 $Y=0 $X2=2.2
+ $Y2=1.285
cc_73 N_GND_c_47_p N_A_342_442#_c_618_n 0.00470355f $X=2.07 $Y=0.74 $X2=2.2
+ $Y2=1.285
cc_74 N_GND_M1021_b N_A_342_442#_c_620_n 0.00198494f $X=-0.05 $Y=0 $X2=3.365
+ $Y2=1.2
cc_75 N_GND_M1021_b N_A_342_442#_c_621_n 0.0066411f $X=-0.05 $Y=0 $X2=1.94
+ $Y2=2.375
cc_76 N_GND_M1021_b N_A_342_442#_c_622_n 0.00311983f $X=-0.05 $Y=0 $X2=3.365
+ $Y2=0.755
cc_77 N_GND_c_50_p N_A_342_442#_c_622_n 0.0147897f $X=4.255 $Y=0.152 $X2=3.365
+ $Y2=0.755
cc_78 N_GND_c_5_p N_A_342_442#_c_622_n 0.0098977f $X=9.175 $Y=0.19 $X2=3.365
+ $Y2=0.755
cc_79 N_GND_M1021_b N_D_M1007_g 0.0418787f $X=-0.05 $Y=0 $X2=2.805 $Y2=0.835
cc_80 N_GND_c_49_p N_D_M1007_g 0.00509529f $X=2.59 $Y=0.755 $X2=2.805 $Y2=0.835
cc_81 N_GND_c_50_p N_D_M1007_g 0.00606474f $X=4.255 $Y=0.152 $X2=2.805 $Y2=0.835
cc_82 N_GND_c_5_p N_D_M1007_g 0.00468827f $X=9.175 $Y=0.19 $X2=2.805 $Y2=0.835
cc_83 N_GND_M1021_b N_D_M1028_g 0.0359102f $X=-0.05 $Y=0 $X2=2.805 $Y2=3.235
cc_84 N_GND_M1021_b N_D_c_698_n 0.0324288f $X=-0.05 $Y=0 $X2=2.865 $Y2=1.74
cc_85 N_GND_M1021_b N_D_c_699_n 0.00311208f $X=-0.05 $Y=0 $X2=2.865 $Y2=1.74
cc_86 N_GND_M1021_b D 0.00973922f $X=-0.05 $Y=0 $X2=2.865 $Y2=1.74
cc_87 N_GND_M1021_b N_CK_c_735_n 0.0183851f $X=-0.05 $Y=0 $X2=6.305 $Y2=1.205
cc_88 N_GND_c_53_p N_CK_c_735_n 0.00311745f $X=6.09 $Y=0.755 $X2=6.305 $Y2=1.205
cc_89 N_GND_c_54_p N_CK_c_735_n 0.00606474f $X=6.955 $Y=0.152 $X2=6.305
+ $Y2=1.205
cc_90 N_GND_c_55_p N_CK_c_735_n 0.00359543f $X=7.04 $Y=0.74 $X2=6.305 $Y2=1.205
cc_91 N_GND_c_5_p N_CK_c_735_n 0.00468827f $X=9.175 $Y=0.19 $X2=6.305 $Y2=1.205
cc_92 N_GND_M1021_b N_CK_c_740_n 0.0306664f $X=-0.05 $Y=0 $X2=6.305 $Y2=2.45
cc_93 N_GND_M1021_b N_CK_c_741_n 0.0428261f $X=-0.05 $Y=0 $X2=6.385 $Y2=2.12
cc_94 N_GND_M1021_b N_CK_c_742_n 0.0244095f $X=-0.05 $Y=0 $X2=3.225 $Y2=2.285
cc_95 N_GND_M1021_b N_CK_c_743_n 0.0254608f $X=-0.05 $Y=0 $X2=3.705 $Y2=1.37
cc_96 N_GND_M1021_b N_CK_c_744_n 0.0173906f $X=-0.05 $Y=0 $X2=3.705 $Y2=1.205
cc_97 N_GND_c_50_p N_CK_c_744_n 0.00606474f $X=4.255 $Y=0.152 $X2=3.705
+ $Y2=1.205
cc_98 N_GND_c_5_p N_CK_c_744_n 0.00468827f $X=9.175 $Y=0.19 $X2=3.705 $Y2=1.205
cc_99 N_GND_M1021_b N_CK_c_747_n 0.0267352f $X=-0.05 $Y=0 $X2=4.975 $Y2=1.37
cc_100 N_GND_M1021_b N_CK_c_748_n 0.0174883f $X=-0.05 $Y=0 $X2=4.975 $Y2=1.205
cc_101 N_GND_c_52_p N_CK_c_748_n 0.00606474f $X=6.005 $Y=0.152 $X2=4.975
+ $Y2=1.205
cc_102 N_GND_c_5_p N_CK_c_748_n 0.00468827f $X=9.175 $Y=0.19 $X2=4.975 $Y2=1.205
cc_103 N_GND_M1021_b N_CK_c_751_n 0.022014f $X=-0.05 $Y=0 $X2=5.455 $Y2=2.285
cc_104 N_GND_M1021_b N_CK_c_752_n 0.014732f $X=-0.05 $Y=0 $X2=6.385 $Y2=1.28
cc_105 N_GND_M1021_b N_CK_c_753_n 0.00609317f $X=-0.05 $Y=0 $X2=3.62 $Y2=2.11
cc_106 N_GND_M1021_b N_CK_c_754_n 0.00920685f $X=-0.05 $Y=0 $X2=3.705 $Y2=1.37
cc_107 N_GND_M1021_b N_CK_c_755_n 0.008127f $X=-0.05 $Y=0 $X2=4.975 $Y2=1.37
cc_108 N_GND_M1021_b N_CK_c_756_n 0.00482713f $X=-0.05 $Y=0 $X2=5.37 $Y2=2.11
cc_109 N_GND_M1021_b N_CK_c_757_n 5.00459e-19 $X=-0.05 $Y=0 $X2=5.06 $Y2=2.11
cc_110 N_GND_M1021_b N_CK_c_758_n 6.15269e-19 $X=-0.05 $Y=0 $X2=6.45 $Y2=2.11
cc_111 N_GND_M1021_b N_CK_c_759_n 0.00276905f $X=-0.05 $Y=0 $X2=3.225 $Y2=2.11
cc_112 N_GND_M1021_b N_CK_c_760_n 0.00119864f $X=-0.05 $Y=0 $X2=5.455 $Y2=2.11
cc_113 N_GND_M1021_b N_CK_c_761_n 0.0338168f $X=-0.05 $Y=0 $X2=5.31 $Y2=2.11
cc_114 N_GND_M1021_b N_CK_c_762_n 0.00714094f $X=-0.05 $Y=0 $X2=3.37 $Y2=2.11
cc_115 N_GND_M1021_b N_CK_c_763_n 0.0138229f $X=-0.05 $Y=0 $X2=6.305 $Y2=2.11
cc_116 N_GND_M1021_b N_CK_c_764_n 0.0025628f $X=-0.05 $Y=0 $X2=5.6 $Y2=2.11
cc_117 N_GND_M1021_b CK 0.0016917f $X=-0.05 $Y=0 $X2=6.45 $Y2=2.11
cc_118 N_GND_M1021_b N_A_217_605#_M1027_g 0.0171926f $X=-0.05 $Y=0 $X2=4.125
+ $Y2=0.835
cc_119 N_GND_c_50_p N_A_217_605#_M1027_g 0.00606474f $X=4.255 $Y=0.152 $X2=4.125
+ $Y2=0.835
cc_120 N_GND_c_51_p N_A_217_605#_M1027_g 0.00308284f $X=4.34 $Y=0.74 $X2=4.125
+ $Y2=0.835
cc_121 N_GND_c_5_p N_A_217_605#_M1027_g 0.00468827f $X=9.175 $Y=0.19 $X2=4.125
+ $Y2=0.835
cc_122 N_GND_M1021_b N_A_217_605#_c_990_n 0.0240311f $X=-0.05 $Y=0 $X2=4.48
+ $Y2=1.37
cc_123 N_GND_c_51_p N_A_217_605#_c_990_n 9.93645e-19 $X=4.34 $Y=0.74 $X2=4.48
+ $Y2=1.37
cc_124 N_GND_M1021_b N_A_217_605#_c_992_n 0.0105855f $X=-0.05 $Y=0 $X2=4.2
+ $Y2=1.37
cc_125 N_GND_M1021_b N_A_217_605#_c_993_n 0.0232417f $X=-0.05 $Y=0 $X2=4.48
+ $Y2=2.285
cc_126 N_GND_M1021_b N_A_217_605#_c_994_n 0.0105265f $X=-0.05 $Y=0 $X2=4.2
+ $Y2=2.285
cc_127 N_GND_M1021_b N_A_217_605#_M1025_g 0.0170177f $X=-0.05 $Y=0 $X2=4.555
+ $Y2=0.835
cc_128 N_GND_c_51_p N_A_217_605#_M1025_g 0.00308284f $X=4.34 $Y=0.74 $X2=4.555
+ $Y2=0.835
cc_129 N_GND_c_52_p N_A_217_605#_M1025_g 0.00606474f $X=6.005 $Y=0.152 $X2=4.555
+ $Y2=0.835
cc_130 N_GND_c_5_p N_A_217_605#_M1025_g 0.00468827f $X=9.175 $Y=0.19 $X2=4.555
+ $Y2=0.835
cc_131 N_GND_M1021_b N_A_217_605#_c_999_n 0.011276f $X=-0.05 $Y=0 $X2=1.21
+ $Y2=3.275
cc_132 N_GND_M1021_b N_A_217_605#_c_1000_n 0.0127277f $X=-0.05 $Y=0 $X2=1.555
+ $Y2=1.81
cc_133 N_GND_M1021_b N_A_217_605#_c_1001_n 0.00259716f $X=-0.05 $Y=0 $X2=1.295
+ $Y2=1.81
cc_134 N_GND_M1021_b N_A_217_605#_c_1002_n 0.017579f $X=-0.05 $Y=0 $X2=1.64
+ $Y2=0.74
cc_135 N_GND_c_12_p N_A_217_605#_c_1002_n 0.00734006f $X=1.985 $Y=0.152 $X2=1.64
+ $Y2=0.74
cc_136 N_GND_c_5_p N_A_217_605#_c_1002_n 0.00475776f $X=9.175 $Y=0.19 $X2=1.64
+ $Y2=0.74
cc_137 N_GND_M1021_b N_A_217_605#_c_1005_n 0.00871176f $X=-0.05 $Y=0 $X2=4.295
+ $Y2=2.285
cc_138 N_GND_M1021_b N_A_217_605#_c_1006_n 0.00210386f $X=-0.05 $Y=0 $X2=4.295
+ $Y2=1.37
cc_139 N_GND_c_51_p N_A_217_605#_c_1006_n 0.00441035f $X=4.34 $Y=0.74 $X2=4.295
+ $Y2=1.37
cc_140 N_GND_M1021_b N_A_217_605#_c_1008_n 0.0335787f $X=-0.05 $Y=0 $X2=4.06
+ $Y2=1.37
cc_141 N_GND_M1021_b N_A_217_605#_c_1009_n 0.00340906f $X=-0.05 $Y=0 $X2=1.78
+ $Y2=1.372
cc_142 N_GND_M1021_b N_A_618_89#_c_1124_n 0.0173059f $X=-0.05 $Y=0 $X2=3.165
+ $Y2=1.205
cc_143 N_GND_c_50_p N_A_618_89#_c_1124_n 0.00606474f $X=4.255 $Y=0.152 $X2=3.165
+ $Y2=1.205
cc_144 N_GND_c_5_p N_A_618_89#_c_1124_n 0.00468827f $X=9.175 $Y=0.19 $X2=3.165
+ $Y2=1.205
cc_145 N_GND_M1021_b N_A_618_89#_c_1127_n 0.0203057f $X=-0.05 $Y=0 $X2=3.285
+ $Y2=1.745
cc_146 N_GND_M1021_b N_A_618_89#_c_1128_n 0.0187566f $X=-0.05 $Y=0 $X2=3.69
+ $Y2=1.82
cc_147 N_GND_M1021_b N_A_618_89#_c_1129_n 0.00755029f $X=-0.05 $Y=0 $X2=3.36
+ $Y2=1.82
cc_148 N_GND_M1021_b N_A_618_89#_M1017_g 0.032457f $X=-0.05 $Y=0 $X2=3.765
+ $Y2=3.235
cc_149 N_GND_M1021_b N_A_618_89#_c_1131_n 0.0559794f $X=-0.05 $Y=0 $X2=4.84
+ $Y2=1.82
cc_150 N_GND_M1021_b N_A_618_89#_M1003_g 0.0319667f $X=-0.05 $Y=0 $X2=4.915
+ $Y2=3.235
cc_151 N_GND_M1021_b N_A_618_89#_c_1133_n 0.0187483f $X=-0.05 $Y=0 $X2=5.32
+ $Y2=1.82
cc_152 N_GND_M1021_b N_A_618_89#_M1020_g 0.0322593f $X=-0.05 $Y=0 $X2=5.515
+ $Y2=0.835
cc_153 N_GND_c_52_p N_A_618_89#_M1020_g 0.00606474f $X=6.005 $Y=0.152 $X2=5.515
+ $Y2=0.835
cc_154 N_GND_c_5_p N_A_618_89#_M1020_g 0.00468827f $X=9.175 $Y=0.19 $X2=5.515
+ $Y2=0.835
cc_155 N_GND_M1021_b N_A_618_89#_c_1137_n 0.0141736f $X=-0.05 $Y=0 $X2=3.285
+ $Y2=1.28
cc_156 N_GND_M1021_b N_A_618_89#_c_1138_n 0.00426512f $X=-0.05 $Y=0 $X2=3.765
+ $Y2=1.82
cc_157 N_GND_M1021_b N_A_618_89#_c_1139_n 0.00426512f $X=-0.05 $Y=0 $X2=4.915
+ $Y2=1.82
cc_158 N_GND_M1021_b N_A_618_89#_c_1140_n 0.0333891f $X=-0.05 $Y=0 $X2=5.455
+ $Y2=1.725
cc_159 N_GND_M1021_b N_A_618_89#_c_1141_n 0.00141731f $X=-0.05 $Y=0 $X2=5.455
+ $Y2=1.725
cc_160 N_GND_M1021_b N_A_618_89#_c_1142_n 0.00795998f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=0.755
cc_161 N_GND_c_53_p N_A_618_89#_c_1142_n 4.65312e-19 $X=6.09 $Y=0.755 $X2=6.52
+ $Y2=0.755
cc_162 N_GND_c_54_p N_A_618_89#_c_1142_n 0.00736239f $X=6.955 $Y=0.152 $X2=6.52
+ $Y2=0.755
cc_163 N_GND_c_55_p N_A_618_89#_c_1142_n 0.0140971f $X=7.04 $Y=0.74 $X2=6.52
+ $Y2=0.755
cc_164 N_GND_c_5_p N_A_618_89#_c_1142_n 0.00476261f $X=9.175 $Y=0.19 $X2=6.52
+ $Y2=0.755
cc_165 N_GND_M1021_b N_A_618_89#_c_1147_n 0.012459f $X=-0.05 $Y=0 $X2=6.795
+ $Y2=2.62
cc_166 N_GND_M1021_b N_A_618_89#_c_1148_n 0.0110734f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=1.725
cc_167 N_GND_M1021_b N_A_618_89#_c_1149_n 0.0056826f $X=-0.05 $Y=0 $X2=6.215
+ $Y2=1.74
cc_168 N_GND_M1021_b N_A_618_89#_c_1150_n 0.0019581f $X=-0.05 $Y=0 $X2=6.36
+ $Y2=1.74
cc_169 N_GND_M1021_b N_A_1160_89#_M1009_g 0.00746385f $X=-0.05 $Y=0 $X2=5.875
+ $Y2=3.235
cc_170 N_GND_M1021_b N_A_1160_89#_M1016_g 0.0259924f $X=-0.05 $Y=0 $X2=8.635
+ $Y2=0.755
cc_171 N_GND_c_16_p N_A_1160_89#_M1016_g 0.00359543f $X=7.9 $Y=0.74 $X2=8.635
+ $Y2=0.755
cc_172 N_GND_c_172_p N_A_1160_89#_M1016_g 0.00606474f $X=8.765 $Y=0.152
+ $X2=8.635 $Y2=0.755
cc_173 N_GND_c_173_p N_A_1160_89#_M1016_g 0.00308284f $X=8.85 $Y=0.74 $X2=8.635
+ $Y2=0.755
cc_174 N_GND_c_5_p N_A_1160_89#_M1016_g 0.00468827f $X=9.175 $Y=0.19 $X2=8.635
+ $Y2=0.755
cc_175 N_GND_M1021_b N_A_1160_89#_c_1326_n 0.016106f $X=-0.05 $Y=0 $X2=5.89
+ $Y2=1.205
cc_176 N_GND_c_52_p N_A_1160_89#_c_1326_n 0.00606474f $X=6.005 $Y=0.152 $X2=5.89
+ $Y2=1.205
cc_177 N_GND_c_53_p N_A_1160_89#_c_1326_n 0.00315235f $X=6.09 $Y=0.755 $X2=5.89
+ $Y2=1.205
cc_178 N_GND_c_5_p N_A_1160_89#_c_1326_n 0.00468827f $X=9.175 $Y=0.19 $X2=5.89
+ $Y2=1.205
cc_179 N_GND_M1021_b N_A_1160_89#_c_1330_n 0.00990642f $X=-0.05 $Y=0 $X2=5.89
+ $Y2=1.365
cc_180 N_GND_M1021_b N_A_1160_89#_c_1331_n 0.0116478f $X=-0.05 $Y=0 $X2=5.89
+ $Y2=2.105
cc_181 N_GND_M1021_b N_A_1160_89#_c_1332_n 0.00919812f $X=-0.05 $Y=0 $X2=5.89
+ $Y2=2.255
cc_182 N_GND_M1021_b N_A_1160_89#_c_1333_n 0.0272598f $X=-0.05 $Y=0 $X2=5.965
+ $Y2=1.77
cc_183 N_GND_c_53_p N_A_1160_89#_c_1333_n 0.00110843f $X=6.09 $Y=0.755 $X2=5.965
+ $Y2=1.77
cc_184 N_GND_M1021_b N_A_1160_89#_c_1335_n 0.0119095f $X=-0.05 $Y=0 $X2=5.965
+ $Y2=1.605
cc_185 N_GND_M1021_b N_A_1160_89#_c_1336_n 0.0294757f $X=-0.05 $Y=0 $X2=8.52
+ $Y2=1.74
cc_186 N_GND_M1021_b N_A_1160_89#_c_1337_n 0.0171478f $X=-0.05 $Y=0 $X2=8.522
+ $Y2=1.575
cc_187 N_GND_M1021_b N_A_1160_89#_c_1338_n 0.0136411f $X=-0.05 $Y=0 $X2=8.61
+ $Y2=1.32
cc_188 N_GND_M1021_b N_A_1160_89#_c_1339_n 0.0341464f $X=-0.05 $Y=0 $X2=8.61
+ $Y2=2.375
cc_189 N_GND_M1021_b N_A_1160_89#_c_1340_n 0.00495925f $X=-0.05 $Y=0 $X2=8.61
+ $Y2=2.525
cc_190 N_GND_M1021_b N_A_1160_89#_c_1341_n 0.00212375f $X=-0.05 $Y=0 $X2=5.935
+ $Y2=2.025
cc_191 N_GND_c_53_p N_A_1160_89#_c_1341_n 4.59543e-19 $X=6.09 $Y=0.755 $X2=5.935
+ $Y2=2.025
cc_192 N_GND_M1021_b N_A_1160_89#_c_1343_n 0.00271797f $X=-0.05 $Y=0 $X2=5.935
+ $Y2=2.48
cc_193 N_GND_M1021_b N_A_1160_89#_c_1344_n 0.0119722f $X=-0.05 $Y=0 $X2=7.47
+ $Y2=0.74
cc_194 N_GND_c_19_p N_A_1160_89#_c_1344_n 0.0075556f $X=7.815 $Y=0.152 $X2=7.47
+ $Y2=0.74
cc_195 N_GND_c_5_p N_A_1160_89#_c_1344_n 0.00475776f $X=9.175 $Y=0.19 $X2=7.47
+ $Y2=0.74
cc_196 N_GND_M1021_b N_A_1160_89#_c_1347_n 0.00449369f $X=-0.05 $Y=0 $X2=7.47
+ $Y2=2.96
cc_197 N_GND_M1021_b N_A_1160_89#_c_1348_n 0.0181474f $X=-0.05 $Y=0 $X2=8.52
+ $Y2=1.74
cc_198 N_GND_M1021_b N_A_1160_89#_c_1349_n 0.00134922f $X=-0.05 $Y=0 $X2=7.47
+ $Y2=1.74
cc_199 N_GND_M1021_b N_A_1160_89#_c_1350_n 0.00284861f $X=-0.05 $Y=0 $X2=6.735
+ $Y2=2.48
cc_200 N_GND_M1021_b N_A_1160_89#_c_1351_n 0.0011503f $X=-0.05 $Y=0 $X2=6.08
+ $Y2=2.48
cc_201 N_GND_M1021_b N_A_1160_89#_c_1352_n 0.00577273f $X=-0.05 $Y=0 $X2=6.825
+ $Y2=2.395
cc_202 N_GND_M1021_b N_A_1160_89#_c_1353_n 2.49257e-19 $X=-0.05 $Y=0 $X2=6.915
+ $Y2=1.737
cc_203 N_GND_M1021_b N_A_1160_89#_c_1354_n 0.00280684f $X=-0.05 $Y=0 $X2=8.52
+ $Y2=1.74
cc_204 N_GND_M1021_b N_A_1160_89#_c_1355_n 0.0497022f $X=-0.05 $Y=0 $X2=8.375
+ $Y2=1.74
cc_205 N_GND_M1021_b N_A_998_115#_M1012_g 0.0283844f $X=-0.05 $Y=0 $X2=7.255
+ $Y2=0.755
cc_206 N_GND_c_55_p N_A_998_115#_M1012_g 0.00502587f $X=7.04 $Y=0.74 $X2=7.255
+ $Y2=0.755
cc_207 N_GND_c_19_p N_A_998_115#_M1012_g 0.00606474f $X=7.815 $Y=0.152 $X2=7.255
+ $Y2=0.755
cc_208 N_GND_c_5_p N_A_998_115#_M1012_g 0.00468827f $X=9.175 $Y=0.19 $X2=7.255
+ $Y2=0.755
cc_209 N_GND_M1021_b N_A_998_115#_M1006_g 0.0532683f $X=-0.05 $Y=0 $X2=7.255
+ $Y2=3.445
cc_210 N_GND_M1021_b N_A_998_115#_c_1538_n 0.0362825f $X=-0.05 $Y=0 $X2=7.13
+ $Y2=1.37
cc_211 N_GND_c_55_p N_A_998_115#_c_1538_n 0.00254427f $X=7.04 $Y=0.74 $X2=7.13
+ $Y2=1.37
cc_212 N_GND_M1021_b N_A_998_115#_c_1540_n 0.0113462f $X=-0.05 $Y=0 $X2=4.635
+ $Y2=1.37
cc_213 N_GND_M1021_b N_A_998_115#_c_1541_n 0.00904057f $X=-0.05 $Y=0 $X2=5.315
+ $Y2=1.37
cc_214 N_GND_M1021_b N_A_998_115#_c_1542_n 0.00285975f $X=-0.05 $Y=0 $X2=7.13
+ $Y2=1.37
cc_215 N_GND_c_55_p N_A_998_115#_c_1542_n 0.00241953f $X=7.04 $Y=0.74 $X2=7.13
+ $Y2=1.37
cc_216 N_GND_M1021_b N_A_998_115#_c_1544_n 0.00312748f $X=-0.05 $Y=0 $X2=5.215
+ $Y2=0.755
cc_217 N_GND_c_52_p N_A_998_115#_c_1544_n 0.0150341f $X=6.005 $Y=0.152 $X2=5.215
+ $Y2=0.755
cc_218 N_GND_c_5_p N_A_998_115#_c_1544_n 0.00994746f $X=9.175 $Y=0.19 $X2=5.215
+ $Y2=0.755
cc_219 N_GND_M1021_b N_A_998_115#_c_1547_n 0.00241727f $X=-0.05 $Y=0 $X2=5.18
+ $Y2=1.37
cc_220 N_GND_M1021_b N_A_998_115#_c_1548_n 0.00125111f $X=-0.05 $Y=0 $X2=4.78
+ $Y2=1.37
cc_221 N_GND_M1021_b N_A_998_115#_c_1549_n 0.0136427f $X=-0.05 $Y=0 $X2=6.985
+ $Y2=1.37
cc_222 N_GND_c_53_p N_A_998_115#_c_1549_n 7.83815e-19 $X=6.09 $Y=0.755 $X2=6.985
+ $Y2=1.37
cc_223 N_GND_M1021_b N_A_998_115#_c_1551_n 0.00209768f $X=-0.05 $Y=0 $X2=5.44
+ $Y2=1.37
cc_224 N_GND_M1021_b N_A_998_115#_c_1552_n 6.94251e-19 $X=-0.05 $Y=0 $X2=7.13
+ $Y2=1.37
cc_225 N_GND_M1021_b N_QN_M1008_g 0.0651437f $X=-0.05 $Y=0 $X2=9.065 $Y2=0.755
cc_226 N_GND_c_173_p N_QN_M1008_g 0.00308284f $X=8.85 $Y=0.74 $X2=9.065
+ $Y2=0.755
cc_227 N_GND_c_5_p N_QN_M1008_g 0.00468827f $X=9.175 $Y=0.19 $X2=9.065 $Y2=0.755
cc_228 N_GND_M1021_b N_QN_M1001_g 0.0186095f $X=-0.05 $Y=0 $X2=9.065 $Y2=3.445
cc_229 N_GND_M1021_b N_QN_c_1680_n 0.0291868f $X=-0.05 $Y=0 $X2=9.005 $Y2=1.915
cc_230 N_GND_M1021_b N_QN_c_1681_n 0.00776412f $X=-0.05 $Y=0 $X2=8.42 $Y2=0.74
cc_231 N_GND_c_16_p N_QN_c_1681_n 0.0140971f $X=7.9 $Y=0.74 $X2=8.42 $Y2=0.74
cc_232 N_GND_c_172_p N_QN_c_1681_n 0.00736239f $X=8.765 $Y=0.152 $X2=8.42
+ $Y2=0.74
cc_233 N_GND_c_5_p N_QN_c_1681_n 0.00476261f $X=9.175 $Y=0.19 $X2=8.42 $Y2=0.74
cc_234 N_GND_M1021_b N_QN_c_1685_n 0.00138285f $X=-0.05 $Y=0 $X2=8.42 $Y2=2.48
cc_235 N_GND_M1021_b N_QN_c_1686_n 0.0134367f $X=-0.05 $Y=0 $X2=8.92 $Y2=1.37
cc_236 N_GND_c_173_p N_QN_c_1686_n 0.00779875f $X=8.85 $Y=0.74 $X2=8.92 $Y2=1.37
cc_237 N_GND_M1021_b N_QN_c_1688_n 0.00232247f $X=-0.05 $Y=0 $X2=8.505 $Y2=1.37
cc_238 N_GND_M1021_b N_QN_c_1689_n 0.0138306f $X=-0.05 $Y=0 $X2=8.92 $Y2=2.285
cc_239 N_GND_M1021_b N_QN_c_1690_n 0.00434805f $X=-0.05 $Y=0 $X2=8.505 $Y2=2.285
cc_240 N_GND_M1021_b N_QN_c_1691_n 0.00362324f $X=-0.05 $Y=0 $X2=9.005 $Y2=1.915
cc_241 N_GND_M1021_b QN 0.00270537f $X=-0.05 $Y=0 $X2=8.425 $Y2=2.48
cc_242 N_GND_M1021_b N_Q_c_1771_n 0.0098062f $X=-0.05 $Y=0 $X2=9.28 $Y2=0.74
cc_243 N_GND_c_5_p N_Q_c_1771_n 0.00467398f $X=9.175 $Y=0.19 $X2=9.28 $Y2=0.74
cc_244 N_GND_M1021_b N_Q_c_1773_n 0.0625704f $X=-0.05 $Y=0 $X2=9.395 $Y2=2.68
cc_245 N_GND_M1021_b N_Q_c_1774_n 0.0189963f $X=-0.05 $Y=0 $X2=9.395 $Y2=1.035
cc_246 N_VDD_M1004_b N_RN_M1004_g 0.0266406f $X=-0.05 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_247 N_VDD_c_247_p N_RN_M1004_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_248 N_VDD_c_248_p N_RN_M1004_g 0.00606474f $X=1.915 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_249 N_VDD_c_249_p N_RN_M1004_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.475
+ $Y2=3.235
cc_250 N_VDD_M1004_s N_RN_c_382_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32
+ $Y2=2.85
cc_251 N_VDD_M1004_b N_RN_c_382_n 0.00618364f $X=-0.05 $Y=2.425 $X2=0.32
+ $Y2=2.85
cc_252 N_VDD_c_247_p N_RN_c_382_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_253 N_VDD_M1004_s RN 0.016276f $X=0.135 $Y=2.605 $X2=0.325 $Y2=2.85
cc_254 N_VDD_c_247_p RN 0.00522047f $X=0.26 $Y=3.635 $X2=0.325 $Y2=2.85
cc_255 N_VDD_M1004_b N_A_110_115#_M1015_g 0.0463013f $X=-0.05 $Y=2.425 $X2=1.425
+ $Y2=3.445
cc_256 N_VDD_c_248_p N_A_110_115#_M1015_g 0.00606474f $X=1.915 $Y=4.287
+ $X2=1.425 $Y2=3.445
cc_257 N_VDD_c_249_p N_A_110_115#_M1015_g 0.00468827f $X=9.175 $Y=4.25 $X2=1.425
+ $Y2=3.445
cc_258 N_VDD_M1004_b N_A_110_115#_M1030_g 0.0450837f $X=-0.05 $Y=2.425 $X2=7.615
+ $Y2=3.445
cc_259 N_VDD_c_259_p N_A_110_115#_M1030_g 0.00606474f $X=7.745 $Y=4.287
+ $X2=7.615 $Y2=3.445
cc_260 N_VDD_c_260_p N_A_110_115#_M1030_g 0.00713292f $X=7.83 $Y=3.275 $X2=7.615
+ $Y2=3.445
cc_261 N_VDD_c_249_p N_A_110_115#_M1030_g 0.00468827f $X=9.175 $Y=4.25 $X2=7.615
+ $Y2=3.445
cc_262 N_VDD_M1004_b N_A_110_115#_c_431_n 0.00549797f $X=-0.05 $Y=2.425 $X2=0.69
+ $Y2=2.95
cc_263 N_VDD_c_248_p N_A_110_115#_c_431_n 0.00757793f $X=1.915 $Y=4.287 $X2=0.69
+ $Y2=2.95
cc_264 N_VDD_c_249_p N_A_110_115#_c_431_n 0.00476261f $X=9.175 $Y=4.25 $X2=0.69
+ $Y2=2.95
cc_265 N_VDD_M1004_b N_A_342_442#_M1002_g 0.0430317f $X=-0.05 $Y=2.425 $X2=1.785
+ $Y2=3.445
cc_266 N_VDD_c_248_p N_A_342_442#_M1002_g 0.00606474f $X=1.915 $Y=4.287
+ $X2=1.785 $Y2=3.445
cc_267 N_VDD_c_267_p N_A_342_442#_M1002_g 0.00713292f $X=2 $Y=3.275 $X2=1.785
+ $Y2=3.445
cc_268 N_VDD_c_249_p N_A_342_442#_M1002_g 0.00468827f $X=9.175 $Y=4.25 $X2=1.785
+ $Y2=3.445
cc_269 N_VDD_M1004_b N_A_342_442#_c_614_n 0.015181f $X=-0.05 $Y=2.425 $X2=1.94
+ $Y2=2.375
cc_270 N_VDD_c_267_p N_A_342_442#_c_614_n 9.61776e-19 $X=2 $Y=3.275 $X2=1.94
+ $Y2=2.375
cc_271 N_VDD_M1028_s N_A_342_442#_c_631_n 0.0125004f $X=2.465 $Y=2.605 $X2=3.295
+ $Y2=2.705
cc_272 N_VDD_M1004_b N_A_342_442#_c_631_n 0.0199377f $X=-0.05 $Y=2.425 $X2=3.295
+ $Y2=2.705
cc_273 N_VDD_c_273_p N_A_342_442#_c_631_n 0.00952036f $X=2.59 $Y=3.295 $X2=3.295
+ $Y2=2.705
cc_274 N_VDD_M1004_b N_A_342_442#_c_634_n 0.00313975f $X=-0.05 $Y=2.425
+ $X2=3.465 $Y2=2.955
cc_275 N_VDD_c_275_p N_A_342_442#_c_634_n 0.0151129f $X=4.255 $Y=4.287 $X2=3.465
+ $Y2=2.955
cc_276 N_VDD_c_249_p N_A_342_442#_c_634_n 0.00958198f $X=9.175 $Y=4.25 $X2=3.465
+ $Y2=2.955
cc_277 N_VDD_M1004_b N_A_342_442#_c_621_n 0.0146567f $X=-0.05 $Y=2.425 $X2=1.94
+ $Y2=2.375
cc_278 N_VDD_c_267_p N_A_342_442#_c_621_n 0.00826787f $X=2 $Y=3.275 $X2=1.94
+ $Y2=2.375
cc_279 N_VDD_M1004_b N_D_M1028_g 0.0219788f $X=-0.05 $Y=2.425 $X2=2.805
+ $Y2=3.235
cc_280 N_VDD_c_267_p N_D_M1028_g 0.00284049f $X=2 $Y=3.275 $X2=2.805 $Y2=3.235
cc_281 N_VDD_c_273_p N_D_M1028_g 0.00636672f $X=2.59 $Y=3.295 $X2=2.805
+ $Y2=3.235
cc_282 N_VDD_c_275_p N_D_M1028_g 0.00606474f $X=4.255 $Y=4.287 $X2=2.805
+ $Y2=3.235
cc_283 N_VDD_c_249_p N_D_M1028_g 0.00468827f $X=9.175 $Y=4.25 $X2=2.805
+ $Y2=3.235
cc_284 N_VDD_M1004_b N_CK_M1024_g 0.020128f $X=-0.05 $Y=2.425 $X2=3.165
+ $Y2=3.235
cc_285 N_VDD_c_275_p N_CK_M1024_g 0.00606474f $X=4.255 $Y=4.287 $X2=3.165
+ $Y2=3.235
cc_286 N_VDD_c_249_p N_CK_M1024_g 0.00468827f $X=9.175 $Y=4.25 $X2=3.165
+ $Y2=3.235
cc_287 N_VDD_M1004_b N_CK_M1000_g 0.0201163f $X=-0.05 $Y=2.425 $X2=5.515
+ $Y2=3.235
cc_288 N_VDD_c_288_p N_CK_M1000_g 0.00606474f $X=6.005 $Y=4.287 $X2=5.515
+ $Y2=3.235
cc_289 N_VDD_c_249_p N_CK_M1000_g 0.00468827f $X=9.175 $Y=4.25 $X2=5.515
+ $Y2=3.235
cc_290 N_VDD_M1004_b N_CK_c_740_n 0.00796681f $X=-0.05 $Y=2.425 $X2=6.305
+ $Y2=2.45
cc_291 N_VDD_M1004_b N_CK_M1029_g 0.0241399f $X=-0.05 $Y=2.425 $X2=6.305
+ $Y2=3.235
cc_292 N_VDD_c_292_p N_CK_M1029_g 0.00409291f $X=6.09 $Y=3.21 $X2=6.305
+ $Y2=3.235
cc_293 N_VDD_c_259_p N_CK_M1029_g 0.00606474f $X=7.745 $Y=4.287 $X2=6.305
+ $Y2=3.235
cc_294 N_VDD_c_249_p N_CK_M1029_g 0.00468827f $X=9.175 $Y=4.25 $X2=6.305
+ $Y2=3.235
cc_295 N_VDD_M1004_b N_CK_c_742_n 0.00487135f $X=-0.05 $Y=2.425 $X2=3.225
+ $Y2=2.285
cc_296 N_VDD_M1004_b N_CK_c_751_n 0.00486793f $X=-0.05 $Y=2.425 $X2=5.455
+ $Y2=2.285
cc_297 N_VDD_M1004_b N_CK_c_758_n 0.0010436f $X=-0.05 $Y=2.425 $X2=6.45 $Y2=2.11
cc_298 N_VDD_M1004_b N_CK_c_759_n 6.42499e-19 $X=-0.05 $Y=2.425 $X2=3.225
+ $Y2=2.11
cc_299 N_VDD_M1004_b N_CK_c_760_n 0.0022456f $X=-0.05 $Y=2.425 $X2=5.455
+ $Y2=2.11
cc_300 N_VDD_M1004_b N_A_217_605#_M1022_g 0.0192219f $X=-0.05 $Y=2.425 $X2=4.125
+ $Y2=3.235
cc_301 N_VDD_c_275_p N_A_217_605#_M1022_g 0.00606474f $X=4.255 $Y=4.287
+ $X2=4.125 $Y2=3.235
cc_302 N_VDD_c_302_p N_A_217_605#_M1022_g 0.00337744f $X=4.34 $Y=3.295 $X2=4.125
+ $Y2=3.235
cc_303 N_VDD_c_249_p N_A_217_605#_M1022_g 0.00468827f $X=9.175 $Y=4.25 $X2=4.125
+ $Y2=3.235
cc_304 N_VDD_c_302_p N_A_217_605#_c_993_n 8.24975e-19 $X=4.34 $Y=3.295 $X2=4.48
+ $Y2=2.285
cc_305 N_VDD_M1004_b N_A_217_605#_M1014_g 0.0181098f $X=-0.05 $Y=2.425 $X2=4.555
+ $Y2=3.235
cc_306 N_VDD_c_302_p N_A_217_605#_M1014_g 0.00337744f $X=4.34 $Y=3.295 $X2=4.555
+ $Y2=3.235
cc_307 N_VDD_c_288_p N_A_217_605#_M1014_g 0.00606474f $X=6.005 $Y=4.287
+ $X2=4.555 $Y2=3.235
cc_308 N_VDD_c_249_p N_A_217_605#_M1014_g 0.00468827f $X=9.175 $Y=4.25 $X2=4.555
+ $Y2=3.235
cc_309 N_VDD_M1004_b N_A_217_605#_c_999_n 0.0163203f $X=-0.05 $Y=2.425 $X2=1.21
+ $Y2=3.275
cc_310 N_VDD_c_248_p N_A_217_605#_c_999_n 0.00745733f $X=1.915 $Y=4.287 $X2=1.21
+ $Y2=3.275
cc_311 N_VDD_c_249_p N_A_217_605#_c_999_n 0.00476261f $X=9.175 $Y=4.25 $X2=1.21
+ $Y2=3.275
cc_312 N_VDD_M1004_b N_A_217_605#_c_1005_n 0.00424346f $X=-0.05 $Y=2.425
+ $X2=4.295 $Y2=2.285
cc_313 N_VDD_c_302_p N_A_217_605#_c_1005_n 0.004428f $X=4.34 $Y=3.295 $X2=4.295
+ $Y2=2.285
cc_314 N_VDD_M1004_b N_A_618_89#_M1017_g 0.0215131f $X=-0.05 $Y=2.425 $X2=3.765
+ $Y2=3.235
cc_315 N_VDD_c_275_p N_A_618_89#_M1017_g 0.00606474f $X=4.255 $Y=4.287 $X2=3.765
+ $Y2=3.235
cc_316 N_VDD_c_249_p N_A_618_89#_M1017_g 0.00468827f $X=9.175 $Y=4.25 $X2=3.765
+ $Y2=3.235
cc_317 N_VDD_M1004_b N_A_618_89#_M1003_g 0.0214821f $X=-0.05 $Y=2.425 $X2=4.915
+ $Y2=3.235
cc_318 N_VDD_c_288_p N_A_618_89#_M1003_g 0.00606474f $X=6.005 $Y=4.287 $X2=4.915
+ $Y2=3.235
cc_319 N_VDD_c_249_p N_A_618_89#_M1003_g 0.00468827f $X=9.175 $Y=4.25 $X2=4.915
+ $Y2=3.235
cc_320 N_VDD_M1004_b N_A_618_89#_c_1157_n 0.00156053f $X=-0.05 $Y=2.425 $X2=6.52
+ $Y2=2.955
cc_321 N_VDD_c_259_p N_A_618_89#_c_1157_n 0.00736239f $X=7.745 $Y=4.287 $X2=6.52
+ $Y2=2.955
cc_322 N_VDD_c_249_p N_A_618_89#_c_1157_n 0.00476261f $X=9.175 $Y=4.25 $X2=6.52
+ $Y2=2.955
cc_323 N_VDD_M1004_b N_A_618_89#_c_1147_n 0.00552543f $X=-0.05 $Y=2.425
+ $X2=6.795 $Y2=2.62
cc_324 N_VDD_M1004_b N_A_618_89#_c_1161_n 0.0123356f $X=-0.05 $Y=2.425 $X2=6.795
+ $Y2=2.705
cc_325 N_VDD_M1004_b N_A_1160_89#_M1009_g 0.0178558f $X=-0.05 $Y=2.425 $X2=5.875
+ $Y2=3.235
cc_326 N_VDD_c_288_p N_A_1160_89#_M1009_g 0.00606474f $X=6.005 $Y=4.287
+ $X2=5.875 $Y2=3.235
cc_327 N_VDD_c_292_p N_A_1160_89#_M1009_g 0.00409291f $X=6.09 $Y=3.21 $X2=5.875
+ $Y2=3.235
cc_328 N_VDD_c_249_p N_A_1160_89#_M1009_g 0.00468827f $X=9.175 $Y=4.25 $X2=5.875
+ $Y2=3.235
cc_329 N_VDD_M1004_b N_A_1160_89#_M1011_g 0.0412931f $X=-0.05 $Y=2.425 $X2=8.635
+ $Y2=3.445
cc_330 N_VDD_c_260_p N_A_1160_89#_M1011_g 0.00453298f $X=7.83 $Y=3.275 $X2=8.635
+ $Y2=3.445
cc_331 N_VDD_c_331_p N_A_1160_89#_M1011_g 0.00606474f $X=8.765 $Y=4.287
+ $X2=8.635 $Y2=3.445
cc_332 N_VDD_c_332_p N_A_1160_89#_M1011_g 0.00602599f $X=8.85 $Y=3.265 $X2=8.635
+ $Y2=3.445
cc_333 N_VDD_c_249_p N_A_1160_89#_M1011_g 0.00468827f $X=9.175 $Y=4.25 $X2=8.635
+ $Y2=3.445
cc_334 N_VDD_M1004_b N_A_1160_89#_c_1340_n 0.00913729f $X=-0.05 $Y=2.425
+ $X2=8.61 $Y2=2.525
cc_335 N_VDD_M1004_b N_A_1160_89#_c_1343_n 0.00242843f $X=-0.05 $Y=2.425
+ $X2=5.935 $Y2=2.48
cc_336 N_VDD_c_292_p N_A_1160_89#_c_1343_n 4.62798e-19 $X=6.09 $Y=3.21 $X2=5.935
+ $Y2=2.48
cc_337 N_VDD_M1004_b N_A_1160_89#_c_1368_n 0.00156053f $X=-0.05 $Y=2.425
+ $X2=7.04 $Y2=3.275
cc_338 N_VDD_c_259_p N_A_1160_89#_c_1368_n 0.00736239f $X=7.745 $Y=4.287
+ $X2=7.04 $Y2=3.275
cc_339 N_VDD_c_249_p N_A_1160_89#_c_1368_n 0.00476261f $X=9.175 $Y=4.25 $X2=7.04
+ $Y2=3.275
cc_340 N_VDD_M1004_b N_A_1160_89#_c_1371_n 0.00371018f $X=-0.05 $Y=2.425
+ $X2=7.385 $Y2=3.045
cc_341 N_VDD_M1004_b N_A_1160_89#_c_1372_n 0.00767127f $X=-0.05 $Y=2.425
+ $X2=7.125 $Y2=3.045
cc_342 N_VDD_M1004_b N_A_1160_89#_c_1347_n 0.00448797f $X=-0.05 $Y=2.425
+ $X2=7.47 $Y2=2.96
cc_343 N_VDD_M1004_b N_A_1160_89#_c_1350_n 0.00938985f $X=-0.05 $Y=2.425
+ $X2=6.735 $Y2=2.48
cc_344 N_VDD_c_292_p N_A_1160_89#_c_1350_n 0.00425473f $X=6.09 $Y=3.21 $X2=6.735
+ $Y2=2.48
cc_345 N_VDD_M1004_b N_A_1160_89#_c_1351_n 0.00604093f $X=-0.05 $Y=2.425
+ $X2=6.08 $Y2=2.48
cc_346 N_VDD_c_292_p N_A_1160_89#_c_1351_n 0.003295f $X=6.09 $Y=3.21 $X2=6.08
+ $Y2=2.48
cc_347 N_VDD_M1004_b N_A_998_115#_M1006_g 0.0487838f $X=-0.05 $Y=2.425 $X2=7.255
+ $Y2=3.445
cc_348 N_VDD_c_259_p N_A_998_115#_M1006_g 0.00606474f $X=7.745 $Y=4.287
+ $X2=7.255 $Y2=3.445
cc_349 N_VDD_c_249_p N_A_998_115#_M1006_g 0.00468827f $X=9.175 $Y=4.25 $X2=7.255
+ $Y2=3.445
cc_350 N_VDD_M1004_b N_A_998_115#_c_1540_n 0.00168314f $X=-0.05 $Y=2.425
+ $X2=4.635 $Y2=1.37
cc_351 N_VDD_M1004_b N_A_998_115#_c_1557_n 0.00313975f $X=-0.05 $Y=2.425
+ $X2=5.215 $Y2=3.295
cc_352 N_VDD_c_288_p N_A_998_115#_c_1557_n 0.0149205f $X=6.005 $Y=4.287
+ $X2=5.215 $Y2=3.295
cc_353 N_VDD_c_249_p N_A_998_115#_c_1557_n 0.00958198f $X=9.175 $Y=4.25
+ $X2=5.215 $Y2=3.295
cc_354 N_VDD_M1004_b N_QN_M1001_g 0.051339f $X=-0.05 $Y=2.425 $X2=9.065
+ $Y2=3.445
cc_355 N_VDD_c_332_p N_QN_M1001_g 0.00601131f $X=8.85 $Y=3.265 $X2=9.065
+ $Y2=3.445
cc_356 N_VDD_c_356_p N_QN_M1001_g 0.00606474f $X=9.175 $Y=4.22 $X2=9.065
+ $Y2=3.445
cc_357 N_VDD_c_249_p N_QN_M1001_g 0.00468827f $X=9.175 $Y=4.25 $X2=9.065
+ $Y2=3.445
cc_358 N_VDD_c_332_p N_QN_c_1680_n 2.00737e-19 $X=8.85 $Y=3.265 $X2=9.005
+ $Y2=1.915
cc_359 N_VDD_M1004_b N_QN_c_1685_n 0.0181975f $X=-0.05 $Y=2.425 $X2=8.42
+ $Y2=2.48
cc_360 N_VDD_c_260_p N_QN_c_1685_n 0.0313352f $X=7.83 $Y=3.275 $X2=8.42 $Y2=2.48
cc_361 N_VDD_c_331_p N_QN_c_1685_n 0.00736239f $X=8.765 $Y=4.287 $X2=8.42
+ $Y2=2.48
cc_362 N_VDD_c_332_p N_QN_c_1685_n 0.0159141f $X=8.85 $Y=3.265 $X2=8.42 $Y2=2.48
cc_363 N_VDD_c_249_p N_QN_c_1685_n 0.00476261f $X=9.175 $Y=4.25 $X2=8.42
+ $Y2=2.48
cc_364 N_VDD_c_332_p N_QN_c_1689_n 0.00856258f $X=8.85 $Y=3.265 $X2=8.92
+ $Y2=2.285
cc_365 N_VDD_M1004_b QN 0.0110801f $X=-0.05 $Y=2.425 $X2=8.425 $Y2=2.48
cc_366 N_VDD_M1004_b N_Q_c_1775_n 0.00508086f $X=-0.05 $Y=2.425 $X2=9.28
+ $Y2=3.265
cc_367 N_VDD_c_332_p N_Q_c_1775_n 0.00454099f $X=8.85 $Y=3.265 $X2=9.28
+ $Y2=3.265
cc_368 N_VDD_c_356_p N_Q_c_1775_n 0.00736239f $X=9.175 $Y=4.22 $X2=9.28
+ $Y2=3.265
cc_369 N_VDD_c_249_p N_Q_c_1775_n 0.00476261f $X=9.175 $Y=4.25 $X2=9.28
+ $Y2=3.265
cc_370 N_VDD_M1004_b N_Q_c_1773_n 0.0127419f $X=-0.05 $Y=2.425 $X2=9.395
+ $Y2=2.68
cc_371 N_VDD_M1004_b N_Q_c_1780_n 0.0190821f $X=-0.05 $Y=2.425 $X2=9.28
+ $Y2=2.807
cc_372 N_VDD_c_332_p N_Q_c_1780_n 0.00905719f $X=8.85 $Y=3.265 $X2=9.28
+ $Y2=2.807
cc_373 N_VDD_M1004_b Q 0.0106945f $X=-0.05 $Y=2.425 $X2=9.275 $Y2=2.85
cc_374 N_VDD_c_332_p Q 0.00675808f $X=8.85 $Y=3.265 $X2=9.275 $Y2=2.85
cc_375 RN N_A_110_115#_M1004_d 0.00410657f $X=0.325 $Y=2.85 $X2=0.55 $Y2=2.605
cc_376 N_RN_c_380_n N_A_110_115#_M1015_g 0.00315143f $X=0.475 $Y=1.99 $X2=1.425
+ $Y2=3.445
cc_377 N_RN_M1021_g N_A_110_115#_c_425_n 0.00524963f $X=0.475 $Y=0.835 $X2=1.425
+ $Y2=1.21
cc_378 N_RN_M1004_g N_A_110_115#_c_431_n 0.00968001f $X=0.475 $Y=3.235 $X2=0.69
+ $Y2=2.95
cc_379 N_RN_c_382_n N_A_110_115#_c_431_n 0.0281933f $X=0.32 $Y=2.85 $X2=0.69
+ $Y2=2.95
cc_380 RN N_A_110_115#_c_431_n 0.0097626f $X=0.325 $Y=2.85 $X2=0.69 $Y2=2.95
cc_381 N_RN_M1021_g N_A_110_115#_c_432_n 0.0107733f $X=0.475 $Y=0.835 $X2=0.87
+ $Y2=2.175
cc_382 N_RN_c_380_n N_A_110_115#_c_432_n 0.00370757f $X=0.475 $Y=1.99 $X2=0.87
+ $Y2=2.175
cc_383 N_RN_M1004_g N_A_110_115#_c_432_n 0.00363549f $X=0.475 $Y=3.235 $X2=0.87
+ $Y2=2.175
cc_384 N_RN_c_382_n N_A_110_115#_c_432_n 0.0072511f $X=0.32 $Y=2.85 $X2=0.87
+ $Y2=2.175
cc_385 N_RN_c_383_n N_A_110_115#_c_432_n 0.0248372f $X=0.32 $Y=1.825 $X2=0.87
+ $Y2=2.175
cc_386 N_RN_M1021_g N_A_110_115#_c_435_n 0.0067448f $X=0.475 $Y=0.835 $X2=0.955
+ $Y2=1.21
cc_387 N_RN_c_380_n N_A_110_115#_c_435_n 0.00166615f $X=0.475 $Y=1.99 $X2=0.955
+ $Y2=1.21
cc_388 N_RN_c_383_n N_A_110_115#_c_435_n 3.95917e-19 $X=0.32 $Y=1.825 $X2=0.955
+ $Y2=1.21
cc_389 N_RN_c_380_n N_A_110_115#_c_436_n 0.00191737f $X=0.475 $Y=1.99 $X2=0.87
+ $Y2=2.26
cc_390 N_RN_M1004_g N_A_110_115#_c_436_n 0.00385986f $X=0.475 $Y=3.235 $X2=0.87
+ $Y2=2.26
cc_391 N_RN_c_382_n N_A_110_115#_c_436_n 0.0113366f $X=0.32 $Y=2.85 $X2=0.87
+ $Y2=2.26
cc_392 N_RN_c_383_n N_A_110_115#_c_436_n 7.08415e-19 $X=0.32 $Y=1.825 $X2=0.87
+ $Y2=2.26
cc_393 N_RN_M1004_g N_A_217_605#_c_999_n 0.0035258f $X=0.475 $Y=3.235 $X2=1.21
+ $Y2=3.275
cc_394 RN N_A_217_605#_c_999_n 8.83853e-19 $X=0.325 $Y=2.85 $X2=1.21 $Y2=3.275
cc_395 N_A_110_115#_c_441_n N_A_342_442#_M1031_d 0.0032387f $X=7.805 $Y=1
+ $X2=3.24 $Y2=0.575
cc_396 N_A_110_115#_c_413_n N_A_342_442#_M1005_g 0.0597799f $X=1.425 $Y=1.045
+ $X2=1.855 $Y2=0.755
cc_397 N_A_110_115#_c_441_n N_A_342_442#_M1005_g 0.00770937f $X=7.805 $Y=1
+ $X2=1.855 $Y2=0.755
cc_398 N_A_110_115#_M1015_g N_A_342_442#_c_614_n 0.106726f $X=1.425 $Y=3.445
+ $X2=1.94 $Y2=2.375
cc_399 N_A_110_115#_c_441_n N_A_342_442#_c_616_n 0.0257941f $X=7.805 $Y=1
+ $X2=3.28 $Y2=1.285
cc_400 N_A_110_115#_c_441_n N_A_342_442#_c_618_n 0.00300956f $X=7.805 $Y=1
+ $X2=2.2 $Y2=1.285
cc_401 N_A_110_115#_c_441_n N_A_342_442#_c_620_n 0.0151351f $X=7.805 $Y=1
+ $X2=3.365 $Y2=1.2
cc_402 N_A_110_115#_M1015_g N_A_342_442#_c_621_n 9.08764e-19 $X=1.425 $Y=3.445
+ $X2=1.94 $Y2=2.375
cc_403 N_A_110_115#_c_441_n N_A_342_442#_c_622_n 0.0133869f $X=7.805 $Y=1
+ $X2=3.365 $Y2=0.755
cc_404 N_A_110_115#_c_441_n N_D_M1007_g 0.00683925f $X=7.805 $Y=1 $X2=2.805
+ $Y2=0.835
cc_405 N_A_110_115#_c_441_n N_CK_c_735_n 0.00692639f $X=7.805 $Y=1 $X2=6.305
+ $Y2=1.205
cc_406 N_A_110_115#_c_441_n N_CK_c_743_n 8.06574e-19 $X=7.805 $Y=1 $X2=3.705
+ $Y2=1.37
cc_407 N_A_110_115#_c_441_n N_CK_c_744_n 0.0064255f $X=7.805 $Y=1 $X2=3.705
+ $Y2=1.205
cc_408 N_A_110_115#_c_441_n N_CK_c_747_n 8.06574e-19 $X=7.805 $Y=1 $X2=4.975
+ $Y2=1.37
cc_409 N_A_110_115#_c_441_n N_CK_c_748_n 0.00633231f $X=7.805 $Y=1 $X2=4.975
+ $Y2=1.205
cc_410 N_A_110_115#_c_441_n N_CK_c_752_n 0.00109675f $X=7.805 $Y=1 $X2=6.385
+ $Y2=1.28
cc_411 N_A_110_115#_c_441_n N_CK_c_754_n 0.00493929f $X=7.805 $Y=1 $X2=3.705
+ $Y2=1.37
cc_412 N_A_110_115#_c_441_n N_CK_c_755_n 0.00493657f $X=7.805 $Y=1 $X2=4.975
+ $Y2=1.37
cc_413 N_A_110_115#_c_441_n N_A_217_605#_M1018_d 0.00142852f $X=7.805 $Y=1
+ $X2=1.5 $Y2=0.575
cc_414 N_A_110_115#_c_441_n N_A_217_605#_M1027_g 0.00607163f $X=7.805 $Y=1
+ $X2=4.125 $Y2=0.835
cc_415 N_A_110_115#_c_441_n N_A_217_605#_c_990_n 2.42482e-19 $X=7.805 $Y=1
+ $X2=4.48 $Y2=1.37
cc_416 N_A_110_115#_c_441_n N_A_217_605#_M1025_g 0.00632589f $X=7.805 $Y=1
+ $X2=4.555 $Y2=0.835
cc_417 N_A_110_115#_M1015_g N_A_217_605#_c_999_n 0.0409873f $X=1.425 $Y=3.445
+ $X2=1.21 $Y2=3.275
cc_418 N_A_110_115#_c_431_n N_A_217_605#_c_999_n 0.0652498f $X=0.69 $Y=2.95
+ $X2=1.21 $Y2=3.275
cc_419 N_A_110_115#_c_432_n N_A_217_605#_c_999_n 0.0210459f $X=0.87 $Y=2.175
+ $X2=1.21 $Y2=3.275
cc_420 N_A_110_115#_c_436_n N_A_217_605#_c_999_n 0.0134441f $X=0.87 $Y=2.26
+ $X2=1.21 $Y2=3.275
cc_421 N_A_110_115#_M1015_g N_A_217_605#_c_1000_n 0.0188678f $X=1.425 $Y=3.445
+ $X2=1.555 $Y2=1.81
cc_422 N_A_110_115#_c_425_n N_A_217_605#_c_1000_n 6.98912e-19 $X=1.425 $Y=1.21
+ $X2=1.555 $Y2=1.81
cc_423 N_A_110_115#_c_437_n N_A_217_605#_c_1000_n 0.00235169f $X=1.22 $Y=1.21
+ $X2=1.555 $Y2=1.81
cc_424 N_A_110_115#_c_465_n N_A_217_605#_c_1000_n 0.00181457f $X=1.22 $Y=1.37
+ $X2=1.555 $Y2=1.81
cc_425 N_A_110_115#_c_425_n N_A_217_605#_c_1001_n 0.00117358f $X=1.425 $Y=1.21
+ $X2=1.295 $Y2=1.81
cc_426 N_A_110_115#_c_432_n N_A_217_605#_c_1001_n 0.0142099f $X=0.87 $Y=2.175
+ $X2=1.295 $Y2=1.81
cc_427 N_A_110_115#_c_433_n N_A_217_605#_c_1001_n 2.13728e-19 $X=1.135 $Y=1.21
+ $X2=1.295 $Y2=1.81
cc_428 N_A_110_115#_c_437_n N_A_217_605#_c_1001_n 0.00732624f $X=1.22 $Y=1.21
+ $X2=1.295 $Y2=1.81
cc_429 N_A_110_115#_c_465_n N_A_217_605#_c_1001_n 0.00574122f $X=1.22 $Y=1.37
+ $X2=1.295 $Y2=1.81
cc_430 N_A_110_115#_c_413_n N_A_217_605#_c_1002_n 0.00886891f $X=1.425 $Y=1.045
+ $X2=1.64 $Y2=0.74
cc_431 N_A_110_115#_c_432_n N_A_217_605#_c_1002_n 0.00730421f $X=0.87 $Y=2.175
+ $X2=1.64 $Y2=0.74
cc_432 N_A_110_115#_c_435_n N_A_217_605#_c_1002_n 0.00143173f $X=0.955 $Y=1.21
+ $X2=1.64 $Y2=0.74
cc_433 N_A_110_115#_c_437_n N_A_217_605#_c_1002_n 0.0197974f $X=1.22 $Y=1.21
+ $X2=1.64 $Y2=0.74
cc_434 N_A_110_115#_c_534_p N_A_217_605#_c_1002_n 0.00177859f $X=1.22 $Y=1.255
+ $X2=1.64 $Y2=0.74
cc_435 N_A_110_115#_c_441_n N_A_217_605#_c_1002_n 0.0195703f $X=7.805 $Y=1
+ $X2=1.64 $Y2=0.74
cc_436 N_A_110_115#_c_465_n N_A_217_605#_c_1002_n 0.00122345f $X=1.22 $Y=1.37
+ $X2=1.64 $Y2=0.74
cc_437 N_A_110_115#_c_441_n N_A_217_605#_c_1006_n 0.00476535f $X=7.805 $Y=1
+ $X2=4.295 $Y2=1.37
cc_438 N_A_110_115#_c_441_n N_A_217_605#_c_1008_n 0.184203f $X=7.805 $Y=1
+ $X2=4.06 $Y2=1.37
cc_439 N_A_110_115#_M1015_g N_A_217_605#_c_1009_n 0.00152013f $X=1.425 $Y=3.445
+ $X2=1.78 $Y2=1.372
cc_440 N_A_110_115#_c_425_n N_A_217_605#_c_1009_n 0.0015251f $X=1.425 $Y=1.21
+ $X2=1.78 $Y2=1.372
cc_441 N_A_110_115#_c_437_n N_A_217_605#_c_1009_n 9.3821e-19 $X=1.22 $Y=1.21
+ $X2=1.78 $Y2=1.372
cc_442 N_A_110_115#_c_534_p N_A_217_605#_c_1009_n 3.8078e-19 $X=1.22 $Y=1.255
+ $X2=1.78 $Y2=1.372
cc_443 N_A_110_115#_c_441_n N_A_217_605#_c_1009_n 0.0254104f $X=7.805 $Y=1
+ $X2=1.78 $Y2=1.372
cc_444 N_A_110_115#_c_465_n N_A_217_605#_c_1009_n 0.0252399f $X=1.22 $Y=1.37
+ $X2=1.78 $Y2=1.372
cc_445 N_A_110_115#_c_441_n N_A_217_605#_c_1058_n 0.0259207f $X=7.805 $Y=1
+ $X2=4.205 $Y2=1.37
cc_446 N_A_110_115#_c_441_n N_A_618_89#_M1010_d 0.00188999f $X=7.805 $Y=1
+ $X2=6.38 $Y2=0.575
cc_447 N_A_110_115#_c_441_n N_A_618_89#_c_1124_n 0.00599689f $X=7.805 $Y=1
+ $X2=3.165 $Y2=1.205
cc_448 N_A_110_115#_c_441_n N_A_618_89#_M1020_g 0.00631256f $X=7.805 $Y=1
+ $X2=5.515 $Y2=0.835
cc_449 N_A_110_115#_c_441_n N_A_618_89#_c_1142_n 0.0198218f $X=7.805 $Y=1
+ $X2=6.52 $Y2=0.755
cc_450 N_A_110_115#_c_441_n N_A_1160_89#_M1012_d 0.00142852f $X=7.805 $Y=1
+ $X2=7.33 $Y2=0.575
cc_451 N_A_110_115#_c_418_n N_A_1160_89#_M1016_g 0.00187137f $X=7.615 $Y=1.52
+ $X2=8.635 $Y2=0.755
cc_452 N_A_110_115#_c_441_n N_A_1160_89#_c_1326_n 0.00599085f $X=7.805 $Y=1
+ $X2=5.89 $Y2=1.205
cc_453 N_A_110_115#_c_441_n N_A_1160_89#_c_1330_n 5.89421e-19 $X=7.805 $Y=1
+ $X2=5.89 $Y2=1.365
cc_454 N_A_110_115#_M1030_g N_A_1160_89#_c_1336_n 0.00507506f $X=7.615 $Y=3.445
+ $X2=8.52 $Y2=1.74
cc_455 N_A_110_115#_c_439_n N_A_1160_89#_c_1337_n 2.80323e-19 $X=7.89 $Y=1.21
+ $X2=8.522 $Y2=1.575
cc_456 N_A_110_115#_c_466_n N_A_1160_89#_c_1337_n 6.06666e-19 $X=7.89 $Y=1.37
+ $X2=8.522 $Y2=1.575
cc_457 N_A_110_115#_c_418_n N_A_1160_89#_c_1338_n 0.00416492f $X=7.615 $Y=1.52
+ $X2=8.61 $Y2=1.32
cc_458 N_A_110_115#_c_439_n N_A_1160_89#_c_1338_n 4.20096e-19 $X=7.89 $Y=1.21
+ $X2=8.61 $Y2=1.32
cc_459 N_A_110_115#_M1030_g N_A_1160_89#_c_1371_n 0.00633587f $X=7.615 $Y=3.445
+ $X2=7.385 $Y2=3.045
cc_460 N_A_110_115#_c_418_n N_A_1160_89#_c_1344_n 0.00411162f $X=7.615 $Y=1.52
+ $X2=7.47 $Y2=0.74
cc_461 N_A_110_115#_M1030_g N_A_1160_89#_c_1344_n 0.00587172f $X=7.615 $Y=3.445
+ $X2=7.47 $Y2=0.74
cc_462 N_A_110_115#_c_421_n N_A_1160_89#_c_1344_n 0.00633298f $X=7.685 $Y=1.045
+ $X2=7.47 $Y2=0.74
cc_463 N_A_110_115#_c_439_n N_A_1160_89#_c_1344_n 0.0182754f $X=7.89 $Y=1.21
+ $X2=7.47 $Y2=0.74
cc_464 N_A_110_115#_c_441_n N_A_1160_89#_c_1344_n 0.026518f $X=7.805 $Y=1
+ $X2=7.47 $Y2=0.74
cc_465 N_A_110_115#_c_565_p N_A_1160_89#_c_1344_n 0.00235259f $X=7.89 $Y=1.255
+ $X2=7.47 $Y2=0.74
cc_466 N_A_110_115#_c_466_n N_A_1160_89#_c_1344_n 0.00254925f $X=7.89 $Y=1.37
+ $X2=7.47 $Y2=0.74
cc_467 N_A_110_115#_M1030_g N_A_1160_89#_c_1347_n 0.0483827f $X=7.615 $Y=3.445
+ $X2=7.47 $Y2=2.96
cc_468 N_A_110_115#_c_418_n N_A_1160_89#_c_1348_n 0.00465519f $X=7.615 $Y=1.52
+ $X2=8.52 $Y2=1.74
cc_469 N_A_110_115#_M1030_g N_A_1160_89#_c_1348_n 0.0118805f $X=7.615 $Y=3.445
+ $X2=8.52 $Y2=1.74
cc_470 N_A_110_115#_c_439_n N_A_1160_89#_c_1348_n 0.0151944f $X=7.89 $Y=1.21
+ $X2=8.52 $Y2=1.74
cc_471 N_A_110_115#_c_441_n N_A_1160_89#_c_1348_n 0.00335122f $X=7.805 $Y=1
+ $X2=8.52 $Y2=1.74
cc_472 N_A_110_115#_c_466_n N_A_1160_89#_c_1348_n 0.00122291f $X=7.89 $Y=1.37
+ $X2=8.52 $Y2=1.74
cc_473 N_A_110_115#_M1030_g N_A_1160_89#_c_1349_n 0.00122231f $X=7.615 $Y=3.445
+ $X2=7.47 $Y2=1.74
cc_474 N_A_110_115#_c_418_n N_A_1160_89#_c_1355_n 0.00234211f $X=7.615 $Y=1.52
+ $X2=8.375 $Y2=1.74
cc_475 N_A_110_115#_M1030_g N_A_1160_89#_c_1355_n 0.0111655f $X=7.615 $Y=3.445
+ $X2=8.375 $Y2=1.74
cc_476 N_A_110_115#_c_439_n N_A_1160_89#_c_1355_n 0.00196064f $X=7.89 $Y=1.21
+ $X2=8.375 $Y2=1.74
cc_477 N_A_110_115#_c_466_n N_A_1160_89#_c_1355_n 0.028449f $X=7.89 $Y=1.37
+ $X2=8.375 $Y2=1.74
cc_478 N_A_110_115#_c_441_n N_A_998_115#_M1019_d 0.0032738f $X=7.805 $Y=1
+ $X2=4.99 $Y2=0.575
cc_479 N_A_110_115#_c_421_n N_A_998_115#_M1012_g 0.0121747f $X=7.685 $Y=1.045
+ $X2=7.255 $Y2=0.755
cc_480 N_A_110_115#_c_441_n N_A_998_115#_M1012_g 0.00926356f $X=7.805 $Y=1
+ $X2=7.255 $Y2=0.755
cc_481 N_A_110_115#_M1030_g N_A_998_115#_M1006_g 0.0780098f $X=7.615 $Y=3.445
+ $X2=7.255 $Y2=3.445
cc_482 N_A_110_115#_c_418_n N_A_998_115#_c_1538_n 0.0901845f $X=7.615 $Y=1.52
+ $X2=7.13 $Y2=1.37
cc_483 N_A_110_115#_c_441_n N_A_998_115#_c_1538_n 7.9412e-19 $X=7.805 $Y=1
+ $X2=7.13 $Y2=1.37
cc_484 N_A_110_115#_c_441_n N_A_998_115#_c_1540_n 0.00554379f $X=7.805 $Y=1
+ $X2=4.635 $Y2=1.37
cc_485 N_A_110_115#_c_441_n N_A_998_115#_c_1541_n 0.00648735f $X=7.805 $Y=1
+ $X2=5.315 $Y2=1.37
cc_486 N_A_110_115#_c_441_n N_A_998_115#_c_1542_n 0.00307345f $X=7.805 $Y=1
+ $X2=7.13 $Y2=1.37
cc_487 N_A_110_115#_c_441_n N_A_998_115#_c_1544_n 0.0230872f $X=7.805 $Y=1
+ $X2=5.215 $Y2=0.755
cc_488 N_A_110_115#_c_441_n N_A_998_115#_c_1547_n 0.0328521f $X=7.805 $Y=1
+ $X2=5.18 $Y2=1.37
cc_489 N_A_110_115#_c_441_n N_A_998_115#_c_1548_n 0.0259499f $X=7.805 $Y=1
+ $X2=4.78 $Y2=1.37
cc_490 N_A_110_115#_c_441_n N_A_998_115#_c_1549_n 0.12896f $X=7.805 $Y=1
+ $X2=6.985 $Y2=1.37
cc_491 N_A_110_115#_c_441_n N_A_998_115#_c_1551_n 0.0224792f $X=7.805 $Y=1
+ $X2=5.44 $Y2=1.37
cc_492 N_A_110_115#_c_441_n N_A_998_115#_c_1552_n 0.0259663f $X=7.805 $Y=1
+ $X2=7.13 $Y2=1.37
cc_493 N_A_110_115#_c_466_n N_A_998_115#_c_1552_n 0.0127174f $X=7.89 $Y=1.37
+ $X2=7.13 $Y2=1.37
cc_494 N_A_110_115#_c_418_n N_QN_c_1681_n 0.00222227f $X=7.615 $Y=1.52 $X2=8.42
+ $Y2=0.74
cc_495 N_A_110_115#_c_421_n N_QN_c_1681_n 0.00298655f $X=7.685 $Y=1.045 $X2=8.42
+ $Y2=0.74
cc_496 N_A_110_115#_c_439_n N_QN_c_1681_n 0.00781846f $X=7.89 $Y=1.21 $X2=8.42
+ $Y2=0.74
cc_497 N_A_110_115#_c_441_n N_QN_c_1681_n 0.00875851f $X=7.805 $Y=1 $X2=8.42
+ $Y2=0.74
cc_498 N_A_110_115#_c_565_p N_QN_c_1681_n 7.96604e-19 $X=7.89 $Y=1.255 $X2=8.42
+ $Y2=0.74
cc_499 N_A_110_115#_c_466_n N_QN_c_1681_n 2.00168e-19 $X=7.89 $Y=1.37 $X2=8.42
+ $Y2=0.74
cc_500 N_A_110_115#_M1030_g N_QN_c_1685_n 0.0144714f $X=7.615 $Y=3.445 $X2=8.42
+ $Y2=2.48
cc_501 N_A_110_115#_c_418_n N_QN_c_1688_n 6.86262e-19 $X=7.615 $Y=1.52 $X2=8.505
+ $Y2=1.37
cc_502 N_A_110_115#_c_439_n N_QN_c_1688_n 0.00565014f $X=7.89 $Y=1.21 $X2=8.505
+ $Y2=1.37
cc_503 N_A_110_115#_c_466_n N_QN_c_1688_n 0.00464864f $X=7.89 $Y=1.37 $X2=8.505
+ $Y2=1.37
cc_504 N_A_110_115#_M1030_g N_QN_c_1690_n 0.00423893f $X=7.615 $Y=3.445
+ $X2=8.505 $Y2=2.285
cc_505 N_A_110_115#_M1030_g QN 0.00472165f $X=7.615 $Y=3.445 $X2=8.425 $Y2=2.48
cc_506 N_A_110_115#_c_441_n A_576_115# 0.00381028f $X=7.805 $Y=1 $X2=2.88
+ $Y2=0.575
cc_507 N_A_110_115#_c_441_n A_768_115# 0.00473401f $X=7.805 $Y=1 $X2=3.84
+ $Y2=0.575
cc_508 N_A_110_115#_c_441_n A_926_115# 0.00429254f $X=7.805 $Y=1 $X2=4.63
+ $Y2=0.575
cc_509 N_A_110_115#_c_441_n A_1118_115# 0.00465218f $X=7.805 $Y=1 $X2=5.59
+ $Y2=0.575
cc_510 N_A_342_442#_c_615_n N_D_M1007_g 0.0137346f $X=2.11 $Y=2.21 $X2=2.805
+ $Y2=0.835
cc_511 N_A_342_442#_c_616_n N_D_M1007_g 0.0122665f $X=3.28 $Y=1.285 $X2=2.805
+ $Y2=0.835
cc_512 N_A_342_442#_c_618_n N_D_M1007_g 0.00158134f $X=2.2 $Y=1.285 $X2=2.805
+ $Y2=0.835
cc_513 N_A_342_442#_c_614_n N_D_M1028_g 0.00395324f $X=1.94 $Y=2.375 $X2=2.805
+ $Y2=3.235
cc_514 N_A_342_442#_c_631_n N_D_M1028_g 0.0211478f $X=3.295 $Y=2.705 $X2=2.805
+ $Y2=3.235
cc_515 N_A_342_442#_c_621_n N_D_M1028_g 0.00767395f $X=1.94 $Y=2.375 $X2=2.805
+ $Y2=3.235
cc_516 N_A_342_442#_c_616_n N_D_c_698_n 0.00207628f $X=3.28 $Y=1.285 $X2=2.865
+ $Y2=1.74
cc_517 N_A_342_442#_c_615_n N_D_c_699_n 0.00613892f $X=2.11 $Y=2.21 $X2=2.865
+ $Y2=1.74
cc_518 N_A_342_442#_c_616_n N_D_c_699_n 0.0086486f $X=3.28 $Y=1.285 $X2=2.865
+ $Y2=1.74
cc_519 N_A_342_442#_c_615_n D 0.0055149f $X=2.11 $Y=2.21 $X2=2.865 $Y2=1.74
cc_520 N_A_342_442#_c_616_n D 0.00200799f $X=3.28 $Y=1.285 $X2=2.865 $Y2=1.74
cc_521 N_A_342_442#_c_631_n N_CK_M1024_g 0.0153421f $X=3.295 $Y=2.705 $X2=3.165
+ $Y2=3.235
cc_522 N_A_342_442#_c_631_n N_CK_c_742_n 0.00150627f $X=3.295 $Y=2.705 $X2=3.225
+ $Y2=2.285
cc_523 N_A_342_442#_c_616_n N_CK_c_743_n 9.45214e-19 $X=3.28 $Y=1.285 $X2=3.705
+ $Y2=1.37
cc_524 N_A_342_442#_c_622_n N_CK_c_743_n 0.00165184f $X=3.365 $Y=0.755 $X2=3.705
+ $Y2=1.37
cc_525 N_A_342_442#_c_620_n N_CK_c_744_n 0.00464203f $X=3.365 $Y=1.2 $X2=3.705
+ $Y2=1.205
cc_526 N_A_342_442#_c_622_n N_CK_c_744_n 0.00243799f $X=3.365 $Y=0.755 $X2=3.705
+ $Y2=1.205
cc_527 N_A_342_442#_c_631_n N_CK_c_753_n 0.00883015f $X=3.295 $Y=2.705 $X2=3.62
+ $Y2=2.11
cc_528 N_A_342_442#_c_616_n N_CK_c_753_n 0.0019742f $X=3.28 $Y=1.285 $X2=3.62
+ $Y2=2.11
cc_529 N_A_342_442#_c_616_n N_CK_c_754_n 0.012316f $X=3.28 $Y=1.285 $X2=3.705
+ $Y2=1.37
cc_530 N_A_342_442#_c_622_n N_CK_c_754_n 5.6626e-19 $X=3.365 $Y=0.755 $X2=3.705
+ $Y2=1.37
cc_531 N_A_342_442#_c_631_n N_CK_c_759_n 0.0101098f $X=3.295 $Y=2.705 $X2=3.225
+ $Y2=2.11
cc_532 N_A_342_442#_c_616_n N_CK_c_759_n 0.00224443f $X=3.28 $Y=1.285 $X2=3.225
+ $Y2=2.11
cc_533 N_A_342_442#_c_631_n N_CK_c_761_n 0.00601583f $X=3.295 $Y=2.705 $X2=5.31
+ $Y2=2.11
cc_534 N_A_342_442#_c_631_n N_CK_c_762_n 0.00409373f $X=3.295 $Y=2.705 $X2=3.37
+ $Y2=2.11
cc_535 N_A_342_442#_c_621_n N_A_217_605#_c_999_n 0.0100421f $X=1.94 $Y=2.375
+ $X2=1.21 $Y2=3.275
cc_536 N_A_342_442#_M1005_g N_A_217_605#_c_1000_n 0.00176497f $X=1.855 $Y=0.755
+ $X2=1.555 $Y2=1.81
cc_537 N_A_342_442#_c_614_n N_A_217_605#_c_1000_n 6.21732e-19 $X=1.94 $Y=2.375
+ $X2=1.555 $Y2=1.81
cc_538 N_A_342_442#_c_615_n N_A_217_605#_c_1000_n 0.00954176f $X=2.11 $Y=2.21
+ $X2=1.555 $Y2=1.81
cc_539 N_A_342_442#_M1005_g N_A_217_605#_c_1002_n 0.0102637f $X=1.855 $Y=0.755
+ $X2=1.64 $Y2=0.74
cc_540 N_A_342_442#_c_615_n N_A_217_605#_c_1002_n 0.012524f $X=2.11 $Y=2.21
+ $X2=1.64 $Y2=0.74
cc_541 N_A_342_442#_c_618_n N_A_217_605#_c_1002_n 0.011766f $X=2.2 $Y=1.285
+ $X2=1.64 $Y2=0.74
cc_542 N_A_342_442#_M1005_g N_A_217_605#_c_1008_n 0.0112415f $X=1.855 $Y=0.755
+ $X2=4.06 $Y2=1.37
cc_543 N_A_342_442#_c_616_n N_A_217_605#_c_1008_n 0.0476148f $X=3.28 $Y=1.285
+ $X2=4.06 $Y2=1.37
cc_544 N_A_342_442#_c_618_n N_A_217_605#_c_1008_n 0.0198865f $X=2.2 $Y=1.285
+ $X2=4.06 $Y2=1.37
cc_545 N_A_342_442#_c_622_n N_A_217_605#_c_1008_n 8.84066e-19 $X=3.365 $Y=0.755
+ $X2=4.06 $Y2=1.37
cc_546 N_A_342_442#_M1005_g N_A_217_605#_c_1009_n 0.00236248f $X=1.855 $Y=0.755
+ $X2=1.78 $Y2=1.372
cc_547 N_A_342_442#_c_615_n N_A_217_605#_c_1009_n 6.00227e-19 $X=2.11 $Y=2.21
+ $X2=1.78 $Y2=1.372
cc_548 N_A_342_442#_c_618_n N_A_217_605#_c_1009_n 0.00125688f $X=2.2 $Y=1.285
+ $X2=1.78 $Y2=1.372
cc_549 N_A_342_442#_c_616_n N_A_618_89#_c_1124_n 0.0022787f $X=3.28 $Y=1.285
+ $X2=3.165 $Y2=1.205
cc_550 N_A_342_442#_c_620_n N_A_618_89#_c_1124_n 0.00492892f $X=3.365 $Y=1.2
+ $X2=3.165 $Y2=1.205
cc_551 N_A_342_442#_c_622_n N_A_618_89#_c_1124_n 0.00116801f $X=3.365 $Y=0.755
+ $X2=3.165 $Y2=1.205
cc_552 N_A_342_442#_c_616_n N_A_618_89#_c_1127_n 0.00326059f $X=3.28 $Y=1.285
+ $X2=3.285 $Y2=1.745
cc_553 N_A_342_442#_c_616_n N_A_618_89#_c_1137_n 0.00984832f $X=3.28 $Y=1.285
+ $X2=3.285 $Y2=1.28
cc_554 N_A_342_442#_c_631_n A_576_521# 0.00732587f $X=3.295 $Y=2.705 $X2=2.88
+ $Y2=2.605
cc_555 N_D_M1028_g N_CK_c_742_n 0.11474f $X=2.805 $Y=3.235 $X2=3.225 $Y2=2.285
cc_556 N_D_c_698_n N_CK_c_754_n 2.89615e-19 $X=2.865 $Y=1.74 $X2=3.705 $Y2=1.37
cc_557 N_D_c_699_n N_CK_c_754_n 0.00478177f $X=2.865 $Y=1.74 $X2=3.705 $Y2=1.37
cc_558 D N_CK_c_754_n 0.00551577f $X=2.865 $Y=1.74 $X2=3.705 $Y2=1.37
cc_559 N_D_M1028_g N_CK_c_759_n 0.00494364f $X=2.805 $Y=3.235 $X2=3.225 $Y2=2.11
cc_560 N_D_M1028_g N_CK_c_762_n 0.00515433f $X=2.805 $Y=3.235 $X2=3.37 $Y2=2.11
cc_561 D N_CK_c_762_n 0.00375733f $X=2.865 $Y=1.74 $X2=3.37 $Y2=2.11
cc_562 N_D_M1007_g N_A_217_605#_c_1008_n 0.0030176f $X=2.805 $Y=0.835 $X2=4.06
+ $Y2=1.37
cc_563 N_D_c_698_n N_A_217_605#_c_1008_n 7.9412e-19 $X=2.865 $Y=1.74 $X2=4.06
+ $Y2=1.37
cc_564 N_D_c_699_n N_A_217_605#_c_1008_n 0.00111625f $X=2.865 $Y=1.74 $X2=4.06
+ $Y2=1.37
cc_565 D N_A_217_605#_c_1008_n 0.0353362f $X=2.865 $Y=1.74 $X2=4.06 $Y2=1.37
cc_566 N_D_M1007_g N_A_618_89#_c_1124_n 0.0567053f $X=2.805 $Y=0.835 $X2=3.165
+ $Y2=1.205
cc_567 N_D_M1007_g N_A_618_89#_c_1127_n 0.00932846f $X=2.805 $Y=0.835 $X2=3.285
+ $Y2=1.745
cc_568 N_D_c_698_n N_A_618_89#_c_1127_n 0.0210215f $X=2.865 $Y=1.74 $X2=3.285
+ $Y2=1.745
cc_569 N_D_c_699_n N_A_618_89#_c_1127_n 0.00164409f $X=2.865 $Y=1.74 $X2=3.285
+ $Y2=1.745
cc_570 D N_A_618_89#_c_1127_n 0.00342011f $X=2.865 $Y=1.74 $X2=3.285 $Y2=1.745
cc_571 D N_A_618_89#_c_1129_n 4.62757e-19 $X=2.865 $Y=1.74 $X2=3.36 $Y2=1.82
cc_572 N_CK_c_744_n N_A_217_605#_M1027_g 0.0338208f $X=3.705 $Y=1.205 $X2=4.125
+ $Y2=0.835
cc_573 N_CK_c_754_n N_A_217_605#_M1027_g 0.00109079f $X=3.705 $Y=1.37 $X2=4.125
+ $Y2=0.835
cc_574 N_CK_c_747_n N_A_217_605#_c_990_n 0.0333732f $X=4.975 $Y=1.37 $X2=4.48
+ $Y2=1.37
cc_575 N_CK_c_743_n N_A_217_605#_c_992_n 0.0338208f $X=3.705 $Y=1.37 $X2=4.2
+ $Y2=1.37
cc_576 N_CK_c_761_n N_A_217_605#_c_993_n 0.00772879f $X=5.31 $Y=2.11 $X2=4.48
+ $Y2=2.285
cc_577 N_CK_c_761_n N_A_217_605#_c_994_n 0.00679967f $X=5.31 $Y=2.11 $X2=4.2
+ $Y2=2.285
cc_578 N_CK_c_748_n N_A_217_605#_M1025_g 0.0333732f $X=4.975 $Y=1.205 $X2=4.555
+ $Y2=0.835
cc_579 N_CK_c_755_n N_A_217_605#_M1025_g 3.67139e-19 $X=4.975 $Y=1.37 $X2=4.555
+ $Y2=0.835
cc_580 N_CK_c_743_n N_A_217_605#_c_1005_n 7.30049e-19 $X=3.705 $Y=1.37 $X2=4.295
+ $Y2=2.285
cc_581 N_CK_c_753_n N_A_217_605#_c_1005_n 0.00401809f $X=3.62 $Y=2.11 $X2=4.295
+ $Y2=2.285
cc_582 N_CK_c_754_n N_A_217_605#_c_1005_n 0.0203851f $X=3.705 $Y=1.37 $X2=4.295
+ $Y2=2.285
cc_583 N_CK_c_761_n N_A_217_605#_c_1005_n 0.0206884f $X=5.31 $Y=2.11 $X2=4.295
+ $Y2=2.285
cc_584 N_CK_c_743_n N_A_217_605#_c_1006_n 7.18106e-19 $X=3.705 $Y=1.37 $X2=4.295
+ $Y2=1.37
cc_585 N_CK_c_754_n N_A_217_605#_c_1006_n 0.00742068f $X=3.705 $Y=1.37 $X2=4.295
+ $Y2=1.37
cc_586 N_CK_c_761_n N_A_217_605#_c_1006_n 0.00102309f $X=5.31 $Y=2.11 $X2=4.295
+ $Y2=1.37
cc_587 N_CK_c_743_n N_A_217_605#_c_1008_n 0.00383172f $X=3.705 $Y=1.37 $X2=4.06
+ $Y2=1.37
cc_588 N_CK_c_753_n N_A_217_605#_c_1008_n 0.00443421f $X=3.62 $Y=2.11 $X2=4.06
+ $Y2=1.37
cc_589 N_CK_c_754_n N_A_217_605#_c_1008_n 0.0149971f $X=3.705 $Y=1.37 $X2=4.06
+ $Y2=1.37
cc_590 N_CK_c_759_n N_A_217_605#_c_1008_n 7.12046e-19 $X=3.225 $Y=2.11 $X2=4.06
+ $Y2=1.37
cc_591 N_CK_c_762_n N_A_217_605#_c_1008_n 0.0126164f $X=3.37 $Y=2.11 $X2=4.06
+ $Y2=1.37
cc_592 N_CK_c_743_n N_A_217_605#_c_1058_n 3.3031e-19 $X=3.705 $Y=1.37 $X2=4.205
+ $Y2=1.37
cc_593 N_CK_c_754_n N_A_217_605#_c_1058_n 0.00143592f $X=3.705 $Y=1.37 $X2=4.205
+ $Y2=1.37
cc_594 N_CK_c_761_n N_A_217_605#_c_1058_n 0.0129652f $X=5.31 $Y=2.11 $X2=4.205
+ $Y2=1.37
cc_595 N_CK_c_744_n N_A_618_89#_c_1124_n 0.0171207f $X=3.705 $Y=1.205 $X2=3.165
+ $Y2=1.205
cc_596 N_CK_c_754_n N_A_618_89#_c_1127_n 0.00613747f $X=3.705 $Y=1.37 $X2=3.285
+ $Y2=1.745
cc_597 N_CK_c_743_n N_A_618_89#_c_1128_n 0.0183603f $X=3.705 $Y=1.37 $X2=3.69
+ $Y2=1.82
cc_598 N_CK_c_754_n N_A_618_89#_c_1128_n 0.00630484f $X=3.705 $Y=1.37 $X2=3.69
+ $Y2=1.82
cc_599 N_CK_c_761_n N_A_618_89#_c_1128_n 0.00613485f $X=5.31 $Y=2.11 $X2=3.69
+ $Y2=1.82
cc_600 N_CK_c_742_n N_A_618_89#_c_1129_n 0.00904036f $X=3.225 $Y=2.285 $X2=3.36
+ $Y2=1.82
cc_601 N_CK_c_753_n N_A_618_89#_c_1129_n 0.00878348f $X=3.62 $Y=2.11 $X2=3.36
+ $Y2=1.82
cc_602 N_CK_c_759_n N_A_618_89#_c_1129_n 0.00109468f $X=3.225 $Y=2.11 $X2=3.36
+ $Y2=1.82
cc_603 N_CK_c_762_n N_A_618_89#_c_1129_n 0.00137501f $X=3.37 $Y=2.11 $X2=3.36
+ $Y2=1.82
cc_604 N_CK_M1024_g N_A_618_89#_M1017_g 0.0316011f $X=3.165 $Y=3.235 $X2=3.765
+ $Y2=3.235
cc_605 N_CK_c_742_n N_A_618_89#_M1017_g 0.0128384f $X=3.225 $Y=2.285 $X2=3.765
+ $Y2=3.235
cc_606 N_CK_c_753_n N_A_618_89#_M1017_g 0.0081071f $X=3.62 $Y=2.11 $X2=3.765
+ $Y2=3.235
cc_607 N_CK_c_754_n N_A_618_89#_M1017_g 0.00478024f $X=3.705 $Y=1.37 $X2=3.765
+ $Y2=3.235
cc_608 N_CK_c_759_n N_A_618_89#_M1017_g 0.00184124f $X=3.225 $Y=2.11 $X2=3.765
+ $Y2=3.235
cc_609 N_CK_c_761_n N_A_618_89#_M1017_g 0.00938974f $X=5.31 $Y=2.11 $X2=3.765
+ $Y2=3.235
cc_610 N_CK_c_762_n N_A_618_89#_M1017_g 4.2e-19 $X=3.37 $Y=2.11 $X2=3.765
+ $Y2=3.235
cc_611 N_CK_c_761_n N_A_618_89#_c_1131_n 0.00607908f $X=5.31 $Y=2.11 $X2=4.84
+ $Y2=1.82
cc_612 N_CK_M1000_g N_A_618_89#_M1003_g 0.0316011f $X=5.515 $Y=3.235 $X2=4.915
+ $Y2=3.235
cc_613 N_CK_c_751_n N_A_618_89#_M1003_g 0.0118393f $X=5.455 $Y=2.285 $X2=4.915
+ $Y2=3.235
cc_614 N_CK_c_755_n N_A_618_89#_M1003_g 0.00399495f $X=4.975 $Y=1.37 $X2=4.915
+ $Y2=3.235
cc_615 N_CK_c_757_n N_A_618_89#_M1003_g 0.00654233f $X=5.06 $Y=2.11 $X2=4.915
+ $Y2=3.235
cc_616 N_CK_c_760_n N_A_618_89#_M1003_g 0.00128351f $X=5.455 $Y=2.11 $X2=4.915
+ $Y2=3.235
cc_617 N_CK_c_761_n N_A_618_89#_M1003_g 0.00497421f $X=5.31 $Y=2.11 $X2=4.915
+ $Y2=3.235
cc_618 N_CK_c_764_n N_A_618_89#_M1003_g 4.2e-19 $X=5.6 $Y=2.11 $X2=4.915
+ $Y2=3.235
cc_619 N_CK_c_755_n N_A_618_89#_c_1133_n 0.00635358f $X=4.975 $Y=1.37 $X2=5.32
+ $Y2=1.82
cc_620 N_CK_c_756_n N_A_618_89#_c_1133_n 0.00842176f $X=5.37 $Y=2.11 $X2=5.32
+ $Y2=1.82
cc_621 N_CK_c_761_n N_A_618_89#_c_1133_n 0.00519056f $X=5.31 $Y=2.11 $X2=5.32
+ $Y2=1.82
cc_622 N_CK_c_764_n N_A_618_89#_c_1133_n 0.00150125f $X=5.6 $Y=2.11 $X2=5.32
+ $Y2=1.82
cc_623 N_CK_c_747_n N_A_618_89#_M1020_g 0.012357f $X=4.975 $Y=1.37 $X2=5.515
+ $Y2=0.835
cc_624 N_CK_c_748_n N_A_618_89#_M1020_g 0.017109f $X=4.975 $Y=1.205 $X2=5.515
+ $Y2=0.835
cc_625 N_CK_c_755_n N_A_618_89#_M1020_g 4.67639e-19 $X=4.975 $Y=1.37 $X2=5.515
+ $Y2=0.835
cc_626 N_CK_c_743_n N_A_618_89#_c_1137_n 0.0216263f $X=3.705 $Y=1.37 $X2=3.285
+ $Y2=1.28
cc_627 N_CK_c_759_n N_A_618_89#_c_1137_n 2.45465e-19 $X=3.225 $Y=2.11 $X2=3.285
+ $Y2=1.28
cc_628 N_CK_c_754_n N_A_618_89#_c_1138_n 0.00568091f $X=3.705 $Y=1.37 $X2=3.765
+ $Y2=1.82
cc_629 N_CK_c_747_n N_A_618_89#_c_1139_n 0.0183603f $X=4.975 $Y=1.37 $X2=4.915
+ $Y2=1.82
cc_630 N_CK_c_755_n N_A_618_89#_c_1139_n 0.00436024f $X=4.975 $Y=1.37 $X2=4.915
+ $Y2=1.82
cc_631 N_CK_c_747_n N_A_618_89#_c_1140_n 9.99307e-19 $X=4.975 $Y=1.37 $X2=5.455
+ $Y2=1.725
cc_632 N_CK_c_751_n N_A_618_89#_c_1140_n 0.0165037f $X=5.455 $Y=2.285 $X2=5.455
+ $Y2=1.725
cc_633 N_CK_c_755_n N_A_618_89#_c_1140_n 0.003871f $X=4.975 $Y=1.37 $X2=5.455
+ $Y2=1.725
cc_634 N_CK_c_760_n N_A_618_89#_c_1140_n 0.0010914f $X=5.455 $Y=2.11 $X2=5.455
+ $Y2=1.725
cc_635 N_CK_c_763_n N_A_618_89#_c_1140_n 3.23651e-19 $X=6.305 $Y=2.11 $X2=5.455
+ $Y2=1.725
cc_636 N_CK_c_751_n N_A_618_89#_c_1141_n 7.90579e-19 $X=5.455 $Y=2.285 $X2=5.455
+ $Y2=1.725
cc_637 N_CK_c_755_n N_A_618_89#_c_1141_n 0.0107188f $X=4.975 $Y=1.37 $X2=5.455
+ $Y2=1.725
cc_638 N_CK_c_756_n N_A_618_89#_c_1141_n 0.00447505f $X=5.37 $Y=2.11 $X2=5.455
+ $Y2=1.725
cc_639 N_CK_c_760_n N_A_618_89#_c_1141_n 0.00985566f $X=5.455 $Y=2.11 $X2=5.455
+ $Y2=1.725
cc_640 N_CK_c_763_n N_A_618_89#_c_1141_n 2.90862e-19 $X=6.305 $Y=2.11 $X2=5.455
+ $Y2=1.725
cc_641 N_CK_c_764_n N_A_618_89#_c_1141_n 0.0019318f $X=5.6 $Y=2.11 $X2=5.455
+ $Y2=1.725
cc_642 N_CK_c_735_n N_A_618_89#_c_1142_n 0.00793442f $X=6.305 $Y=1.205 $X2=6.52
+ $Y2=0.755
cc_643 N_CK_c_741_n N_A_618_89#_c_1142_n 0.00847232f $X=6.385 $Y=2.12 $X2=6.52
+ $Y2=0.755
cc_644 N_CK_c_752_n N_A_618_89#_c_1142_n 0.00540063f $X=6.385 $Y=1.28 $X2=6.52
+ $Y2=0.755
cc_645 N_CK_c_740_n N_A_618_89#_c_1147_n 0.0031983f $X=6.305 $Y=2.45 $X2=6.795
+ $Y2=2.62
cc_646 N_CK_M1029_g N_A_618_89#_c_1147_n 0.00397698f $X=6.305 $Y=3.235 $X2=6.795
+ $Y2=2.62
cc_647 N_CK_c_741_n N_A_618_89#_c_1147_n 0.0027512f $X=6.385 $Y=2.12 $X2=6.795
+ $Y2=2.62
cc_648 N_CK_c_758_n N_A_618_89#_c_1147_n 0.02768f $X=6.45 $Y=2.11 $X2=6.795
+ $Y2=2.62
cc_649 CK N_A_618_89#_c_1147_n 0.00176523f $X=6.45 $Y=2.11 $X2=6.795 $Y2=2.62
cc_650 N_CK_c_740_n N_A_618_89#_c_1148_n 0.00296017f $X=6.305 $Y=2.45 $X2=6.52
+ $Y2=1.725
cc_651 N_CK_c_741_n N_A_618_89#_c_1148_n 0.0119539f $X=6.385 $Y=2.12 $X2=6.52
+ $Y2=1.725
cc_652 N_CK_c_752_n N_A_618_89#_c_1148_n 8.36012e-19 $X=6.385 $Y=1.28 $X2=6.52
+ $Y2=1.725
cc_653 N_CK_c_758_n N_A_618_89#_c_1148_n 0.00983573f $X=6.45 $Y=2.11 $X2=6.52
+ $Y2=1.725
cc_654 N_CK_c_763_n N_A_618_89#_c_1148_n 2.10751e-19 $X=6.305 $Y=2.11 $X2=6.52
+ $Y2=1.725
cc_655 CK N_A_618_89#_c_1148_n 0.00406363f $X=6.45 $Y=2.11 $X2=6.52 $Y2=1.725
cc_656 N_CK_c_740_n N_A_618_89#_c_1161_n 0.00233159f $X=6.305 $Y=2.45 $X2=6.795
+ $Y2=2.705
cc_657 N_CK_c_758_n N_A_618_89#_c_1161_n 0.00601935f $X=6.45 $Y=2.11 $X2=6.795
+ $Y2=2.705
cc_658 N_CK_c_763_n N_A_618_89#_c_1149_n 0.0504038f $X=6.305 $Y=2.11 $X2=6.215
+ $Y2=1.74
cc_659 N_CK_c_755_n N_A_618_89#_c_1241_n 0.00243046f $X=4.975 $Y=1.37 $X2=5.6
+ $Y2=1.74
cc_660 N_CK_c_760_n N_A_618_89#_c_1241_n 4.75808e-19 $X=5.455 $Y=2.11 $X2=5.6
+ $Y2=1.74
cc_661 N_CK_c_764_n N_A_618_89#_c_1241_n 0.0296144f $X=5.6 $Y=2.11 $X2=5.6
+ $Y2=1.74
cc_662 N_CK_c_741_n N_A_618_89#_c_1150_n 0.00233584f $X=6.385 $Y=2.12 $X2=6.36
+ $Y2=1.74
cc_663 N_CK_c_752_n N_A_618_89#_c_1150_n 3.99064e-19 $X=6.385 $Y=1.28 $X2=6.36
+ $Y2=1.74
cc_664 N_CK_c_758_n N_A_618_89#_c_1150_n 5.59009e-19 $X=6.45 $Y=2.11 $X2=6.36
+ $Y2=1.74
cc_665 N_CK_c_763_n N_A_618_89#_c_1150_n 0.0083989f $X=6.305 $Y=2.11 $X2=6.36
+ $Y2=1.74
cc_666 CK N_A_618_89#_c_1150_n 0.0208541f $X=6.45 $Y=2.11 $X2=6.36 $Y2=1.74
cc_667 N_CK_M1000_g N_A_1160_89#_M1009_g 0.0565466f $X=5.515 $Y=3.235 $X2=5.875
+ $Y2=3.235
cc_668 N_CK_c_740_n N_A_1160_89#_M1009_g 0.042164f $X=6.305 $Y=2.45 $X2=5.875
+ $Y2=3.235
cc_669 N_CK_c_758_n N_A_1160_89#_M1009_g 2.2703e-19 $X=6.45 $Y=2.11 $X2=5.875
+ $Y2=3.235
cc_670 N_CK_c_735_n N_A_1160_89#_c_1326_n 0.0168538f $X=6.305 $Y=1.205 $X2=5.89
+ $Y2=1.205
cc_671 N_CK_c_741_n N_A_1160_89#_c_1330_n 0.0099158f $X=6.385 $Y=2.12 $X2=5.89
+ $Y2=1.365
cc_672 N_CK_c_752_n N_A_1160_89#_c_1330_n 0.00839284f $X=6.385 $Y=1.28 $X2=5.89
+ $Y2=1.365
cc_673 N_CK_c_741_n N_A_1160_89#_c_1331_n 0.00681852f $X=6.385 $Y=2.12 $X2=5.89
+ $Y2=2.105
cc_674 N_CK_c_758_n N_A_1160_89#_c_1331_n 3.88594e-19 $X=6.45 $Y=2.11 $X2=5.89
+ $Y2=2.105
cc_675 N_CK_c_760_n N_A_1160_89#_c_1331_n 0.00103465f $X=5.455 $Y=2.11 $X2=5.89
+ $Y2=2.105
cc_676 N_CK_c_763_n N_A_1160_89#_c_1331_n 0.00145834f $X=6.305 $Y=2.11 $X2=5.89
+ $Y2=2.105
cc_677 N_CK_c_764_n N_A_1160_89#_c_1331_n 6.89974e-19 $X=5.6 $Y=2.11 $X2=5.89
+ $Y2=2.105
cc_678 N_CK_c_740_n N_A_1160_89#_c_1332_n 0.00559821f $X=6.305 $Y=2.45 $X2=5.89
+ $Y2=2.255
cc_679 N_CK_c_751_n N_A_1160_89#_c_1332_n 0.0565466f $X=5.455 $Y=2.285 $X2=5.89
+ $Y2=2.255
cc_680 N_CK_c_760_n N_A_1160_89#_c_1332_n 0.0011802f $X=5.455 $Y=2.11 $X2=5.89
+ $Y2=2.255
cc_681 N_CK_c_763_n N_A_1160_89#_c_1332_n 0.00136902f $X=6.305 $Y=2.11 $X2=5.89
+ $Y2=2.255
cc_682 N_CK_c_764_n N_A_1160_89#_c_1332_n 4.36292e-19 $X=5.6 $Y=2.11 $X2=5.89
+ $Y2=2.255
cc_683 N_CK_c_741_n N_A_1160_89#_c_1333_n 0.021525f $X=6.385 $Y=2.12 $X2=5.965
+ $Y2=1.77
cc_684 N_CK_c_763_n N_A_1160_89#_c_1333_n 8.07535e-19 $X=6.305 $Y=2.11 $X2=5.965
+ $Y2=1.77
cc_685 N_CK_c_741_n N_A_1160_89#_c_1341_n 0.00163452f $X=6.385 $Y=2.12 $X2=5.935
+ $Y2=2.025
cc_686 N_CK_c_763_n N_A_1160_89#_c_1341_n 0.00382734f $X=6.305 $Y=2.11 $X2=5.935
+ $Y2=2.025
cc_687 N_CK_c_764_n N_A_1160_89#_c_1341_n 0.00126344f $X=5.6 $Y=2.11 $X2=5.935
+ $Y2=2.025
cc_688 CK N_A_1160_89#_c_1341_n 9.59297e-19 $X=6.45 $Y=2.11 $X2=5.935 $Y2=2.025
cc_689 N_CK_c_740_n N_A_1160_89#_c_1343_n 0.0038598f $X=6.305 $Y=2.45 $X2=5.935
+ $Y2=2.48
cc_690 N_CK_c_741_n N_A_1160_89#_c_1343_n 4.37212e-19 $X=6.385 $Y=2.12 $X2=5.935
+ $Y2=2.48
cc_691 N_CK_c_751_n N_A_1160_89#_c_1343_n 0.00225243f $X=5.455 $Y=2.285
+ $X2=5.935 $Y2=2.48
cc_692 N_CK_c_758_n N_A_1160_89#_c_1343_n 0.0147004f $X=6.45 $Y=2.11 $X2=5.935
+ $Y2=2.48
cc_693 N_CK_c_760_n N_A_1160_89#_c_1343_n 0.0150485f $X=5.455 $Y=2.11 $X2=5.935
+ $Y2=2.48
cc_694 N_CK_c_763_n N_A_1160_89#_c_1343_n 0.011095f $X=6.305 $Y=2.11 $X2=5.935
+ $Y2=2.48
cc_695 N_CK_c_764_n N_A_1160_89#_c_1343_n 8.19742e-19 $X=5.6 $Y=2.11 $X2=5.935
+ $Y2=2.48
cc_696 CK N_A_1160_89#_c_1343_n 7.07735e-19 $X=6.45 $Y=2.11 $X2=5.935 $Y2=2.48
cc_697 N_CK_c_740_n N_A_1160_89#_c_1350_n 0.00414649f $X=6.305 $Y=2.45 $X2=6.735
+ $Y2=2.48
cc_698 N_CK_M1029_g N_A_1160_89#_c_1350_n 0.00886306f $X=6.305 $Y=3.235
+ $X2=6.735 $Y2=2.48
cc_699 N_CK_c_758_n N_A_1160_89#_c_1350_n 0.00641049f $X=6.45 $Y=2.11 $X2=6.735
+ $Y2=2.48
cc_700 N_CK_c_763_n N_A_1160_89#_c_1350_n 0.0190773f $X=6.305 $Y=2.11 $X2=6.735
+ $Y2=2.48
cc_701 CK N_A_1160_89#_c_1350_n 0.025144f $X=6.45 $Y=2.11 $X2=6.735 $Y2=2.48
cc_702 N_CK_c_740_n N_A_1160_89#_c_1351_n 4.83733e-19 $X=6.305 $Y=2.45 $X2=6.08
+ $Y2=2.48
cc_703 N_CK_M1029_g N_A_1160_89#_c_1351_n 4.63789e-19 $X=6.305 $Y=3.235 $X2=6.08
+ $Y2=2.48
cc_704 N_CK_c_751_n N_A_1160_89#_c_1351_n 0.00405956f $X=5.455 $Y=2.285 $X2=6.08
+ $Y2=2.48
cc_705 N_CK_c_758_n N_A_1160_89#_c_1351_n 7.98697e-19 $X=6.45 $Y=2.11 $X2=6.08
+ $Y2=2.48
cc_706 N_CK_c_760_n N_A_1160_89#_c_1351_n 0.0025579f $X=5.455 $Y=2.11 $X2=6.08
+ $Y2=2.48
cc_707 N_CK_c_763_n N_A_1160_89#_c_1351_n 0.0253083f $X=6.305 $Y=2.11 $X2=6.08
+ $Y2=2.48
cc_708 N_CK_c_758_n N_A_1160_89#_c_1352_n 0.00141357f $X=6.45 $Y=2.11 $X2=6.825
+ $Y2=2.395
cc_709 CK N_A_1160_89#_c_1352_n 0.0233707f $X=6.45 $Y=2.11 $X2=6.825 $Y2=2.395
cc_710 N_CK_c_740_n N_A_998_115#_M1006_g 0.00467255f $X=6.305 $Y=2.45 $X2=7.255
+ $Y2=3.445
cc_711 N_CK_c_741_n N_A_998_115#_M1006_g 0.00591235f $X=6.385 $Y=2.12 $X2=7.255
+ $Y2=3.445
cc_712 N_CK_c_752_n N_A_998_115#_c_1538_n 0.00638002f $X=6.385 $Y=1.28 $X2=7.13
+ $Y2=1.37
cc_713 N_CK_c_747_n N_A_998_115#_c_1540_n 0.00215979f $X=4.975 $Y=1.37 $X2=4.635
+ $Y2=1.37
cc_714 N_CK_c_755_n N_A_998_115#_c_1540_n 0.0571231f $X=4.975 $Y=1.37 $X2=4.635
+ $Y2=1.37
cc_715 N_CK_c_757_n N_A_998_115#_c_1540_n 0.0116326f $X=5.06 $Y=2.11 $X2=4.635
+ $Y2=1.37
cc_716 N_CK_c_760_n N_A_998_115#_c_1540_n 0.00613815f $X=5.455 $Y=2.11 $X2=4.635
+ $Y2=1.37
cc_717 N_CK_c_761_n N_A_998_115#_c_1540_n 0.020361f $X=5.31 $Y=2.11 $X2=4.635
+ $Y2=1.37
cc_718 N_CK_c_764_n N_A_998_115#_c_1540_n 6.61118e-19 $X=5.6 $Y=2.11 $X2=4.635
+ $Y2=1.37
cc_719 N_CK_c_751_n N_A_998_115#_c_1585_n 0.00150627f $X=5.455 $Y=2.285
+ $X2=5.045 $Y2=2.705
cc_720 N_CK_c_756_n N_A_998_115#_c_1585_n 0.00843004f $X=5.37 $Y=2.11 $X2=5.045
+ $Y2=2.705
cc_721 N_CK_c_757_n N_A_998_115#_c_1585_n 0.00323798f $X=5.06 $Y=2.11 $X2=5.045
+ $Y2=2.705
cc_722 N_CK_c_760_n N_A_998_115#_c_1585_n 0.00103871f $X=5.455 $Y=2.11 $X2=5.045
+ $Y2=2.705
cc_723 N_CK_c_761_n N_A_998_115#_c_1585_n 0.012754f $X=5.31 $Y=2.11 $X2=5.045
+ $Y2=2.705
cc_724 N_CK_c_764_n N_A_998_115#_c_1585_n 0.00146098f $X=5.6 $Y=2.11 $X2=5.045
+ $Y2=2.705
cc_725 N_CK_c_747_n N_A_998_115#_c_1541_n 0.00154744f $X=4.975 $Y=1.37 $X2=5.315
+ $Y2=1.37
cc_726 N_CK_c_748_n N_A_998_115#_c_1541_n 0.00321467f $X=4.975 $Y=1.205
+ $X2=5.315 $Y2=1.37
cc_727 N_CK_c_755_n N_A_998_115#_c_1541_n 0.0169532f $X=4.975 $Y=1.37 $X2=5.315
+ $Y2=1.37
cc_728 N_CK_c_756_n N_A_998_115#_c_1541_n 0.00114215f $X=5.37 $Y=2.11 $X2=5.315
+ $Y2=1.37
cc_729 N_CK_c_761_n N_A_998_115#_c_1541_n 2.84338e-19 $X=5.31 $Y=2.11 $X2=5.315
+ $Y2=1.37
cc_730 N_CK_c_752_n N_A_998_115#_c_1542_n 4.3075e-19 $X=6.385 $Y=1.28 $X2=7.13
+ $Y2=1.37
cc_731 N_CK_c_747_n N_A_998_115#_c_1544_n 0.00191034f $X=4.975 $Y=1.37 $X2=5.215
+ $Y2=0.755
cc_732 N_CK_c_748_n N_A_998_115#_c_1544_n 0.00389012f $X=4.975 $Y=1.205
+ $X2=5.215 $Y2=0.755
cc_733 N_CK_c_755_n N_A_998_115#_c_1544_n 9.01642e-19 $X=4.975 $Y=1.37 $X2=5.215
+ $Y2=0.755
cc_734 N_CK_c_747_n N_A_998_115#_c_1547_n 0.0042095f $X=4.975 $Y=1.37 $X2=5.18
+ $Y2=1.37
cc_735 N_CK_c_755_n N_A_998_115#_c_1547_n 0.0123759f $X=4.975 $Y=1.37 $X2=5.18
+ $Y2=1.37
cc_736 N_CK_c_756_n N_A_998_115#_c_1547_n 0.00195757f $X=5.37 $Y=2.11 $X2=5.18
+ $Y2=1.37
cc_737 N_CK_c_747_n N_A_998_115#_c_1548_n 3.88864e-19 $X=4.975 $Y=1.37 $X2=4.78
+ $Y2=1.37
cc_738 N_CK_c_755_n N_A_998_115#_c_1548_n 6.325e-19 $X=4.975 $Y=1.37 $X2=4.78
+ $Y2=1.37
cc_739 N_CK_c_761_n N_A_998_115#_c_1548_n 0.0128239f $X=5.31 $Y=2.11 $X2=4.78
+ $Y2=1.37
cc_740 N_CK_c_741_n N_A_998_115#_c_1549_n 0.00155926f $X=6.385 $Y=2.12 $X2=6.985
+ $Y2=1.37
cc_741 N_CK_c_752_n N_A_998_115#_c_1549_n 0.00331314f $X=6.385 $Y=1.28 $X2=6.985
+ $Y2=1.37
cc_742 CK N_A_998_115#_c_1549_n 0.00379778f $X=6.45 $Y=2.11 $X2=6.985 $Y2=1.37
cc_743 N_CK_c_747_n N_A_998_115#_c_1551_n 4.42421e-19 $X=4.975 $Y=1.37 $X2=5.44
+ $Y2=1.37
cc_744 N_CK_c_755_n N_A_998_115#_c_1551_n 0.00114522f $X=4.975 $Y=1.37 $X2=5.44
+ $Y2=1.37
cc_745 N_CK_c_756_n N_A_998_115#_c_1551_n 6.62932e-19 $X=5.37 $Y=2.11 $X2=5.44
+ $Y2=1.37
cc_746 N_CK_c_761_n N_A_998_115#_c_1551_n 0.00662656f $X=5.31 $Y=2.11 $X2=5.44
+ $Y2=1.37
cc_747 N_A_217_605#_c_1008_n N_A_618_89#_c_1127_n 0.00253253f $X=4.06 $Y=1.37
+ $X2=3.285 $Y2=1.745
cc_748 N_A_217_605#_c_1008_n N_A_618_89#_c_1128_n 0.00296105f $X=4.06 $Y=1.37
+ $X2=3.69 $Y2=1.82
cc_749 N_A_217_605#_c_994_n N_A_618_89#_M1017_g 0.114035f $X=4.2 $Y=2.285
+ $X2=3.765 $Y2=3.235
cc_750 N_A_217_605#_c_1005_n N_A_618_89#_M1017_g 0.00486364f $X=4.295 $Y=2.285
+ $X2=3.765 $Y2=3.235
cc_751 N_A_217_605#_c_992_n N_A_618_89#_c_1131_n 0.0342351f $X=4.2 $Y=1.37
+ $X2=4.84 $Y2=1.82
cc_752 N_A_217_605#_c_994_n N_A_618_89#_c_1131_n 0.0307748f $X=4.2 $Y=2.285
+ $X2=4.84 $Y2=1.82
cc_753 N_A_217_605#_c_1005_n N_A_618_89#_c_1131_n 0.0113171f $X=4.295 $Y=2.285
+ $X2=4.84 $Y2=1.82
cc_754 N_A_217_605#_c_1006_n N_A_618_89#_c_1131_n 8.69982e-19 $X=4.295 $Y=1.37
+ $X2=4.84 $Y2=1.82
cc_755 N_A_217_605#_c_1008_n N_A_618_89#_c_1131_n 0.00486036f $X=4.06 $Y=1.37
+ $X2=4.84 $Y2=1.82
cc_756 N_A_217_605#_c_1058_n N_A_618_89#_c_1131_n 4.12801e-19 $X=4.205 $Y=1.37
+ $X2=4.84 $Y2=1.82
cc_757 N_A_217_605#_c_993_n N_A_618_89#_M1003_g 0.110621f $X=4.48 $Y=2.285
+ $X2=4.915 $Y2=3.235
cc_758 N_A_217_605#_M1022_g N_A_998_115#_c_1540_n 9.36754e-19 $X=4.125 $Y=3.235
+ $X2=4.635 $Y2=1.37
cc_759 N_A_217_605#_c_990_n N_A_998_115#_c_1540_n 0.0061959f $X=4.48 $Y=1.37
+ $X2=4.635 $Y2=1.37
cc_760 N_A_217_605#_c_993_n N_A_998_115#_c_1540_n 0.00738718f $X=4.48 $Y=2.285
+ $X2=4.635 $Y2=1.37
cc_761 N_A_217_605#_M1025_g N_A_998_115#_c_1540_n 0.00190555f $X=4.555 $Y=0.835
+ $X2=4.635 $Y2=1.37
cc_762 N_A_217_605#_M1014_g N_A_998_115#_c_1540_n 0.00479454f $X=4.555 $Y=3.235
+ $X2=4.635 $Y2=1.37
cc_763 N_A_217_605#_c_1005_n N_A_998_115#_c_1540_n 0.0702347f $X=4.295 $Y=2.285
+ $X2=4.635 $Y2=1.37
cc_764 N_A_217_605#_c_1006_n N_A_998_115#_c_1540_n 0.0157315f $X=4.295 $Y=1.37
+ $X2=4.635 $Y2=1.37
cc_765 N_A_217_605#_c_1058_n N_A_998_115#_c_1540_n 4.18442e-19 $X=4.205 $Y=1.37
+ $X2=4.635 $Y2=1.37
cc_766 N_A_217_605#_M1022_g N_A_998_115#_c_1621_n 9.13132e-19 $X=4.125 $Y=3.235
+ $X2=4.72 $Y2=2.705
cc_767 N_A_217_605#_M1014_g N_A_998_115#_c_1621_n 0.0096885f $X=4.555 $Y=3.235
+ $X2=4.72 $Y2=2.705
cc_768 N_A_217_605#_c_990_n N_A_998_115#_c_1548_n 0.00229064f $X=4.48 $Y=1.37
+ $X2=4.78 $Y2=1.37
cc_769 N_A_217_605#_c_1006_n N_A_998_115#_c_1548_n 0.0012094f $X=4.295 $Y=1.37
+ $X2=4.78 $Y2=1.37
cc_770 N_A_217_605#_c_1058_n N_A_998_115#_c_1548_n 0.0241863f $X=4.205 $Y=1.37
+ $X2=4.78 $Y2=1.37
cc_771 N_A_618_89#_M1020_g N_A_1160_89#_c_1326_n 0.0575597f $X=5.515 $Y=0.835
+ $X2=5.89 $Y2=1.205
cc_772 N_A_618_89#_c_1142_n N_A_1160_89#_c_1330_n 0.00221914f $X=6.52 $Y=0.755
+ $X2=5.89 $Y2=1.365
cc_773 N_A_618_89#_c_1141_n N_A_1160_89#_c_1333_n 7.17123e-19 $X=5.455 $Y=1.725
+ $X2=5.965 $Y2=1.77
cc_774 N_A_618_89#_c_1148_n N_A_1160_89#_c_1333_n 9.21617e-19 $X=6.52 $Y=1.725
+ $X2=5.965 $Y2=1.77
cc_775 N_A_618_89#_c_1149_n N_A_1160_89#_c_1333_n 0.00307203f $X=6.215 $Y=1.74
+ $X2=5.965 $Y2=1.77
cc_776 N_A_618_89#_c_1150_n N_A_1160_89#_c_1333_n 9.45235e-19 $X=6.36 $Y=1.74
+ $X2=5.965 $Y2=1.77
cc_777 N_A_618_89#_M1020_g N_A_1160_89#_c_1335_n 0.00905991f $X=5.515 $Y=0.835
+ $X2=5.965 $Y2=1.605
cc_778 N_A_618_89#_c_1140_n N_A_1160_89#_c_1335_n 0.0260042f $X=5.455 $Y=1.725
+ $X2=5.965 $Y2=1.605
cc_779 N_A_618_89#_c_1140_n N_A_1160_89#_c_1341_n 0.00126849f $X=5.455 $Y=1.725
+ $X2=5.935 $Y2=2.025
cc_780 N_A_618_89#_c_1141_n N_A_1160_89#_c_1341_n 0.00810099f $X=5.455 $Y=1.725
+ $X2=5.935 $Y2=2.025
cc_781 N_A_618_89#_c_1142_n N_A_1160_89#_c_1341_n 6.86732e-19 $X=6.52 $Y=0.755
+ $X2=5.935 $Y2=2.025
cc_782 N_A_618_89#_c_1147_n N_A_1160_89#_c_1341_n 0.00444172f $X=6.795 $Y=2.62
+ $X2=5.935 $Y2=2.025
cc_783 N_A_618_89#_c_1148_n N_A_1160_89#_c_1341_n 0.00950295f $X=6.52 $Y=1.725
+ $X2=5.935 $Y2=2.025
cc_784 N_A_618_89#_c_1149_n N_A_1160_89#_c_1341_n 0.0125852f $X=6.215 $Y=1.74
+ $X2=5.935 $Y2=2.025
cc_785 N_A_618_89#_c_1241_n N_A_1160_89#_c_1341_n 0.00127809f $X=5.6 $Y=1.74
+ $X2=5.935 $Y2=2.025
cc_786 N_A_618_89#_c_1150_n N_A_1160_89#_c_1341_n 0.00194798f $X=6.36 $Y=1.74
+ $X2=5.935 $Y2=2.025
cc_787 N_A_618_89#_c_1157_n N_A_1160_89#_c_1368_n 0.0313767f $X=6.52 $Y=2.955
+ $X2=7.04 $Y2=3.275
cc_788 N_A_618_89#_c_1157_n N_A_1160_89#_c_1372_n 0.00815518f $X=6.52 $Y=2.955
+ $X2=7.125 $Y2=3.045
cc_789 N_A_618_89#_c_1148_n N_A_1160_89#_c_1344_n 0.00106098f $X=6.52 $Y=1.725
+ $X2=7.47 $Y2=0.74
cc_790 N_A_618_89#_c_1147_n N_A_1160_89#_c_1347_n 0.0178263f $X=6.795 $Y=2.62
+ $X2=7.47 $Y2=2.96
cc_791 N_A_618_89#_c_1161_n N_A_1160_89#_c_1347_n 0.00644034f $X=6.795 $Y=2.705
+ $X2=7.47 $Y2=2.96
cc_792 N_A_618_89#_c_1148_n N_A_1160_89#_c_1349_n 0.00398388f $X=6.52 $Y=1.725
+ $X2=7.47 $Y2=1.74
cc_793 N_A_618_89#_c_1147_n N_A_1160_89#_c_1350_n 0.013021f $X=6.795 $Y=2.62
+ $X2=6.735 $Y2=2.48
cc_794 N_A_618_89#_c_1148_n N_A_1160_89#_c_1350_n 0.00366675f $X=6.52 $Y=1.725
+ $X2=6.735 $Y2=2.48
cc_795 N_A_618_89#_c_1161_n N_A_1160_89#_c_1350_n 0.0134869f $X=6.795 $Y=2.705
+ $X2=6.735 $Y2=2.48
cc_796 N_A_618_89#_c_1147_n N_A_1160_89#_c_1352_n 0.0215237f $X=6.795 $Y=2.62
+ $X2=6.825 $Y2=2.395
cc_797 N_A_618_89#_c_1148_n N_A_1160_89#_c_1353_n 0.0109407f $X=6.52 $Y=1.725
+ $X2=6.915 $Y2=1.737
cc_798 N_A_618_89#_c_1150_n N_A_1160_89#_c_1353_n 0.0166008f $X=6.36 $Y=1.74
+ $X2=6.915 $Y2=1.737
cc_799 N_A_618_89#_c_1142_n N_A_998_115#_M1012_g 0.00559858f $X=6.52 $Y=0.755
+ $X2=7.255 $Y2=0.755
cc_800 N_A_618_89#_c_1142_n N_A_998_115#_M1006_g 0.0013415f $X=6.52 $Y=0.755
+ $X2=7.255 $Y2=3.445
cc_801 N_A_618_89#_c_1157_n N_A_998_115#_M1006_g 0.00441825f $X=6.52 $Y=2.955
+ $X2=7.255 $Y2=3.445
cc_802 N_A_618_89#_c_1147_n N_A_998_115#_M1006_g 0.00857372f $X=6.795 $Y=2.62
+ $X2=7.255 $Y2=3.445
cc_803 N_A_618_89#_c_1148_n N_A_998_115#_M1006_g 0.00170265f $X=6.52 $Y=1.725
+ $X2=7.255 $Y2=3.445
cc_804 N_A_618_89#_c_1161_n N_A_998_115#_M1006_g 0.00343288f $X=6.795 $Y=2.705
+ $X2=7.255 $Y2=3.445
cc_805 N_A_618_89#_c_1142_n N_A_998_115#_c_1538_n 0.00208762f $X=6.52 $Y=0.755
+ $X2=7.13 $Y2=1.37
cc_806 N_A_618_89#_c_1131_n N_A_998_115#_c_1540_n 0.0123066f $X=4.84 $Y=1.82
+ $X2=4.635 $Y2=1.37
cc_807 N_A_618_89#_M1003_g N_A_998_115#_c_1540_n 0.0111407f $X=4.915 $Y=3.235
+ $X2=4.635 $Y2=1.37
cc_808 N_A_618_89#_M1003_g N_A_998_115#_c_1585_n 0.0162544f $X=4.915 $Y=3.235
+ $X2=5.045 $Y2=2.705
cc_809 N_A_618_89#_c_1140_n N_A_998_115#_c_1541_n 0.00206196f $X=5.455 $Y=1.725
+ $X2=5.315 $Y2=1.37
cc_810 N_A_618_89#_c_1141_n N_A_998_115#_c_1541_n 0.00758189f $X=5.455 $Y=1.725
+ $X2=5.315 $Y2=1.37
cc_811 N_A_618_89#_c_1142_n N_A_998_115#_c_1542_n 0.00866447f $X=6.52 $Y=0.755
+ $X2=7.13 $Y2=1.37
cc_812 N_A_618_89#_M1020_g N_A_998_115#_c_1544_n 0.0131134f $X=5.515 $Y=0.835
+ $X2=5.215 $Y2=0.755
cc_813 N_A_618_89#_c_1131_n N_A_998_115#_c_1547_n 0.00156696f $X=4.84 $Y=1.82
+ $X2=5.18 $Y2=1.37
cc_814 N_A_618_89#_c_1133_n N_A_998_115#_c_1547_n 0.00141359f $X=5.32 $Y=1.82
+ $X2=5.18 $Y2=1.37
cc_815 N_A_618_89#_c_1139_n N_A_998_115#_c_1547_n 5.19983e-19 $X=4.915 $Y=1.82
+ $X2=5.18 $Y2=1.37
cc_816 N_A_618_89#_c_1131_n N_A_998_115#_c_1548_n 0.00120486f $X=4.84 $Y=1.82
+ $X2=4.78 $Y2=1.37
cc_817 N_A_618_89#_M1020_g N_A_998_115#_c_1549_n 0.00393577f $X=5.515 $Y=0.835
+ $X2=6.985 $Y2=1.37
cc_818 N_A_618_89#_c_1140_n N_A_998_115#_c_1549_n 5.08054e-19 $X=5.455 $Y=1.725
+ $X2=6.985 $Y2=1.37
cc_819 N_A_618_89#_c_1141_n N_A_998_115#_c_1549_n 0.00283556f $X=5.455 $Y=1.725
+ $X2=6.985 $Y2=1.37
cc_820 N_A_618_89#_c_1142_n N_A_998_115#_c_1549_n 0.0174175f $X=6.52 $Y=0.755
+ $X2=6.985 $Y2=1.37
cc_821 N_A_618_89#_c_1148_n N_A_998_115#_c_1549_n 0.013349f $X=6.52 $Y=1.725
+ $X2=6.985 $Y2=1.37
cc_822 N_A_618_89#_c_1149_n N_A_998_115#_c_1549_n 0.0512581f $X=6.215 $Y=1.74
+ $X2=6.985 $Y2=1.37
cc_823 N_A_618_89#_c_1241_n N_A_998_115#_c_1549_n 0.0139023f $X=5.6 $Y=1.74
+ $X2=6.985 $Y2=1.37
cc_824 N_A_618_89#_c_1150_n N_A_998_115#_c_1549_n 0.0265578f $X=6.36 $Y=1.74
+ $X2=6.985 $Y2=1.37
cc_825 N_A_618_89#_c_1133_n N_A_998_115#_c_1551_n 6.94944e-19 $X=5.32 $Y=1.82
+ $X2=5.44 $Y2=1.37
cc_826 N_A_618_89#_M1020_g N_A_998_115#_c_1551_n 0.00225742f $X=5.515 $Y=0.835
+ $X2=5.44 $Y2=1.37
cc_827 N_A_618_89#_c_1140_n N_A_998_115#_c_1551_n 0.0020361f $X=5.455 $Y=1.725
+ $X2=5.44 $Y2=1.37
cc_828 N_A_618_89#_c_1141_n N_A_998_115#_c_1551_n 0.0012656f $X=5.455 $Y=1.725
+ $X2=5.44 $Y2=1.37
cc_829 N_A_618_89#_c_1241_n N_A_998_115#_c_1551_n 0.0127467f $X=5.6 $Y=1.74
+ $X2=5.44 $Y2=1.37
cc_830 N_A_618_89#_c_1142_n N_A_998_115#_c_1552_n 0.00153931f $X=6.52 $Y=0.755
+ $X2=7.13 $Y2=1.37
cc_831 N_A_1160_89#_c_1344_n N_A_998_115#_M1012_g 0.0108232f $X=7.47 $Y=0.74
+ $X2=7.255 $Y2=0.755
cc_832 N_A_1160_89#_c_1371_n N_A_998_115#_M1006_g 0.0193327f $X=7.385 $Y=3.045
+ $X2=7.255 $Y2=3.445
cc_833 N_A_1160_89#_c_1347_n N_A_998_115#_M1006_g 0.0138402f $X=7.47 $Y=2.96
+ $X2=7.255 $Y2=3.445
cc_834 N_A_1160_89#_c_1349_n N_A_998_115#_M1006_g 0.00169596f $X=7.47 $Y=1.74
+ $X2=7.255 $Y2=3.445
cc_835 N_A_1160_89#_c_1352_n N_A_998_115#_M1006_g 0.0124124f $X=6.825 $Y=2.395
+ $X2=7.255 $Y2=3.445
cc_836 N_A_1160_89#_c_1355_n N_A_998_115#_M1006_g 0.0125592f $X=8.375 $Y=1.74
+ $X2=7.255 $Y2=3.445
cc_837 N_A_1160_89#_c_1355_n N_A_998_115#_c_1538_n 7.95399e-19 $X=8.375 $Y=1.74
+ $X2=7.13 $Y2=1.37
cc_838 N_A_1160_89#_c_1344_n N_A_998_115#_c_1542_n 0.0213712f $X=7.47 $Y=0.74
+ $X2=7.13 $Y2=1.37
cc_839 N_A_1160_89#_c_1355_n N_A_998_115#_c_1542_n 0.00454041f $X=8.375 $Y=1.74
+ $X2=7.13 $Y2=1.37
cc_840 N_A_1160_89#_c_1330_n N_A_998_115#_c_1549_n 0.00346468f $X=5.89 $Y=1.365
+ $X2=6.985 $Y2=1.37
cc_841 N_A_1160_89#_c_1333_n N_A_998_115#_c_1549_n 7.74479e-19 $X=5.965 $Y=1.77
+ $X2=6.985 $Y2=1.37
cc_842 N_A_1160_89#_c_1335_n N_A_998_115#_c_1549_n 0.00274919f $X=5.965 $Y=1.605
+ $X2=6.985 $Y2=1.37
cc_843 N_A_1160_89#_c_1341_n N_A_998_115#_c_1549_n 0.00439053f $X=5.935 $Y=2.025
+ $X2=6.985 $Y2=1.37
cc_844 N_A_1160_89#_c_1353_n N_A_998_115#_c_1549_n 0.0218319f $X=6.915 $Y=1.737
+ $X2=6.985 $Y2=1.37
cc_845 N_A_1160_89#_c_1344_n N_A_998_115#_c_1552_n 0.0027677f $X=7.47 $Y=0.74
+ $X2=7.13 $Y2=1.37
cc_846 N_A_1160_89#_c_1355_n N_A_998_115#_c_1552_n 0.0263691f $X=8.375 $Y=1.74
+ $X2=7.13 $Y2=1.37
cc_847 N_A_1160_89#_M1016_g N_QN_M1008_g 0.0210474f $X=8.635 $Y=0.755 $X2=9.065
+ $Y2=0.755
cc_848 N_A_1160_89#_c_1337_n N_QN_M1008_g 0.0152125f $X=8.522 $Y=1.575 $X2=9.065
+ $Y2=0.755
cc_849 N_A_1160_89#_c_1348_n N_QN_M1008_g 3.6337e-19 $X=8.52 $Y=1.74 $X2=9.065
+ $Y2=0.755
cc_850 N_A_1160_89#_c_1339_n N_QN_M1001_g 0.0102953f $X=8.61 $Y=2.375 $X2=9.065
+ $Y2=3.445
cc_851 N_A_1160_89#_c_1340_n N_QN_M1001_g 0.0339596f $X=8.61 $Y=2.525 $X2=9.065
+ $Y2=3.445
cc_852 N_A_1160_89#_c_1336_n N_QN_c_1680_n 0.0211392f $X=8.52 $Y=1.74 $X2=9.005
+ $Y2=1.915
cc_853 N_A_1160_89#_c_1348_n N_QN_c_1680_n 5.0648e-19 $X=8.52 $Y=1.74 $X2=9.005
+ $Y2=1.915
cc_854 N_A_1160_89#_c_1354_n N_QN_c_1680_n 4.60229e-19 $X=8.52 $Y=1.74 $X2=9.005
+ $Y2=1.915
cc_855 N_A_1160_89#_M1016_g N_QN_c_1681_n 0.00760341f $X=8.635 $Y=0.755 $X2=8.42
+ $Y2=0.74
cc_856 N_A_1160_89#_c_1338_n N_QN_c_1681_n 0.00327645f $X=8.61 $Y=1.32 $X2=8.42
+ $Y2=0.74
cc_857 N_A_1160_89#_M1011_g N_QN_c_1685_n 0.0164234f $X=8.635 $Y=3.445 $X2=8.42
+ $Y2=2.48
cc_858 N_A_1160_89#_c_1339_n N_QN_c_1685_n 0.00567875f $X=8.61 $Y=2.375 $X2=8.42
+ $Y2=2.48
cc_859 N_A_1160_89#_c_1337_n N_QN_c_1686_n 0.00784613f $X=8.522 $Y=1.575
+ $X2=8.92 $Y2=1.37
cc_860 N_A_1160_89#_c_1338_n N_QN_c_1686_n 0.0108281f $X=8.61 $Y=1.32 $X2=8.92
+ $Y2=1.37
cc_861 N_A_1160_89#_c_1348_n N_QN_c_1686_n 0.0093039f $X=8.52 $Y=1.74 $X2=8.92
+ $Y2=1.37
cc_862 N_A_1160_89#_c_1354_n N_QN_c_1686_n 0.0037949f $X=8.52 $Y=1.74 $X2=8.92
+ $Y2=1.37
cc_863 N_A_1160_89#_c_1336_n N_QN_c_1688_n 0.00303508f $X=8.52 $Y=1.74 $X2=8.505
+ $Y2=1.37
cc_864 N_A_1160_89#_c_1348_n N_QN_c_1688_n 0.0101631f $X=8.52 $Y=1.74 $X2=8.505
+ $Y2=1.37
cc_865 N_A_1160_89#_c_1354_n N_QN_c_1688_n 0.00331526f $X=8.52 $Y=1.74 $X2=8.505
+ $Y2=1.37
cc_866 N_A_1160_89#_c_1355_n N_QN_c_1688_n 0.00105631f $X=8.375 $Y=1.74
+ $X2=8.505 $Y2=1.37
cc_867 N_A_1160_89#_c_1339_n N_QN_c_1689_n 0.0159847f $X=8.61 $Y=2.375 $X2=8.92
+ $Y2=2.285
cc_868 N_A_1160_89#_c_1340_n N_QN_c_1689_n 0.00248624f $X=8.61 $Y=2.525 $X2=8.92
+ $Y2=2.285
cc_869 N_A_1160_89#_c_1348_n N_QN_c_1689_n 0.0046698f $X=8.52 $Y=1.74 $X2=8.92
+ $Y2=2.285
cc_870 N_A_1160_89#_c_1354_n N_QN_c_1689_n 0.00258299f $X=8.52 $Y=1.74 $X2=8.92
+ $Y2=2.285
cc_871 N_A_1160_89#_c_1336_n N_QN_c_1690_n 0.00271474f $X=8.52 $Y=1.74 $X2=8.505
+ $Y2=2.285
cc_872 N_A_1160_89#_c_1348_n N_QN_c_1690_n 0.00515207f $X=8.52 $Y=1.74 $X2=8.505
+ $Y2=2.285
cc_873 N_A_1160_89#_c_1354_n N_QN_c_1690_n 0.00139444f $X=8.52 $Y=1.74 $X2=8.505
+ $Y2=2.285
cc_874 N_A_1160_89#_c_1355_n N_QN_c_1690_n 4.39196e-19 $X=8.375 $Y=1.74
+ $X2=8.505 $Y2=2.285
cc_875 N_A_1160_89#_c_1336_n N_QN_c_1691_n 0.0019182f $X=8.52 $Y=1.74 $X2=9.005
+ $Y2=1.915
cc_876 N_A_1160_89#_c_1337_n N_QN_c_1691_n 0.00380475f $X=8.522 $Y=1.575
+ $X2=9.005 $Y2=1.915
cc_877 N_A_1160_89#_c_1339_n N_QN_c_1691_n 0.00226435f $X=8.61 $Y=2.375
+ $X2=9.005 $Y2=1.915
cc_878 N_A_1160_89#_c_1348_n N_QN_c_1691_n 0.00978463f $X=8.52 $Y=1.74 $X2=9.005
+ $Y2=1.915
cc_879 N_A_1160_89#_c_1354_n N_QN_c_1691_n 0.00377829f $X=8.52 $Y=1.74 $X2=9.005
+ $Y2=1.915
cc_880 N_A_1160_89#_M1011_g QN 0.00233857f $X=8.635 $Y=3.445 $X2=8.425 $Y2=2.48
cc_881 N_A_1160_89#_c_1340_n QN 0.00508004f $X=8.61 $Y=2.525 $X2=8.425 $Y2=2.48
cc_882 N_A_1160_89#_c_1347_n QN 0.00513409f $X=7.47 $Y=2.96 $X2=8.425 $Y2=2.48
cc_883 N_A_1160_89#_c_1348_n QN 0.00286804f $X=8.52 $Y=1.74 $X2=8.425 $Y2=2.48
cc_884 N_A_1160_89#_c_1354_n QN 0.00881422f $X=8.52 $Y=1.74 $X2=8.425 $Y2=2.48
cc_885 N_A_1160_89#_c_1355_n QN 0.00487781f $X=8.375 $Y=1.74 $X2=8.425 $Y2=2.48
cc_886 N_A_1160_89#_c_1371_n A_1466_605# 0.00433061f $X=7.385 $Y=3.045 $X2=7.33
+ $Y2=3.025
cc_887 N_A_998_115#_c_1585_n A_926_521# 0.00342591f $X=5.045 $Y=2.705 $X2=4.63
+ $Y2=2.605
cc_888 N_A_998_115#_c_1621_n A_926_521# 0.00144354f $X=4.72 $Y=2.705 $X2=4.63
+ $Y2=2.605
cc_889 N_QN_M1008_g N_Q_c_1771_n 5.62519e-19 $X=9.065 $Y=0.755 $X2=9.28 $Y2=0.74
cc_890 N_QN_M1001_g N_Q_c_1775_n 0.00409136f $X=9.065 $Y=3.445 $X2=9.28
+ $Y2=3.265
cc_891 N_QN_M1008_g N_Q_c_1773_n 0.0383548f $X=9.065 $Y=0.755 $X2=9.395 $Y2=2.68
cc_892 N_QN_c_1686_n N_Q_c_1773_n 0.0111776f $X=8.92 $Y=1.37 $X2=9.395 $Y2=2.68
cc_893 N_QN_c_1689_n N_Q_c_1773_n 0.0111776f $X=8.92 $Y=2.285 $X2=9.395 $Y2=2.68
cc_894 N_QN_c_1691_n N_Q_c_1773_n 0.0438362f $X=9.005 $Y=1.915 $X2=9.395
+ $Y2=2.68
cc_895 N_QN_M1008_g N_Q_c_1774_n 0.00695117f $X=9.065 $Y=0.755 $X2=9.395
+ $Y2=1.035
cc_896 N_QN_M1001_g N_Q_c_1780_n 0.00614447f $X=9.065 $Y=3.445 $X2=9.28
+ $Y2=2.807
cc_897 N_QN_M1001_g Q 0.0131514f $X=9.065 $Y=3.445 $X2=9.275 $Y2=2.85
cc_898 N_QN_c_1689_n Q 0.00245821f $X=8.92 $Y=2.285 $X2=9.275 $Y2=2.85
