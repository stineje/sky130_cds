* File: sky130_osu_sc_12T_ms__or2_2.pex.spice
* Created: Fri Nov 12 15:26:11 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__OR2_2%GND 1 2 3 31 35 37 44 46 54 64 66
r44 64 66 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r45 52 54 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r46 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r47 46 52 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.305
r48 42 60 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r49 42 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r50 37 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r51 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r52 31 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r53 31 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r54 31 33 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r55 31 38 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r56 31 46 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r57 31 47 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r58 31 37 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r59 31 38 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r60 3 54 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84 $Y=0.575
+ $X2=1.98 $Y2=0.755
r61 2 44 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98 $Y=0.575
+ $X2=1.12 $Y2=0.755
r62 1 35 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_2%VDD 1 2 21 23 32 34 41 47 51
r30 47 51 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.7 $Y2=4.287
r31 41 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r32 39 44 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135 $X2=1.98
+ $Y2=3.635
r33 37 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=4.25 $X2=1.7
+ $Y2=4.25
r34 35 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r35 35 37 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r36 34 39 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.135
r37 34 37 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r38 30 45 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r39 30 32 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135 $X2=1.12
+ $Y2=3.635
r40 25 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r41 25 29 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r42 23 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r43 23 29 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r44 21 37 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r45 21 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r46 21 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r47 2 44 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r48 2 41 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r49 1 32 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_2%B 3 7 12 15 21
r28 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.48
r29 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.195
+ $X2=0.27 $Y2=2.48
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.195 $X2=0.27 $Y2=2.195
r31 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.195
+ $X2=0.475 $Y2=2.195
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=2.195
r33 5 7 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.475 $Y=2.36
+ $X2=0.475 $Y2=3.235
r34 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.03
+ $X2=0.475 $Y2=2.195
r35 1 3 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.475 $Y=2.03
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_2%A 3 7 10 14 20
c44 7 0 1.37149e-19 $X=0.905 $Y=3.235
r45 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.85
+ $X2=0.95 $Y2=2.85
r46 14 17 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=2.85
r47 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.905 $X2=0.95 $Y2=1.905
r48 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=2.07
r49 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.905
+ $X2=0.95 $Y2=1.74
r50 7 12 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.07
r51 3 11 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=0.905 $Y=0.835
+ $X2=0.905 $Y2=1.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_2%A_27_521# 1 3 11 13 15 17 18 22 24 26 27
+ 31 35 37 38 40 43 47 49
r87 45 49 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.455
+ $X2=0.65 $Y2=1.455
r88 45 47 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.455
+ $X2=1.43 $Y2=1.455
r89 41 49 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.65 $Y2=1.455
r90 41 43 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.69 $Y2=0.755
r91 39 49 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.65 $Y2=1.455
r92 39 40 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.54
+ $X2=0.61 $Y2=3.065
r93 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.15
+ $X2=0.61 $Y2=3.065
r94 37 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.15
+ $X2=0.345 $Y2=3.15
r95 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.235
+ $X2=0.345 $Y2=3.15
r96 33 35 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.26 $Y=3.235 $X2=0.26
+ $Y2=3.295
r97 31 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.455 $X2=1.43 $Y2=1.455
r98 29 31 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.455 $X2=1.43
+ $Y2=1.455
r99 28 29 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.455
+ $X2=1.37 $Y2=1.455
r100 24 26 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r101 20 31 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.43 $Y2=1.455
r102 20 22 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=0.835
r103 19 27 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.405
+ $X2=1.352 $Y2=2.405
r104 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.48
r105 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.445 $Y2=2.405
r106 17 27 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.33
+ $X2=1.352 $Y2=2.405
r107 16 29 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=1.455
r108 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.62
+ $X2=1.37 $Y2=2.33
r109 13 27 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.352 $Y2=2.405
r110 13 15 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r111 9 28 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=1.455
r112 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.835
r113 3 35 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.295
r114 1 43 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__OR2_2%Y 1 3 10 16 26 29 32
c42 16 0 1.37149e-19 $X=1.55 $Y=2.11
r43 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=2.11
r44 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=1.995
+ $X2=1.55 $Y2=1.74
r45 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r46 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1.74
r47 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r48 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.11
r49 16 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.55 $Y=2.11
+ $X2=1.55 $Y2=2.955
r50 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r51 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r52 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r53 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r54 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41 $Y=0.575
+ $X2=1.55 $Y2=0.755
.ends

