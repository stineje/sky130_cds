* File: sky130_osu_sc_18T_ls__aoi21_l.pex.spice
* Created: Thu Oct 29 17:34:19 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%GND 1 2 15 19 23 29 31 34
c40 15 0 6.36774e-20 $X=-0.045 $Y=0
r41 31 34 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r42 21 29 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.54 $Y=0.305
+ $X2=1.455 $Y2=0.152
r43 21 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.54 $Y=0.305
+ $X2=1.54 $Y2=0.825
r44 17 19 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r45 15 29 16.4365 $w=3.03e-07 $l=4.35e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.455 $Y2=0.152
r46 15 25 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r47 15 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r48 15 17 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r49 15 25 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r50 2 23 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.825
r51 1 19 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%VDD 1 10 12 18 25 28 32
r26 28 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r27 25 28 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r28 22 32 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507 $X2=1.02
+ $Y2=6.507
r29 22 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r30 18 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=4.475
+ $X2=0.69 $Y2=5.835
r31 16 23 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r32 16 21 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r33 12 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r34 12 14 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r35 10 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r36 10 14 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r37 1 21 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r38 1 18 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%A0 2 3 5 8 12 15 22 24
c37 8 0 6.36774e-20 $X=0.475 $Y=4.585
r38 23 24 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.765
+ $X2=0.475 $Y2=2.765
r39 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.765 $X2=0.385 $Y2=2.765
r40 19 23 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.765
+ $X2=0.385 $Y2=2.765
r41 17 22 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.385 $Y2=2.765
r42 15 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=3.33
+ $X2=0.385 $Y2=3.33
r43 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.77
+ $X2=0.475 $Y2=1.77
r44 6 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=2.765
r45 6 8 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=4.585
r46 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.69 $X2=0.475
+ $Y2=1.77
r47 3 5 197.62 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.475 $Y=1.69
+ $X2=0.475 $Y2=1.075
r48 2 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.63
+ $X2=0.295 $Y2=2.765
r49 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.85 $X2=0.295
+ $Y2=1.77
r50 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.85
+ $X2=0.295 $Y2=2.63
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%A1 3 7 13 14 17 19
c50 17 0 1.38614e-19 $X=0.725 $Y=2.96
r51 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.96
+ $X2=0.725 $Y2=2.96
r52 14 23 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=2.255
+ $X2=0.825 $Y2=2.42
r53 14 22 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=2.255
+ $X2=0.825 $Y2=2.09
r54 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=2.255 $X2=0.815 $Y2=2.255
r55 10 19 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.725 $Y=2.42
+ $X2=0.725 $Y2=2.96
r56 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.725 $Y=2.255
+ $X2=0.815 $Y2=2.255
r57 9 10 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=2.255
+ $X2=0.725 $Y2=2.42
r58 7 23 1110.14 $w=1.5e-07 $l=2.165e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.42
r59 3 22 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.09
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%B0 3 7 10 13 15 17 22 24 27
c53 7 0 1.38614e-19 $X=1.335 $Y=4.585
r54 22 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.59
+ $X2=1.165 $Y2=2.59
r55 20 24 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.165 $Y=1.945
+ $X2=1.165 $Y2=2.59
r56 18 27 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.53 $Y=1.86 $X2=1.47
+ $Y2=1.86
r57 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.53
+ $Y=1.86 $X2=1.53 $Y2=1.86
r58 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.25 $Y=1.86
+ $X2=1.165 $Y2=1.945
r59 15 17 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.25 $Y=1.86
+ $X2=1.53 $Y2=1.86
r60 11 13 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.335 $Y=2.82
+ $X2=1.47 $Y2=2.82
r61 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=2.745
+ $X2=1.47 $Y2=2.82
r62 9 27 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=2.025
+ $X2=1.47 $Y2=1.86
r63 9 10 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.47 $Y=2.025
+ $X2=1.47 $Y2=2.745
r64 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.895
+ $X2=1.335 $Y2=2.82
r65 5 7 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=1.335 $Y=2.895
+ $X2=1.335 $Y2=4.585
r66 1 27 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.325 $Y=1.695
+ $X2=1.47 $Y2=1.86
r67 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.325 $Y=1.695
+ $X2=1.325 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%A_27_617# 1 2 9 13 14 17
r16 17 19 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=5.835
r17 15 17 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=4.055 $X2=1.12
+ $Y2=4.135
r18 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.97
+ $X2=1.12 $Y2=4.055
r19 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.97
+ $X2=0.345 $Y2=3.97
r20 9 11 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r21 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=4.055
+ $X2=0.345 $Y2=3.97
r22 7 9 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=4.055 $X2=0.26
+ $Y2=4.135
r23 2 19 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r24 2 17 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=4.135
r25 1 11 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r26 1 9 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI21_L%Y 1 2 7 8 12 19 20 23
r46 30 32 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.55 $Y=3.795
+ $X2=1.55 $Y2=5.835
r47 20 30 102.754 $w=1.68e-07 $l=1.575e-06 $layer=LI1_cond $X=1.55 $Y=2.22
+ $X2=1.55 $Y2=3.795
r48 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.22
+ $X2=1.55 $Y2=2.22
r49 16 23 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.05 $Y=1.48
+ $X2=1.05 $Y2=0.825
r50 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.05 $Y=1.48
+ $X2=1.05 $Y2=1.48
r51 10 19 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.105
+ $X2=1.55 $Y2=2.22
r52 10 12 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.55 $Y=2.105
+ $X2=1.55 $Y2=2.07
r53 9 12 0.486256 $w=1.7e-07 $l=5.05e-07 $layer=MET1_cond $X=1.55 $Y=1.565
+ $X2=1.55 $Y2=2.07
r54 8 15 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.195 $Y=1.48
+ $X2=1.05 $Y2=1.48
r55 7 9 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.465 $Y=1.48
+ $X2=1.55 $Y2=1.565
r56 7 8 0.259978 $w=1.7e-07 $l=2.7e-07 $layer=MET1_cond $X=1.465 $Y=1.48
+ $X2=1.195 $Y2=1.48
r57 2 32 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r58 2 30 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.795
r59 1 23 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

