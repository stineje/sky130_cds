* File: sky130_osu_sc_15T_ls__buf_8.spice
* Created: Fri Nov 12 14:55:15 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__buf_8.pex.spice"
.subckt sky130_osu_sc_15T_ls__buf_8  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_A_M1006_g N_A_27_115#_M1006_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1006_d N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1000_d N_A_27_115#_M1002_g N_GND_M1002_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_A_27_115#_M1007_g N_GND_M1002_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1007_d N_A_27_115#_M1010_g N_GND_M1010_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A_27_115#_M1011_g N_GND_M1010_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.3 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1011_d N_A_27_115#_M1012_g N_GND_M1012_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1014_d N_A_27_115#_M1014_g N_GND_M1012_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1014_d N_A_27_115#_M1016_g N_GND_M1016_s N_GND_M1006_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75003.6 A=0.3 P=4.3 MULT=1
MM1003 N_VDD_M1001_d N_A_27_115#_M1003_g N_Y_M1003_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75003.2 A=0.3 P=4.3 MULT=1
MM1004 N_VDD_M1004_d N_A_27_115#_M1004_g N_Y_M1003_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75001
+ SB=75002.8 A=0.3 P=4.3 MULT=1
MM1005 N_VDD_M1004_d N_A_27_115#_M1005_g N_Y_M1005_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001.5 SB=75002.3 A=0.3 P=4.3 MULT=1
MM1008 N_VDD_M1008_d N_A_27_115#_M1008_g N_Y_M1005_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001.9 SB=75001.9 A=0.3 P=4.3 MULT=1
MM1009 N_VDD_M1008_d N_A_27_115#_M1009_g N_Y_M1009_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.3 SB=75001.5 A=0.3 P=4.3 MULT=1
MM1013 N_VDD_M1013_d N_A_27_115#_M1013_g N_Y_M1009_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.8 SB=75001 A=0.3 P=4.3 MULT=1
MM1015 N_VDD_M1013_d N_A_27_115#_M1015_g N_Y_M1015_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.28 PD=2.28 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1017 N_VDD_M1017_d N_A_27_115#_M1017_g N_Y_M1015_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.6 SB=75000.2 A=0.3 P=4.3 MULT=1
DX18_noxref N_GND_M1006_b N_VDD_M1001_b NWDIODE A=13.4667 P=15.03
pX19_noxref noxref_6 A A PROBETYPE=1
pX20_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__buf_8.pxi.spice"
*
.ends
*
*
