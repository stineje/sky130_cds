* File: sky130_osu_sc_15T_ms__aoi22_l.pxi.spice
* Created: Fri Nov 12 14:41:13 2021
* 
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%GND N_GND_M1005_s N_GND_M1007_d N_GND_M1005_b
+ N_GND_c_3_p N_GND_c_4_p N_GND_c_27_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_15T_MS__AOI22_L%GND
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%VDD N_VDD_M1006_d N_VDD_M1006_b N_VDD_c_47_p
+ N_VDD_c_48_p N_VDD_c_54_p VDD N_VDD_c_49_p
+ PM_SKY130_OSU_SC_15T_MS__AOI22_L%VDD
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%A0 N_A0_c_77_n N_A0_c_78_n N_A0_M1005_g
+ N_A0_M1006_g N_A0_c_82_n N_A0_c_84_n N_A0_c_85_n A0
+ PM_SKY130_OSU_SC_15T_MS__AOI22_L%A0
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%A1 N_A1_M1002_g N_A1_c_115_n N_A1_M1003_g
+ N_A1_c_117_n A1 PM_SKY130_OSU_SC_15T_MS__AOI22_L%A1
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%B0 N_B0_M1001_g N_B0_M1004_g N_B0_c_160_n
+ N_B0_c_161_n N_B0_c_162_n B0 PM_SKY130_OSU_SC_15T_MS__AOI22_L%B0
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%B1 N_B1_M1007_g N_B1_M1000_g N_B1_c_204_n
+ N_B1_c_206_n B1 PM_SKY130_OSU_SC_15T_MS__AOI22_L%B1
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%A_27_565# N_A_27_565#_M1006_s
+ N_A_27_565#_M1003_d N_A_27_565#_M1000_d N_A_27_565#_c_240_n
+ N_A_27_565#_c_226_n N_A_27_565#_c_229_n N_A_27_565#_c_231_n
+ N_A_27_565#_c_234_n PM_SKY130_OSU_SC_15T_MS__AOI22_L%A_27_565#
x_PM_SKY130_OSU_SC_15T_MS__AOI22_L%Y N_Y_M1002_d N_Y_M1004_d N_Y_c_251_n
+ N_Y_c_288_n N_Y_c_254_n N_Y_c_255_n N_Y_c_256_n Y N_Y_c_260_n
+ PM_SKY130_OSU_SC_15T_MS__AOI22_L%Y
cc_1 N_GND_M1005_b N_A0_c_77_n 0.0646163f $X=-0.045 $Y=0 $X2=0.295 $Y2=2.37
cc_2 N_GND_M1005_b N_A0_c_78_n 0.0198745f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.43
cc_3 N_GND_c_3_p N_A0_c_78_n 0.00502587f $X=0.26 $Y=0.74 $X2=0.475 $Y2=1.43
cc_4 N_GND_c_4_p N_A0_c_78_n 0.00606474f $X=1.825 $Y=0.152 $X2=0.475 $Y2=1.43
cc_5 N_GND_c_5_p N_A0_c_78_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=1.43
cc_6 N_GND_M1005_b N_A0_c_82_n 0.0322892f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.51
cc_7 N_GND_c_3_p N_A0_c_82_n 0.00587964f $X=0.26 $Y=0.74 $X2=0.475 $Y2=1.51
cc_8 N_GND_M1005_b N_A0_c_84_n 0.0421132f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.505
cc_9 N_GND_M1005_b N_A0_c_85_n 0.00438599f $X=-0.045 $Y=0 $X2=0.385 $Y2=2.505
cc_10 N_GND_M1005_b N_A1_M1002_g 0.0384231f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_11 N_GND_c_4_p N_A1_M1002_g 0.00606474f $X=1.825 $Y=0.152 $X2=0.835 $Y2=0.945
cc_12 N_GND_c_5_p N_A1_M1002_g 0.00468827f $X=1.7 $Y=0.19 $X2=0.835 $Y2=0.945
cc_13 N_GND_M1005_b N_A1_c_115_n 0.0512047f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.31
cc_14 N_GND_M1005_b N_A1_M1003_g 0.0173082f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_15 N_GND_M1005_b N_A1_c_117_n 0.0119461f $X=-0.045 $Y=0 $X2=0.725 $Y2=1.995
cc_16 N_GND_M1005_b A1 0.00204783f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.7
cc_17 N_GND_M1005_b N_B0_M1001_g 0.0194676f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.945
cc_18 N_GND_c_4_p N_B0_M1001_g 0.00606474f $X=1.825 $Y=0.152 $X2=1.335 $Y2=0.945
cc_19 N_GND_c_5_p N_B0_M1001_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.335 $Y2=0.945
cc_20 N_GND_M1005_b N_B0_M1004_g 0.0444247f $X=-0.045 $Y=0 $X2=1.335 $Y2=3.825
cc_21 N_GND_M1005_b N_B0_c_160_n 0.0272094f $X=-0.045 $Y=0 $X2=1.255 $Y2=1.64
cc_22 N_GND_M1005_b N_B0_c_161_n 0.0123234f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.33
cc_23 N_GND_M1005_b N_B0_c_162_n 0.00417976f $X=-0.045 $Y=0 $X2=1.165 $Y2=1.64
cc_24 N_GND_M1005_b B0 0.014652f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.33
cc_25 N_GND_M1005_b N_B1_M1007_g 0.0434394f $X=-0.045 $Y=0 $X2=1.695 $Y2=0.945
cc_26 N_GND_c_4_p N_B1_M1007_g 0.00606474f $X=1.825 $Y=0.152 $X2=1.695 $Y2=0.945
cc_27 N_GND_c_27_p N_B1_M1007_g 0.00502587f $X=1.91 $Y=0.74 $X2=1.695 $Y2=0.945
cc_28 N_GND_c_5_p N_B1_M1007_g 0.00468827f $X=1.7 $Y=0.19 $X2=1.695 $Y2=0.945
cc_29 N_GND_M1005_b N_B1_M1000_g 0.0420537f $X=-0.045 $Y=0 $X2=1.765 $Y2=3.825
cc_30 N_GND_M1005_b N_B1_c_204_n 0.057746f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.945
cc_31 N_GND_c_27_p N_B1_c_204_n 0.00170921f $X=1.91 $Y=0.74 $X2=1.765 $Y2=1.945
cc_32 N_GND_M1005_b N_B1_c_206_n 0.00941038f $X=-0.045 $Y=0 $X2=1.935 $Y2=1.965
cc_33 N_GND_c_27_p N_B1_c_206_n 0.00365739f $X=1.91 $Y=0.74 $X2=1.935 $Y2=1.965
cc_34 N_GND_M1005_b B1 0.0102806f $X=-0.045 $Y=0 $X2=1.935 $Y2=1.965
cc_35 N_GND_c_27_p B1 0.00183474f $X=1.91 $Y=0.74 $X2=1.935 $Y2=1.965
cc_36 N_GND_M1005_b N_Y_c_251_n 0.00156987f $X=-0.045 $Y=0 $X2=1.085 $Y2=0.74
cc_37 N_GND_c_4_p N_Y_c_251_n 0.00738471f $X=1.825 $Y=0.152 $X2=1.085 $Y2=0.74
cc_38 N_GND_c_5_p N_Y_c_251_n 0.00476747f $X=1.7 $Y=0.19 $X2=1.085 $Y2=0.74
cc_39 N_GND_M1005_b N_Y_c_254_n 0.0173806f $X=-0.045 $Y=0 $X2=1.595 $Y2=1.59
cc_40 N_GND_c_27_p N_Y_c_255_n 0.00410021f $X=1.91 $Y=0.74 $X2=1.52 $Y2=1.22
cc_41 N_GND_M1005_b N_Y_c_256_n 0.00670877f $X=-0.045 $Y=0 $X2=1.23 $Y2=1.22
cc_42 N_GND_c_3_p N_Y_c_256_n 0.00341553f $X=0.26 $Y=0.74 $X2=1.23 $Y2=1.22
cc_43 N_GND_c_27_p N_Y_c_256_n 6.58722e-19 $X=1.91 $Y=0.74 $X2=1.23 $Y2=1.22
cc_44 N_GND_M1005_b Y 0.00206172f $X=-0.045 $Y=0 $X2=1.605 $Y2=1.44
cc_45 N_GND_M1005_b N_Y_c_260_n 0.00421975f $X=-0.045 $Y=0 $X2=1.595 $Y2=1.59
cc_46 N_VDD_M1006_b N_A0_M1006_g 0.0262808f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_47 N_VDD_c_47_p N_A0_M1006_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_48 N_VDD_c_48_p N_A0_M1006_g 0.00308284f $X=0.69 $Y=3.98 $X2=0.475 $Y2=3.825
cc_49 N_VDD_c_49_p N_A0_M1006_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.475 $Y2=3.825
cc_50 N_VDD_M1006_b N_A0_c_85_n 0.00618364f $X=-0.045 $Y=2.645 $X2=0.385
+ $Y2=2.505
cc_51 N_VDD_M1006_d A0 0.00594715f $X=0.55 $Y=2.825 $X2=0.385 $Y2=3.07
cc_52 N_VDD_M1006_b N_A1_M1003_g 0.0193371f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_53 N_VDD_c_48_p N_A1_M1003_g 0.00153861f $X=0.69 $Y=3.98 $X2=0.905 $Y2=3.825
cc_54 N_VDD_c_54_p N_A1_M1003_g 0.00496961f $X=1.7 $Y=5.33 $X2=0.905 $Y2=3.825
cc_55 N_VDD_c_49_p N_A1_M1003_g 0.00429146f $X=1.7 $Y=5.36 $X2=0.905 $Y2=3.825
cc_56 N_VDD_M1006_b N_A1_c_117_n 0.00527425f $X=-0.045 $Y=2.645 $X2=0.725
+ $Y2=1.995
cc_57 N_VDD_M1006_b A1 0.0104103f $X=-0.045 $Y=2.645 $X2=0.725 $Y2=2.7
cc_58 N_VDD_M1006_b N_B0_M1004_g 0.0198136f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=3.825
cc_59 N_VDD_c_54_p N_B0_M1004_g 0.00354967f $X=1.7 $Y=5.33 $X2=1.335 $Y2=3.825
cc_60 N_VDD_c_49_p N_B0_M1004_g 0.00429146f $X=1.7 $Y=5.36 $X2=1.335 $Y2=3.825
cc_61 N_VDD_M1006_b N_B1_M1000_g 0.027205f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=3.825
cc_62 N_VDD_c_54_p N_B1_M1000_g 0.00354967f $X=1.7 $Y=5.33 $X2=1.765 $Y2=3.825
cc_63 N_VDD_c_49_p N_B1_M1000_g 0.00429146f $X=1.7 $Y=5.36 $X2=1.765 $Y2=3.825
cc_64 N_VDD_M1006_b N_A_27_565#_c_226_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=4.66
cc_65 N_VDD_c_47_p N_A_27_565#_c_226_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=4.66
cc_66 N_VDD_c_49_p N_A_27_565#_c_226_n 0.00435496f $X=1.7 $Y=5.36 $X2=0.26
+ $Y2=4.66
cc_67 N_VDD_M1006_d N_A_27_565#_c_229_n 0.00734238f $X=0.55 $Y=2.825 $X2=1.035
+ $Y2=3.56
cc_68 N_VDD_c_48_p N_A_27_565#_c_229_n 0.0135055f $X=0.69 $Y=3.98 $X2=1.035
+ $Y2=3.56
cc_69 N_VDD_M1006_b N_A_27_565#_c_231_n 0.00984781f $X=-0.045 $Y=2.645 $X2=1.895
+ $Y2=4.837
cc_70 N_VDD_c_54_p N_A_27_565#_c_231_n 0.0297366f $X=1.7 $Y=5.33 $X2=1.895
+ $Y2=4.837
cc_71 N_VDD_c_49_p N_A_27_565#_c_231_n 0.0226548f $X=1.7 $Y=5.36 $X2=1.895
+ $Y2=4.837
cc_72 N_VDD_M1006_b N_A_27_565#_c_234_n 0.0025777f $X=-0.045 $Y=2.645 $X2=1.205
+ $Y2=4.837
cc_73 N_VDD_c_48_p N_A_27_565#_c_234_n 0.0062002f $X=0.69 $Y=3.98 $X2=1.205
+ $Y2=4.837
cc_74 N_VDD_c_54_p N_A_27_565#_c_234_n 0.00644532f $X=1.7 $Y=5.33 $X2=1.205
+ $Y2=4.837
cc_75 N_VDD_c_49_p N_A_27_565#_c_234_n 0.0046901f $X=1.7 $Y=5.36 $X2=1.205
+ $Y2=4.837
cc_76 N_VDD_M1006_b N_Y_c_254_n 0.00371086f $X=-0.045 $Y=2.645 $X2=1.595
+ $Y2=1.59
cc_77 N_A0_c_77_n N_A1_M1002_g 0.00899556f $X=0.295 $Y=2.37 $X2=0.835 $Y2=0.945
cc_78 N_A0_c_78_n N_A1_M1002_g 0.0701308f $X=0.475 $Y=1.43 $X2=0.835 $Y2=0.945
cc_79 N_A0_c_77_n N_A1_c_115_n 0.0253071f $X=0.295 $Y=2.37 $X2=0.905 $Y2=2.31
cc_80 N_A0_c_77_n N_A1_M1003_g 0.00107789f $X=0.295 $Y=2.37 $X2=0.905 $Y2=3.825
cc_81 N_A0_c_84_n N_A1_M1003_g 0.0676965f $X=0.475 $Y=2.505 $X2=0.905 $Y2=3.825
cc_82 N_A0_c_85_n N_A1_M1003_g 0.00277246f $X=0.385 $Y=2.505 $X2=0.905 $Y2=3.825
cc_83 A0 N_A1_M1003_g 0.00309207f $X=0.385 $Y=3.07 $X2=0.905 $Y2=3.825
cc_84 N_A0_c_77_n N_A1_c_117_n 0.00549523f $X=0.295 $Y=2.37 $X2=0.725 $Y2=1.995
cc_85 N_A0_c_84_n N_A1_c_117_n 0.00281397f $X=0.475 $Y=2.505 $X2=0.725 $Y2=1.995
cc_86 N_A0_c_85_n N_A1_c_117_n 0.0297299f $X=0.385 $Y=2.505 $X2=0.725 $Y2=1.995
cc_87 N_A0_c_84_n A1 0.00417236f $X=0.475 $Y=2.505 $X2=0.725 $Y2=2.7
cc_88 N_A0_c_85_n A1 0.00775911f $X=0.385 $Y=2.505 $X2=0.725 $Y2=2.7
cc_89 A0 A1 0.00560453f $X=0.385 $Y=3.07 $X2=0.725 $Y2=2.7
cc_90 N_A0_c_85_n N_A_27_565#_M1006_s 0.00871729f $X=0.385 $Y=2.505 $X2=0.135
+ $Y2=2.825
cc_91 A0 N_A_27_565#_M1006_s 0.0121636f $X=0.385 $Y=3.07 $X2=0.135 $Y2=2.825
cc_92 N_A0_c_85_n N_A_27_565#_c_240_n 0.00155667f $X=0.385 $Y=2.505 $X2=0.26
+ $Y2=3.645
cc_93 A0 N_A_27_565#_c_240_n 0.00416599f $X=0.385 $Y=3.07 $X2=0.26 $Y2=3.645
cc_94 N_A0_M1006_g N_A_27_565#_c_229_n 0.0136167f $X=0.475 $Y=3.825 $X2=1.035
+ $Y2=3.56
cc_95 N_A0_c_85_n N_A_27_565#_c_229_n 0.00253579f $X=0.385 $Y=2.505 $X2=1.035
+ $Y2=3.56
cc_96 A0 N_A_27_565#_c_229_n 0.00927475f $X=0.385 $Y=3.07 $X2=1.035 $Y2=3.56
cc_97 N_A1_M1002_g N_B0_M1001_g 0.0129165f $X=0.835 $Y=0.945 $X2=1.335 $Y2=0.945
cc_98 N_A1_M1002_g N_B0_M1004_g 0.00961043f $X=0.835 $Y=0.945 $X2=1.335
+ $Y2=3.825
cc_99 N_A1_c_115_n N_B0_M1004_g 0.0638946f $X=0.905 $Y=2.31 $X2=1.335 $Y2=3.825
cc_100 A1 N_B0_M1004_g 0.0011808f $X=0.725 $Y=2.7 $X2=1.335 $Y2=3.825
cc_101 N_A1_M1002_g N_B0_c_160_n 0.0198874f $X=0.835 $Y=0.945 $X2=1.255 $Y2=1.64
cc_102 N_A1_M1002_g N_B0_c_161_n 0.0032219f $X=0.835 $Y=0.945 $X2=1.165 $Y2=2.33
cc_103 N_A1_c_115_n N_B0_c_161_n 0.0017522f $X=0.905 $Y=2.31 $X2=1.165 $Y2=2.33
cc_104 N_A1_c_117_n N_B0_c_161_n 0.0272019f $X=0.725 $Y=1.995 $X2=1.165 $Y2=2.33
cc_105 N_A1_M1002_g N_B0_c_162_n 0.00591675f $X=0.835 $Y=0.945 $X2=1.165
+ $Y2=1.64
cc_106 N_A1_c_115_n B0 0.0041793f $X=0.905 $Y=2.31 $X2=1.165 $Y2=2.33
cc_107 N_A1_M1003_g B0 0.00301191f $X=0.905 $Y=3.825 $X2=1.165 $Y2=2.33
cc_108 N_A1_c_117_n B0 0.0073589f $X=0.725 $Y=1.995 $X2=1.165 $Y2=2.33
cc_109 A1 B0 0.00582284f $X=0.725 $Y=2.7 $X2=1.165 $Y2=2.33
cc_110 N_A1_M1003_g N_A_27_565#_c_229_n 0.0174975f $X=0.905 $Y=3.825 $X2=1.035
+ $Y2=3.56
cc_111 N_A1_M1003_g N_A_27_565#_c_234_n 9.82882e-19 $X=0.905 $Y=3.825 $X2=1.205
+ $Y2=4.837
cc_112 N_A1_M1002_g N_Y_c_251_n 0.00633102f $X=0.835 $Y=0.945 $X2=1.085 $Y2=0.74
cc_113 A1 N_Y_c_254_n 0.00544969f $X=0.725 $Y=2.7 $X2=1.595 $Y2=1.59
cc_114 N_A1_M1002_g N_Y_c_256_n 0.00425578f $X=0.835 $Y=0.945 $X2=1.23 $Y2=1.22
cc_115 N_B0_M1001_g N_B1_M1007_g 0.0451872f $X=1.335 $Y=0.945 $X2=1.695
+ $Y2=0.945
cc_116 N_B0_c_162_n N_B1_M1007_g 4.28971e-19 $X=1.165 $Y=1.64 $X2=1.695
+ $Y2=0.945
cc_117 N_B0_M1004_g N_B1_c_204_n 0.0743876f $X=1.335 $Y=3.825 $X2=1.765
+ $Y2=1.945
cc_118 N_B0_c_160_n N_B1_c_204_n 0.0451872f $X=1.255 $Y=1.64 $X2=1.765 $Y2=1.945
cc_119 N_B0_M1004_g N_A_27_565#_c_231_n 0.0133618f $X=1.335 $Y=3.825 $X2=1.895
+ $Y2=4.837
cc_120 N_B0_M1001_g N_Y_c_251_n 0.00630825f $X=1.335 $Y=0.945 $X2=1.085 $Y2=0.74
cc_121 N_B0_c_160_n N_Y_c_251_n 0.00113527f $X=1.255 $Y=1.64 $X2=1.085 $Y2=0.74
cc_122 N_B0_c_162_n N_Y_c_251_n 0.00420445f $X=1.165 $Y=1.64 $X2=1.085 $Y2=0.74
cc_123 N_B0_c_160_n N_Y_c_254_n 0.0171279f $X=1.255 $Y=1.64 $X2=1.595 $Y2=1.59
cc_124 N_B0_c_161_n N_Y_c_254_n 0.0300971f $X=1.165 $Y=2.33 $X2=1.595 $Y2=1.59
cc_125 N_B0_c_162_n N_Y_c_254_n 0.0201907f $X=1.165 $Y=1.64 $X2=1.595 $Y2=1.59
cc_126 B0 N_Y_c_254_n 0.00659034f $X=1.165 $Y=2.33 $X2=1.595 $Y2=1.59
cc_127 N_B0_M1001_g N_Y_c_255_n 0.0119352f $X=1.335 $Y=0.945 $X2=1.52 $Y2=1.22
cc_128 N_B0_c_162_n N_Y_c_255_n 0.00477495f $X=1.165 $Y=1.64 $X2=1.52 $Y2=1.22
cc_129 N_B0_c_160_n N_Y_c_256_n 0.00131678f $X=1.255 $Y=1.64 $X2=1.23 $Y2=1.22
cc_130 N_B0_c_162_n N_Y_c_256_n 0.00568984f $X=1.165 $Y=1.64 $X2=1.23 $Y2=1.22
cc_131 N_B0_M1001_g Y 0.0019765f $X=1.335 $Y=0.945 $X2=1.605 $Y2=1.44
cc_132 N_B0_c_160_n N_Y_c_260_n 0.00382225f $X=1.255 $Y=1.64 $X2=1.595 $Y2=1.59
cc_133 N_B0_c_162_n N_Y_c_260_n 0.00751098f $X=1.165 $Y=1.64 $X2=1.595 $Y2=1.59
cc_134 N_B1_M1000_g N_A_27_565#_c_231_n 0.0143205f $X=1.765 $Y=3.825 $X2=1.895
+ $Y2=4.837
cc_135 N_B1_M1007_g N_Y_c_254_n 0.0097422f $X=1.695 $Y=0.945 $X2=1.595 $Y2=1.59
cc_136 N_B1_c_204_n N_Y_c_254_n 0.0264693f $X=1.765 $Y=1.945 $X2=1.595 $Y2=1.59
cc_137 N_B1_c_206_n N_Y_c_254_n 0.0209874f $X=1.935 $Y=1.965 $X2=1.595 $Y2=1.59
cc_138 B1 N_Y_c_254_n 0.00769441f $X=1.935 $Y=1.965 $X2=1.595 $Y2=1.59
cc_139 N_B1_M1007_g N_Y_c_255_n 0.00794679f $X=1.695 $Y=0.945 $X2=1.52 $Y2=1.22
cc_140 N_B1_M1007_g Y 0.00642782f $X=1.695 $Y=0.945 $X2=1.605 $Y2=1.44
cc_141 N_B1_M1007_g N_Y_c_260_n 0.0113776f $X=1.695 $Y=0.945 $X2=1.595 $Y2=1.59
cc_142 B1 N_Y_c_260_n 0.00545275f $X=1.935 $Y=1.965 $X2=1.595 $Y2=1.59
cc_143 N_A_27_565#_c_231_n N_Y_M1004_d 0.00215867f $X=1.895 $Y=4.837 $X2=1.41
+ $Y2=2.825
cc_144 N_A_27_565#_c_231_n N_Y_c_288_n 0.00974313f $X=1.895 $Y=4.837 $X2=1.55
+ $Y2=3.64
cc_145 N_Y_c_255_n A_282_115# 0.0104934f $X=1.52 $Y=1.22 $X2=1.41 $Y2=0.575
