magic
tech sky130A
magscale 1 2
timestamp 1612373740
<< nwell >>
rect -9 529 375 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 238 115 268 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 238 565 268 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 166 243
rect 110 131 121 215
rect 155 131 166 215
rect 110 115 166 131
rect 196 115 238 243
rect 268 215 321 243
rect 268 131 279 215
rect 313 131 321 215
rect 268 115 321 131
<< pdiff >>
rect 27 949 80 965
rect 27 605 35 949
rect 69 605 80 949
rect 27 565 80 605
rect 110 949 166 965
rect 110 673 121 949
rect 155 673 166 949
rect 110 565 166 673
rect 196 565 238 965
rect 268 949 321 965
rect 268 605 279 949
rect 313 605 321 949
rect 268 565 321 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 279 131 313 215
<< pdiffc >>
rect 35 605 69 949
rect 121 673 155 949
rect 279 605 313 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 238 965 268 991
rect 80 550 110 565
rect 39 520 110 550
rect 39 308 69 520
rect 166 477 196 565
rect 133 461 196 477
rect 133 427 143 461
rect 177 427 196 461
rect 133 411 196 427
rect 238 399 268 565
rect 238 383 292 399
rect 111 335 165 351
rect 111 308 121 335
rect 39 301 121 308
rect 155 308 165 335
rect 238 349 248 383
rect 282 349 292 383
rect 238 333 292 349
rect 155 301 196 308
rect 39 278 196 301
rect 80 243 110 278
rect 166 243 196 278
rect 238 243 268 333
rect 80 89 110 115
rect 166 89 196 115
rect 238 89 268 115
<< polycont >>
rect 143 427 177 461
rect 121 301 155 335
rect 248 349 282 383
<< locali >>
rect 0 1089 374 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 374 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 657 155 673
rect 279 949 313 965
rect 35 461 69 605
rect 143 461 177 477
rect 35 427 143 461
rect 35 215 69 427
rect 143 411 177 427
rect 211 383 245 597
rect 279 483 313 605
rect 211 349 248 383
rect 282 349 298 383
rect 103 301 121 335
rect 155 301 171 335
rect 35 115 69 131
rect 121 215 155 231
rect 121 61 155 131
rect 279 215 313 227
rect 279 115 313 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 211 597 245 631
rect 279 449 313 483
rect 121 301 155 335
rect 279 227 313 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 374 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 374 1089
rect 0 1049 374 1055
rect 199 631 257 637
rect 177 597 211 631
rect 245 597 257 631
rect 199 591 257 597
rect 109 557 167 563
rect 109 523 189 557
rect 109 517 167 523
rect 121 341 155 517
rect 267 483 325 489
rect 267 449 279 483
rect 313 449 325 483
rect 267 443 325 449
rect 109 335 167 341
rect 109 301 121 335
rect 155 301 167 335
rect 109 295 167 301
rect 279 267 313 443
rect 267 261 325 267
rect 267 227 279 261
rect 313 227 325 261
rect 267 221 325 227
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 305 312 305 312 1 Y
port 1 n
rlabel viali 228 614 228 614 1 A
port 2 n
rlabel metal1 138 540 138 540 1 OE
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
