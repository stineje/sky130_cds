* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_18T_hs__dffsr_1
** N=32 EP=0 IP=0 FDC=43
M0 4 RN gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=575 $D=19
M1 9 4 gnd gnd nlowvt L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=1360 $Y=575 $D=19
M2 21 SN 9 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1850 $Y=575 $D=19
M3 gnd 6 21 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2210 $Y=575 $D=19
M4 22 D gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3160 $Y=575 $D=19
M5 6 10 22 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3520 $Y=575 $D=19
M6 23 CK 6 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4120 $Y=575 $D=19
M7 gnd 9 23 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4480 $Y=575 $D=19
M8 24 9 gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4910 $Y=575 $D=19
M9 12 CK 24 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5270 $Y=575 $D=19
M10 25 10 12 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5870 $Y=575 $D=19
M11 gnd 11 25 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6230 $Y=575 $D=19
M12 10 CK gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6660 $Y=575 $D=19
M13 26 12 gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7610 $Y=575 $D=19
M14 11 SN 26 gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7970 $Y=575 $D=19
M15 gnd 4 11 gnd nlowvt L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=8460 $Y=575 $D=19
M16 gnd 11 QN gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9420 $Y=575 $D=19
M17 Q QN gnd gnd nlowvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9850 $Y=575 $D=19
M18 4 RN vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=400 $Y=3085 $D=79
M19 14 4 9 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=1350 $Y=3085 $D=79
M20 vdd SN 14 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=1780 $Y=3085 $D=79
M21 14 6 vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=2210 $Y=3085 $D=79
M22 15 D vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=3160 $Y=3085 $D=79
M23 6 CK 15 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=3520 $Y=3085 $D=79
M24 16 10 6 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=4120 $Y=3085 $D=79
M25 vdd 9 16 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=4480 $Y=3085 $D=79
M26 17 9 vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=4910 $Y=3085 $D=79
M27 12 10 17 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=5270 $Y=3085 $D=79
M28 18 CK 12 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=5870 $Y=3085 $D=79
M29 vdd 11 18 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=6230 $Y=3085 $D=79
M30 10 CK vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=6660 $Y=3085 $D=79
M31 vdd 12 19 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=7610 $Y=3085 $D=79
M32 19 SN vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=8040 $Y=3085 $D=79
M33 11 4 19 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=8470 $Y=3085 $D=79
M34 vdd 11 QN vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=9420 $Y=3085 $D=79
M35 Q QN vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=9850 $Y=3085 $D=79
X36 gnd vdd Dpar a=39.9 p=28.6 m=1 $[nwdiode] $X=-50 $Y=2905 $D=185
X37 27 RN Probe probetype=1 $[RN] $X=323 $Y=3328 $D=289
X38 28 D Probe probetype=1 $[D] $X=3293 $Y=2218 $D=289
X39 29 CK Probe probetype=1 $[CK] $X=6878 $Y=2588 $D=289
X40 30 SN Probe probetype=1 $[SN] $X=7933 $Y=2958 $D=289
X41 31 QN Probe probetype=1 $[QN] $X=9283 $Y=2958 $D=289
X42 32 Q Probe probetype=1 $[Q] $X=10138 $Y=3328 $D=289
.ENDS
***************************************
