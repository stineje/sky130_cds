* File: sky130_osu_sc_18T_hs__buf_8.pex.spice
* Created: Fri Nov 12 13:48:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__BUF_8%GND 1 2 3 4 5 57 59 67 69 76 78 85 87 94
+ 96 104 115 117
r119 115 117 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r120 102 104 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.13 $Y=0.305
+ $X2=4.13 $Y2=0.825
r121 97 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.152
+ $X2=3.27 $Y2=0.152
r122 96 102 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.045 $Y=0.152
+ $X2=4.13 $Y2=0.305
r123 92 111 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.152
r124 92 94 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.825
r125 87 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.152
+ $X2=3.27 $Y2=0.152
r126 83 85 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.825
r127 79 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0.152
+ $X2=1.55 $Y2=0.152
r128 74 107 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.152
r129 74 76 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.825
r130 70 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r131 69 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.152
r132 65 106 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r133 65 67 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r134 59 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r135 57 117 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r136 57 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r137 57 83 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.41 $Y2=0.305
r138 57 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.325 $Y2=0.152
r139 57 88 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.495 $Y2=0.152
r140 57 96 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.045 $Y2=0.152
r141 57 97 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.355 $Y2=0.152
r142 57 87 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.185 $Y2=0.152
r143 57 88 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.495 $Y2=0.152
r144 57 78 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r145 57 79 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r146 57 69 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r147 57 70 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r148 57 59 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r149 5 104 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.825
r150 4 94 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.825
r151 3 85 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r152 2 76 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r153 1 67 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_8%VDD 1 2 3 4 5 45 47 54 58 64 68 74 78 84
+ 88 95 105 109
r82 105 109 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.74 $Y2=6.507
r83 95 98 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.13 $Y=3.455
+ $X2=4.13 $Y2=5.835
r84 93 98 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.13 $Y=6.355
+ $X2=4.13 $Y2=5.835
r85 91 109 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=6.47
+ $X2=3.74 $Y2=6.47
r86 89 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=6.507
+ $X2=3.27 $Y2=6.507
r87 89 91 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=3.355 $Y=6.507
+ $X2=3.74 $Y2=6.507
r88 88 93 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.045 $Y=6.507
+ $X2=4.13 $Y2=6.355
r89 88 91 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.045 $Y=6.507
+ $X2=3.74 $Y2=6.507
r90 84 87 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.27 $Y=3.455
+ $X2=3.27 $Y2=5.835
r91 82 103 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.27 $Y=6.355
+ $X2=3.27 $Y2=6.507
r92 82 87 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=6.355
+ $X2=3.27 $Y2=5.835
r93 79 102 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=2.41 $Y2=6.507
r94 79 81 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=3.06 $Y2=6.507
r95 78 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.27 $Y2=6.507
r96 78 81 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.06 $Y2=6.507
r97 74 77 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r98 72 102 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=6.507
r99 72 77 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=5.835
r100 69 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.55 $Y2=6.507
r101 69 71 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.7 $Y2=6.507
r102 68 102 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=2.41 $Y2=6.507
r103 68 71 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=1.7 $Y2=6.507
r104 64 67 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r105 62 100 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=6.507
r106 62 67 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=5.835
r107 59 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r108 59 61 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r109 58 100 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.55 $Y2=6.507
r110 58 61 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.02 $Y2=6.507
r111 54 57 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r112 52 99 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r113 52 57 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r114 49 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r115 47 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r116 47 49 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r117 45 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r118 45 81 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r119 45 102 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r120 45 71 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r121 45 61 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r122 45 49 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r123 5 98 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.99
+ $Y=3.085 $X2=4.13 $Y2=5.835
r124 5 95 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.99
+ $Y=3.085 $X2=4.13 $Y2=3.455
r125 4 87 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=5.835
r126 4 84 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=3.455
r127 3 77 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r128 3 74 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r129 2 67 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r130 2 64 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r131 1 57 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r132 1 54 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_8%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=3.33
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2.48
+ $X2=0.635 $Y2=3.33
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.48 $X2=0.635 $Y2=2.48
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.645
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.315
r45 7 12 994.766 $w=1.5e-07 $l=1.94e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.645
r46 3 11 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.315
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_8%A_27_115# 1 3 11 13 15 17 20 22 24 25 26
+ 27 28 31 33 35 36 38 42 44 46 47 49 53 56 57 59 60 62 66 68 70 71 73 77 79 81
+ 82 84 88 90 92 102 103 104 105 106 107 108 109 110 111 114 118 122 124 127
c232 79 0 1.33323e-19 $X=3.485 $Y=3.01
c233 77 0 1.33323e-19 $X=3.485 $Y=1.075
c234 68 0 1.33323e-19 $X=3.055 $Y=3.01
c235 66 0 1.33323e-19 $X=3.055 $Y=1.075
c236 57 0 1.33323e-19 $X=2.625 $Y=3.01
c237 53 0 1.33323e-19 $X=2.625 $Y=1.075
c238 44 0 1.33323e-19 $X=2.195 $Y=3.01
c239 42 0 1.33323e-19 $X=2.195 $Y=1.075
c240 33 0 1.33323e-19 $X=1.765 $Y=3.01
c241 31 0 1.33323e-19 $X=1.765 $Y=1.075
c242 22 0 1.33323e-19 $X=1.335 $Y=3.01
c243 20 0 1.33323e-19 $X=1.335 $Y=1.075
r244 123 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.935
+ $X2=0.26 $Y2=1.935
r245 122 127 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.965 $Y2=1.935
r246 122 123 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.345 $Y2=1.935
r247 118 120 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r248 116 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=1.935
r249 116 118 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=3.455
r250 112 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=1.935
r251 112 114 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r252 99 127 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.935 $X2=0.965 $Y2=1.935
r253 99 100 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=1.18 $Y2=1.935
r254 97 99 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.935
+ $X2=0.965 $Y2=1.935
r255 95 96 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.935
+ $X2=1.335 $Y2=2.935
r256 93 95 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.935
+ $X2=1.18 $Y2=2.935
r257 90 92 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.915 $Y=3.01
+ $X2=3.915 $Y2=4.585
r258 86 88 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.915 $Y=1.77
+ $X2=3.915 $Y2=1.075
r259 85 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.935
+ $X2=3.485 $Y2=2.935
r260 84 90 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=2.935
+ $X2=3.915 $Y2=3.01
r261 84 85 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.935
+ $X2=3.56 $Y2=2.935
r262 83 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.845
+ $X2=3.485 $Y2=1.845
r263 82 86 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=1.845
+ $X2=3.915 $Y2=1.77
r264 82 83 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.845
+ $X2=3.56 $Y2=1.845
r265 79 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=3.01
+ $X2=3.485 $Y2=2.935
r266 79 81 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.485 $Y=3.01
+ $X2=3.485 $Y2=4.585
r267 75 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.845
r268 75 77 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.075
r269 74 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.935
+ $X2=3.055 $Y2=2.935
r270 73 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.935
+ $X2=3.485 $Y2=2.935
r271 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.935
+ $X2=3.13 $Y2=2.935
r272 72 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.845
+ $X2=3.055 $Y2=1.845
r273 71 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.485 $Y2=1.845
r274 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.13 $Y2=1.845
r275 68 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=3.01
+ $X2=3.055 $Y2=2.935
r276 68 70 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.055 $Y=3.01
+ $X2=3.055 $Y2=4.585
r277 64 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.845
r278 64 66 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.075
r279 63 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.935
+ $X2=2.625 $Y2=2.935
r280 62 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=3.055 $Y2=2.935
r281 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=2.7 $Y2=2.935
r282 61 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.845
+ $X2=2.625 $Y2=1.845
r283 60 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=3.055 $Y2=1.845
r284 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=2.7 $Y2=1.845
r285 57 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=2.935
r286 57 59 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=4.585
r287 56 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.86
+ $X2=2.625 $Y2=2.935
r288 55 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.92
+ $X2=2.625 $Y2=1.845
r289 55 56 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.625 $Y=1.92 $X2=2.625
+ $Y2=2.86
r290 51 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.845
r291 51 53 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.075
r292 50 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.935
+ $X2=2.195 $Y2=2.935
r293 49 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.625 $Y2=2.935
r294 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.27 $Y2=2.935
r295 48 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.195 $Y2=1.845
r296 47 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.625 $Y2=1.845
r297 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.27 $Y2=1.845
r298 44 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=2.935
r299 44 46 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=4.585
r300 40 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.845
r301 40 42 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r302 39 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.935
+ $X2=1.765 $Y2=2.935
r303 38 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=2.195 $Y2=2.935
r304 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=1.84 $Y2=2.935
r305 37 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.765 $Y2=1.845
r306 36 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.845
r307 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r308 33 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=2.935
r309 33 35 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=4.585
r310 29 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.845
r311 29 31 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r312 28 96 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.935
+ $X2=1.335 $Y2=2.935
r313 27 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.765 $Y2=2.935
r314 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.41 $Y2=2.935
r315 25 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.765 $Y2=1.845
r316 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.41 $Y2=1.845
r317 22 96 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=2.935
r318 22 24 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=4.585
r319 18 26 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.41 $Y2=1.845
r320 18 100 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.18 $Y2=1.935
r321 18 20 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r322 17 95 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.86
+ $X2=1.18 $Y2=2.935
r323 16 100 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=1.935
r324 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=2.86
r325 13 93 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=2.935
r326 13 15 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=4.585
r327 9 97 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.935
r328 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.075
r329 3 120 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r330 3 118 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r331 1 114 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68 76
+ 82 89 90 92 94 96 99 100 101 102 103 105 106 107 108 109 110 111
c167 111 0 1.33323e-19 $X=3.7 $Y=2.845
c168 110 0 1.33323e-19 $X=3.7 $Y=1.595
c169 109 0 2.66647e-19 $X=2.985 $Y=2.96
c170 107 0 2.66647e-19 $X=2.985 $Y=1.48
c171 103 0 2.66647e-19 $X=2.125 $Y=2.96
c172 101 0 2.66647e-19 $X=2.125 $Y=1.48
c173 90 0 1.33323e-19 $X=1.12 $Y=2.845
c174 89 0 1.33323e-19 $X=1.12 $Y=1.595
r175 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.7 $Y=2.845
+ $X2=3.7 $Y2=2.96
r176 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.7 $Y=1.595
+ $X2=3.7 $Y2=1.48
r177 110 111 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.7 $Y=1.595
+ $X2=3.7 $Y2=2.845
r178 109 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=2.96
+ $X2=2.84 $Y2=2.96
r179 108 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.555 $Y=2.96
+ $X2=3.7 $Y2=2.96
r180 108 109 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.555 $Y=2.96
+ $X2=2.985 $Y2=2.96
r181 107 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=1.48
+ $X2=2.84 $Y2=1.48
r182 106 125 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.555 $Y=1.48
+ $X2=3.7 $Y2=1.48
r183 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.555 $Y=1.48
+ $X2=2.985 $Y2=1.48
r184 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=2.845
+ $X2=2.84 $Y2=2.96
r185 104 121 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=1.48
r186 104 105 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=2.845
r187 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=2.96
+ $X2=1.98 $Y2=2.96
r188 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.84 $Y2=2.96
r189 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.125 $Y2=2.96
r190 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=1.48
+ $X2=1.98 $Y2=1.48
r191 100 121 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.84 $Y2=1.48
r192 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.125 $Y2=1.48
r193 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.845
+ $X2=1.98 $Y2=2.96
r194 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=1.48
r195 98 99 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=2.845
r196 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.96
+ $X2=1.12 $Y2=2.96
r197 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.98 $Y2=2.96
r198 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.265 $Y2=2.96
r199 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1.48
+ $X2=1.12 $Y2=1.48
r200 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.98 $Y2=1.48
r201 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.265 $Y2=1.48
r202 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.96
r203 90 92 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.27
r204 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=1.48
r205 89 92 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=2.27
r206 85 87 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.7 $Y=3.455
+ $X2=3.7 $Y2=5.835
r207 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=2.96
+ $X2=3.7 $Y2=2.96
r208 82 85 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.7 $Y=2.96
+ $X2=3.7 $Y2=3.455
r209 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=1.48
+ $X2=3.7 $Y2=1.48
r210 76 79 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.7 $Y=0.825
+ $X2=3.7 $Y2=1.48
r211 71 73 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r212 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=2.96
r213 68 71 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=3.455
r214 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=1.48
+ $X2=2.84 $Y2=1.48
r215 62 65 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.84 $Y=0.825
+ $X2=2.84 $Y2=1.48
r216 57 59 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r217 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=2.96
r218 54 57 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=3.455
r219 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=1.48
r220 48 51 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.98 $Y=0.825
+ $X2=1.98 $Y2=1.48
r221 43 45 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r222 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=2.96
r223 40 43 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=3.455
r224 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=1.48
r225 34 37 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.12 $Y=0.825
+ $X2=1.12 $Y2=1.48
r226 12 87 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=5.835
r227 12 85 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=3.455
r228 11 73 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r229 11 71 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r230 10 59 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r231 10 57 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r232 9 45 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r233 9 43 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r234 4 76 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.825
r235 3 62 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r236 2 48 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r237 1 34 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
.ends

