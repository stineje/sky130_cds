* File: sky130_osu_sc_18T_hs__and2_1.spice
* Created: Fri Nov 12 13:46:29 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_hs__and2_1.pex.spice"
.subckt sky130_osu_sc_18T_hs__and2_1  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1005 A_110_115# N_A_M1005_g N_A_27_115#_M1005_s N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1003 N_GND_M1003_d N_B_M1003_g A_110_115# N_GND_M1005_b NLOWVT L=0.15 W=1
+ AD=0.175 AS=0.105 PD=1.35 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75000.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_A_27_115#_M1002_g N_GND_M1003_d N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.265 AS=0.175 PD=2.53 PS=1.35 NRD=0 NRS=8.388 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_27_115#_M1004_d N_A_M1004_g N_VDD_M1004_s N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2 SB=75001
+ A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_B_M1000_g N_A_27_115#_M1004_d N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75000.6
+ A=0.45 P=6.3 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_VDD_M1000_d N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX6_noxref N_GND_M1005_b N_VDD_M1004_b NWDIODE A=7.277 P=11.43
pX7_noxref noxref_8 A A PROBETYPE=1
pX8_noxref noxref_9 B B PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__and2_1.pxi.spice"
*
.ends
*
*
