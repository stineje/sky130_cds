* File: sky130_osu_sc_12T_ms__dff_1.pex.spice
* Created: Fri Nov 12 15:22:21 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%GND 1 2 3 4 5 81 83 91 93 103 105 115 117
+ 124 126 133 152 154
c181 115 0 1.61426e-19 $X=4.215 $Y=0.755
c182 81 0 1.27355e-19 $X=-0.045 $Y=0
r183 152 154 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r184 131 133 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.545 $Y=0.305
+ $X2=6.545 $Y2=0.74
r185 122 124 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.165 $Y=0.305
+ $X2=5.165 $Y2=0.755
r186 118 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.152
+ $X2=4.215 $Y2=0.152
r187 113 141 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.152
r188 113 115 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.755
r189 105 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.152
+ $X2=4.215 $Y2=0.152
r190 101 103 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.465 $Y=0.305
+ $X2=2.465 $Y2=0.74
r191 94 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.152
+ $X2=0.715 $Y2=0.152
r192 89 137 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.152
r193 89 91 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.755
r194 83 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.152
+ $X2=0.715 $Y2=0.152
r195 81 154 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r196 81 152 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r197 81 131 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.545 $Y2=0.305
r198 81 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.46 $Y2=0.152
r199 81 122 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.165 $Y2=0.305
r200 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.08 $Y2=0.152
r201 81 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.25 $Y2=0.152
r202 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.465 $Y2=0.305
r203 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.38 $Y2=0.152
r204 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.55 $Y2=0.152
r205 81 126 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.46 $Y2=0.152
r206 81 127 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.25 $Y2=0.152
r207 81 117 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=5.08 $Y2=0.152
r208 81 118 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.3 $Y2=0.152
r209 81 105 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.13 $Y2=0.152
r210 81 106 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.55 $Y2=0.152
r211 81 93 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.38 $Y2=0.152
r212 81 94 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.8 $Y2=0.152
r213 81 83 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.63 $Y2=0.152
r214 5 133 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.405
+ $Y=0.575 $X2=6.545 $Y2=0.74
r215 4 124 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.575 $X2=5.165 $Y2=0.755
r216 3 115 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.575 $X2=4.215 $Y2=0.755
r217 2 103 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.74
r218 1 91 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.575 $X2=0.715 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%VDD 1 2 3 4 5 61 63 70 72 80 82 90 92 98
+ 100 106 117 120 124
c101 70 0 5.41559e-20 $X=0.715 $Y=3.295
c102 1 0 1.59851e-19 $X=0.575 $Y=2.605
r103 120 124 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=6.46 $Y2=4.287
r104 117 124 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=4.25
+ $X2=6.46 $Y2=4.25
r105 104 117 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=4.135
+ $X2=6.545 $Y2=4.287
r106 104 106 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.545 $Y=4.135
+ $X2=6.545 $Y2=3.615
r107 101 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.25 $Y=4.287
+ $X2=5.165 $Y2=4.287
r108 101 103 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.25 $Y=4.287
+ $X2=5.78 $Y2=4.287
r109 100 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=4.287
+ $X2=6.545 $Y2=4.287
r110 100 103 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.46 $Y=4.287
+ $X2=5.78 $Y2=4.287
r111 96 115 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.165 $Y=4.135
+ $X2=5.165 $Y2=4.287
r112 96 98 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.165 $Y=4.135
+ $X2=5.165 $Y2=3.295
r113 93 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=4.287
+ $X2=4.215 $Y2=4.287
r114 93 95 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.3 $Y=4.287
+ $X2=4.42 $Y2=4.287
r115 92 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=4.287
+ $X2=5.165 $Y2=4.287
r116 92 95 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.08 $Y=4.287
+ $X2=4.42 $Y2=4.287
r117 88 113 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.215 $Y=4.135
+ $X2=4.215 $Y2=4.287
r118 88 90 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.215 $Y=4.135
+ $X2=4.215 $Y2=3.21
r119 85 87 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=4.287
+ $X2=3.74 $Y2=4.287
r120 83 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=4.287
+ $X2=2.465 $Y2=4.287
r121 83 85 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=2.55 $Y=4.287
+ $X2=3.06 $Y2=4.287
r122 82 113 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=4.287
+ $X2=4.215 $Y2=4.287
r123 82 87 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=4.13 $Y=4.287
+ $X2=3.74 $Y2=4.287
r124 78 112 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.465 $Y=4.135
+ $X2=2.465 $Y2=4.287
r125 78 80 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.465 $Y=4.135
+ $X2=2.465 $Y2=3.295
r126 75 77 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r127 73 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=4.287
+ $X2=0.715 $Y2=4.287
r128 73 75 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=0.8 $Y=4.287
+ $X2=1.02 $Y2=4.287
r129 72 112 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=4.287
+ $X2=2.465 $Y2=4.287
r130 72 77 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=4.287
+ $X2=1.7 $Y2=4.287
r131 68 110 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=4.287
r132 68 70 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=3.295
r133 65 120 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r134 63 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=4.287
+ $X2=0.715 $Y2=4.287
r135 63 65 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.63 $Y=4.287
+ $X2=0.34 $Y2=4.287
r136 61 117 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=4.135 $X2=6.46 $Y2=4.22
r137 61 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=4.135 $X2=5.78 $Y2=4.22
r138 61 115 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=4.135 $X2=5.1 $Y2=4.22
r139 61 95 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=4.135 $X2=4.42 $Y2=4.22
r140 61 87 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=4.135 $X2=3.74 $Y2=4.22
r141 61 85 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=4.135 $X2=3.06 $Y2=4.22
r142 61 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r143 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r144 61 75 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r145 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r146 5 106 600 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=2.605 $X2=6.545 $Y2=3.615
r147 4 98 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=2.605 $X2=5.165 $Y2=3.295
r148 3 90 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=4.075
+ $Y=2.605 $X2=4.215 $Y2=3.21
r149 2 80 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=2.605 $X2=2.465 $Y2=3.295
r150 1 70 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.605 $X2=0.715 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%A_75_248# 1 3 13 17 20 22 23 28 29 30 31
+ 32 34 37 42 43 45
c87 29 0 1.29912e-19 $X=1.405 $Y=1.285
c88 28 0 1.59851e-19 $X=0.625 $Y=2.62
c89 22 0 5.41559e-20 $X=0.51 $Y=2.285
r90 45 47 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=1.49 $Y=0.755 $X2=1.59
+ $Y2=0.755
r91 42 44 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.285
+ $X2=0.567 $Y2=2.45
r92 42 43 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.285
+ $X2=0.567 $Y2=2.12
r93 37 39 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=1.59 $Y=2.955
+ $X2=1.59 $Y2=3.635
r94 35 37 2.03372 $w=3.38e-07 $l=6e-08 $layer=LI1_cond $X=1.59 $Y=2.895 $X2=1.59
+ $Y2=2.955
r95 33 45 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.49 $Y=0.935
+ $X2=1.49 $Y2=0.755
r96 33 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.49 $Y=0.935
+ $X2=1.49 $Y2=1.2
r97 31 35 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=1.42 $Y=2.705
+ $X2=1.59 $Y2=2.895
r98 31 32 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.42 $Y=2.705
+ $X2=0.71 $Y2=2.705
r99 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.285
+ $X2=1.49 $Y2=1.2
r100 29 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.405 $Y=1.285
+ $X2=0.71 $Y2=1.285
r101 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=2.62
+ $X2=0.71 $Y2=2.705
r102 28 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.625 $Y=2.62
+ $X2=0.625 $Y2=2.45
r103 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.37
+ $X2=0.71 $Y2=1.285
r104 25 43 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.625 $Y=1.37
+ $X2=0.625 $Y2=2.12
r105 22 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=2.285 $X2=0.51 $Y2=2.285
r106 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.285
+ $X2=0.51 $Y2=2.45
r107 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.285
+ $X2=0.51 $Y2=2.12
r108 20 23 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.45 $Y=1.39
+ $X2=0.45 $Y2=2.12
r109 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.475 $Y=1.24
+ $X2=0.475 $Y2=1.39
r110 17 24 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.5 $Y=3.235
+ $X2=0.5 $Y2=2.45
r111 13 19 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.5 $Y=0.835
+ $X2=0.5 $Y2=1.24
r112 3 39 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.605 $X2=1.59 $Y2=3.635
r113 3 37 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.605 $X2=1.59 $Y2=2.955
r114 1 47 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.575 $X2=1.59 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%D 3 7 10 14 19
c43 19 0 1.41836e-19 $X=0.99 $Y=1.74
c44 10 0 1.12321e-19 $X=0.99 $Y=1.74
r45 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=1.74
+ $X2=0.99 $Y2=1.74
r46 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.74 $X2=0.99 $Y2=1.74
r47 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.74
+ $X2=0.99 $Y2=1.905
r48 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.74
+ $X2=0.99 $Y2=1.575
r49 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.93 $Y=3.235
+ $X2=0.93 $Y2=1.905
r50 3 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.93 $Y=0.835
+ $X2=0.93 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c230 74 0 9.35091e-20 $X=3.435 $Y=2.11
c231 57 0 1.35605e-19 $X=4.575 $Y=2.11
c232 55 0 6.79641e-20 $X=3.185 $Y=2.11
c233 54 0 1.49078e-19 $X=3.495 $Y=2.11
c234 48 0 1.98654e-19 $X=1.83 $Y=1.37
c235 44 0 1.86602e-19 $X=1.745 $Y=2.11
c236 37 0 4.60524e-20 $X=3.58 $Y=2.285
c237 33 0 1.61406e-19 $X=3.1 $Y=1.37
c238 30 0 1.29912e-19 $X=1.83 $Y=1.205
c239 25 0 1.41836e-19 $X=1.35 $Y=2.285
r240 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.725 $Y=2.11
+ $X2=3.58 $Y2=2.11
r241 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.43 $Y=2.11
+ $X2=4.575 $Y2=2.11
r242 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=4.43 $Y=2.11
+ $X2=3.725 $Y2=2.11
r243 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.495 $Y=2.11
+ $X2=1.35 $Y2=2.11
r244 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.435 $Y=2.11
+ $X2=3.58 $Y2=2.11
r245 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=3.435 $Y=2.11
+ $X2=1.495 $Y2=2.11
r246 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.11
+ $X2=3.58 $Y2=2.11
r247 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.58 $Y=2.11
+ $X2=3.58 $Y2=2.285
r248 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.35 $Y=2.11
+ $X2=1.35 $Y2=2.11
r249 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.35 $Y=2.11
+ $X2=1.35 $Y2=2.285
r250 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.575 $Y=2.11
+ $X2=4.575 $Y2=2.11
r251 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.11
+ $X2=4.575 $Y2=2.285
r252 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.11
+ $X2=3.58 $Y2=2.11
r253 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.495 $Y=2.11
+ $X2=3.185 $Y2=2.11
r254 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.025
+ $X2=3.185 $Y2=2.11
r255 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.1 $Y=2.025
+ $X2=3.1 $Y2=1.37
r256 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.83 $Y=2.025
+ $X2=1.83 $Y2=1.37
r257 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.11
+ $X2=1.35 $Y2=2.11
r258 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=2.11
+ $X2=1.83 $Y2=2.025
r259 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.745 $Y=2.11
+ $X2=1.435 $Y2=2.11
r260 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=2.285 $X2=4.575 $Y2=2.285
r261 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=4.457 $Y=1.205
+ $X2=4.457 $Y2=1.355
r262 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=2.285 $X2=3.58 $Y2=2.285
r263 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=2.285
+ $X2=3.58 $Y2=2.45
r264 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.37 $X2=3.1 $Y2=1.37
r265 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.37
+ $X2=3.1 $Y2=1.205
r266 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.37 $X2=1.83 $Y2=1.37
r267 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.37
+ $X2=1.83 $Y2=1.205
r268 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=2.285 $X2=1.35 $Y2=2.285
r269 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=2.285
+ $X2=1.35 $Y2=2.45
r270 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=4.485 $Y=2.12
+ $X2=4.532 $Y2=2.285
r271 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.485 $Y=2.12
+ $X2=4.485 $Y2=1.355
r272 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=4.43 $Y=2.45
+ $X2=4.532 $Y2=2.285
r273 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=4.43 $Y=2.45
+ $X2=4.43 $Y2=3.235
r274 17 40 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.43 $Y=0.835
+ $X2=4.43 $Y2=1.205
r275 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.64 $Y=3.235
+ $X2=3.64 $Y2=2.45
r276 10 34 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.04 $Y=0.835
+ $X2=3.04 $Y2=1.205
r277 7 30 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.89 $Y=0.835
+ $X2=1.89 $Y2=1.205
r278 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.29 $Y=3.235
+ $X2=1.29 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%A_32_115# 1 3 11 15 17 18 21 22 27 31 34
+ 37 41 47 52 56 61 62 63 68
c114 61 0 1.61406e-19 $X=2.42 $Y=1.37
c115 47 0 1.5821e-19 $X=2.42 $Y=2.285
c116 31 0 6.36774e-20 $X=2.68 $Y=3.235
c117 22 0 1.86602e-19 $X=2.325 $Y=2.285
c118 21 0 6.79641e-20 $X=2.605 $Y=2.285
c119 15 0 6.36774e-20 $X=2.25 $Y=3.235
r120 63 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.43 $Y=1.37
+ $X2=0.285 $Y2=1.37
r121 62 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.185 $Y=1.37
+ $X2=2.33 $Y2=1.37
r122 62 63 1.68986 $w=1.7e-07 $l=1.755e-06 $layer=MET1_cond $X=2.185 $Y=1.37
+ $X2=0.43 $Y2=1.37
r123 59 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.33 $Y=1.37
+ $X2=2.33 $Y2=1.37
r124 59 61 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=2.33 $Y=1.33 $X2=2.42
+ $Y2=1.33
r125 54 56 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=2.78
+ $X2=0.285 $Y2=2.78
r126 52 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.285 $Y=1.37
+ $X2=0.285 $Y2=1.37
r127 49 52 4.81931 $w=2.73e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=1.317
+ $X2=0.285 $Y2=1.317
r128 45 61 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.42 $Y=1.455
+ $X2=2.42 $Y2=1.33
r129 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.42 $Y=1.455
+ $X2=2.42 $Y2=2.285
r130 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.285 $Y=2.955
+ $X2=0.285 $Y2=3.635
r131 39 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.865
+ $X2=0.285 $Y2=2.78
r132 39 41 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.285 $Y=2.865
+ $X2=0.285 $Y2=2.955
r133 35 52 3.55113 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.285 $Y=1.18
+ $X2=0.285 $Y2=1.317
r134 35 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.285 $Y=1.18
+ $X2=0.285 $Y2=0.755
r135 34 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=2.695
+ $X2=0.17 $Y2=2.78
r136 33 49 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=1.317
r137 33 34 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=2.695
r138 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.68 $Y=2.42
+ $X2=2.68 $Y2=3.235
r139 25 27 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.68 $Y=1.235
+ $X2=2.68 $Y2=0.835
r140 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=2.285 $X2=2.42 $Y2=2.285
r141 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=2.285
+ $X2=2.42 $Y2=2.285
r142 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=2.285
+ $X2=2.68 $Y2=2.42
r143 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=2.285
+ $X2=2.42 $Y2=2.285
r144 20 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.37 $X2=2.42 $Y2=1.37
r145 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=1.37
+ $X2=2.42 $Y2=1.37
r146 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=1.37
+ $X2=2.68 $Y2=1.235
r147 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=1.37
+ $X2=2.42 $Y2=1.37
r148 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=2.42
+ $X2=2.325 $Y2=2.285
r149 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.25 $Y=2.42
+ $X2=2.25 $Y2=3.235
r150 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=1.235
+ $X2=2.325 $Y2=1.37
r151 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.25 $Y=1.235 $X2=2.25
+ $Y2=0.835
r152 3 43 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.605 $X2=0.285 $Y2=3.635
r153 3 41 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.605 $X2=0.285 $Y2=2.955
r154 1 37 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%A_243_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 50 54 59 63 67 70 74 75
c191 75 0 1.35605e-19 $X=4.5 $Y=1.74
c192 74 0 3.47982e-21 $X=4.645 $Y=1.74
c193 70 0 4.60524e-20 $X=3.725 $Y=1.725
c194 44 0 9.35091e-20 $X=3.58 $Y=1.74
c195 34 0 1.98654e-19 $X=1.41 $Y=1.28
c196 18 0 1.12321e-19 $X=1.89 $Y=3.235
r197 74 75 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.645 $Y=1.74
+ $X2=4.5 $Y2=1.74
r198 70 72 0.0981889 $w=2.26e-07 $l=1.52315e-07 $layer=MET1_cond $X=3.725
+ $Y=1.725 $X2=3.58 $Y2=1.74
r199 70 75 0.959157 $w=1.4e-07 $l=7.75e-07 $layer=MET1_cond $X=3.725 $Y=1.725
+ $X2=4.5 $Y2=1.725
r200 65 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=2.705
+ $X2=4.915 $Y2=2.705
r201 62 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.645 $Y=1.74
+ $X2=4.645 $Y2=1.74
r202 62 63 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=1.725
+ $X2=4.915 $Y2=1.725
r203 59 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.62
+ $X2=4.915 $Y2=2.705
r204 58 63 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.915 $Y=1.825
+ $X2=4.915 $Y2=1.725
r205 58 59 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.915 $Y=1.825
+ $X2=4.915 $Y2=2.62
r206 54 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.645 $Y=2.955
+ $X2=4.645 $Y2=3.635
r207 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=2.79
+ $X2=4.645 $Y2=2.705
r208 52 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=2.79
+ $X2=4.645 $Y2=2.955
r209 48 62 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.645 $Y=1.625
+ $X2=4.645 $Y2=1.725
r210 48 50 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.645 $Y=1.625
+ $X2=4.645 $Y2=0.755
r211 44 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=1.74
+ $X2=3.58 $Y2=1.74
r212 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.74 $X2=3.58 $Y2=1.74
r213 39 41 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=3.58 $Y=1.74
+ $X2=3.58 $Y2=1.825
r214 39 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.74
+ $X2=3.58 $Y2=1.575
r215 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.29 $Y=1.28
+ $X2=1.41 $Y2=1.28
r216 30 40 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.64 $Y=0.835
+ $X2=3.64 $Y2=1.575
r217 27 37 19.8589 $w=1.55e-07 $l=7.5e-08 $layer=POLY_cond $X=3.115 $Y=1.825
+ $X2=3.04 $Y2=1.825
r218 26 41 15.0071 $w=1.6e-07 $l=1.35e-07 $layer=POLY_cond $X=3.445 $Y=1.825
+ $X2=3.58 $Y2=1.825
r219 26 27 152.942 $w=1.6e-07 $l=3.3e-07 $layer=POLY_cond $X=3.445 $Y=1.825
+ $X2=3.115 $Y2=1.825
r220 22 37 5.77175 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=3.04 $Y=1.905
+ $X2=3.04 $Y2=1.825
r221 22 24 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.04 $Y=1.905
+ $X2=3.04 $Y2=3.235
r222 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=1.82
+ $X2=1.89 $Y2=1.82
r223 20 37 19.8589 $w=1.55e-07 $l=7.74597e-08 $layer=POLY_cond $X=2.965 $Y=1.82
+ $X2=3.04 $Y2=1.825
r224 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.965 $Y=1.82
+ $X2=1.965 $Y2=1.82
r225 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=1.895
+ $X2=1.89 $Y2=1.82
r226 16 18 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=1.89 $Y=1.895
+ $X2=1.89 $Y2=3.235
r227 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=1.82
+ $X2=1.89 $Y2=1.82
r228 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.815 $Y=1.82
+ $X2=1.485 $Y2=1.82
r229 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.745
+ $X2=1.485 $Y2=1.82
r230 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.355
+ $X2=1.41 $Y2=1.28
r231 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.41 $Y=1.355
+ $X2=1.41 $Y2=1.745
r232 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.205
+ $X2=1.29 $Y2=1.28
r233 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.29 $Y=1.205
+ $X2=1.29 $Y2=0.835
r234 3 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.605 $X2=4.645 $Y2=3.635
r235 3 54 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.605 $X2=4.645 $Y2=2.955
r236 1 50 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.575 $X2=4.645 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%A_785_89# 1 3 11 15 17 21 25 27 30 31 34
+ 36 40 44 50 55 56 57 59 60 61 66
c164 66 0 7.28655e-20 $X=6.215 $Y=1.74
c165 60 0 1.62658e-19 $X=6.08 $Y=1.74
c166 34 0 1.61426e-19 $X=4.062 $Y=1.812
c167 31 0 1.34149e-19 $X=6.305 $Y=2.49
c168 11 0 1.35097e-19 $X=4 $Y=0.835
r169 60 66 0.0969593 $w=2.3e-07 $l=1.35e-07 $layer=MET1_cond $X=6.08 $Y=1.74
+ $X2=6.215 $Y2=1.74
r170 60 61 0.962882 $w=1.7e-07 $l=1e-06 $layer=MET1_cond $X=6.08 $Y=1.74
+ $X2=5.08 $Y2=1.74
r171 58 61 0.0704148 $w=1.7e-07 $l=1.15888e-07 $layer=MET1_cond $X=5.007
+ $Y=1.825 $X2=5.08 $Y2=1.74
r172 58 59 0.664026 $w=1.45e-07 $l=5.7e-07 $layer=MET1_cond $X=5.007 $Y=1.825
+ $X2=5.007 $Y2=2.395
r173 57 63 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.205 $Y=2.48
+ $X2=4.06 $Y2=2.48
r174 56 59 0.0704148 $w=1.7e-07 $l=1.15521e-07 $layer=MET1_cond $X=4.935 $Y=2.48
+ $X2=5.007 $Y2=2.395
r175 56 57 0.702904 $w=1.7e-07 $l=7.3e-07 $layer=MET1_cond $X=4.935 $Y=2.48
+ $X2=4.205 $Y2=2.48
r176 50 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=1.74
+ $X2=6.215 $Y2=1.74
r177 48 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=1.74
+ $X2=5.595 $Y2=1.74
r178 48 50 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.68 $Y=1.74
+ $X2=6.215 $Y2=1.74
r179 44 46 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.595 $Y=2.955
+ $X2=5.595 $Y2=3.635
r180 42 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.825
+ $X2=5.595 $Y2=1.74
r181 42 44 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=5.595 $Y=1.825
+ $X2=5.595 $Y2=2.955
r182 38 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.655
+ $X2=5.595 $Y2=1.74
r183 38 40 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.595 $Y=1.655
+ $X2=5.595 $Y2=0.755
r184 36 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.06 $Y=2.48
+ $X2=4.06 $Y2=2.48
r185 34 54 5.01943 $w=1.75e-07 $l=7.2e-08 $layer=LI1_cond $X=4.062 $Y=1.812
+ $X2=4.062 $Y2=1.74
r186 34 36 42.3356 $w=1.73e-07 $l=6.68e-07 $layer=LI1_cond $X=4.062 $Y=1.812
+ $X2=4.062 $Y2=2.48
r187 33 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.74 $X2=6.215 $Y2=1.74
r188 30 31 43.105 $w=2e-07 $l=1.3e-07 $layer=POLY_cond $X=6.305 $Y=2.36
+ $X2=6.305 $Y2=2.49
r189 27 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.74 $X2=4.06 $Y2=1.74
r190 27 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.74
+ $X2=4.06 $Y2=1.905
r191 27 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.74
+ $X2=4.06 $Y2=1.575
r192 25 31 239.393 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=6.33 $Y=3.235
+ $X2=6.33 $Y2=2.49
r193 19 33 105.348 $w=2.27e-07 $l=5.12113e-07 $layer=POLY_cond $X=6.33 $Y=1.27
+ $X2=6.242 $Y2=1.74
r194 19 21 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.33 $Y=1.27
+ $X2=6.33 $Y2=0.835
r195 17 33 40.5863 $w=2.27e-07 $l=1.83016e-07 $layer=POLY_cond $X=6.28 $Y=1.905
+ $X2=6.242 $Y2=1.74
r196 17 30 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.28 $Y=1.905
+ $X2=6.28 $Y2=2.36
r197 15 29 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=4 $Y=3.235 $X2=4
+ $Y2=1.905
r198 11 28 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4 $Y=0.835 $X2=4
+ $Y2=1.575
r199 3 46 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=2.605 $X2=5.595 $Y2=3.635
r200 3 44 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=2.605 $X2=5.595 $Y2=2.955
r201 1 40 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.575 $X2=5.595 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%A_623_115# 1 3 9 11 14 19 23 25 26 29 33
+ 36 41 44 45 46 47 54
c120 47 0 2.84175e-19 $X=3.585 $Y=1.37
c121 45 0 1.5821e-19 $X=2.905 $Y=1.37
c122 23 0 1.57671e-19 $X=2.76 $Y=1.37
c123 14 0 3.47982e-21 $X=5.38 $Y=3.235
r124 47 52 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=3.585
+ $Y=1.37 $X2=3.44 $Y2=1.34
r125 46 54 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.37
+ $X2=5.175 $Y2=1.37
r126 46 47 1.39137 $w=1.7e-07 $l=1.445e-06 $layer=MET1_cond $X=5.03 $Y=1.37
+ $X2=3.585 $Y2=1.37
r127 45 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.905 $Y=1.37
+ $X2=2.76 $Y2=1.37
r128 44 52 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=3.295
+ $Y=1.37 $X2=3.44 $Y2=1.34
r129 44 45 0.375524 $w=1.7e-07 $l=3.9e-07 $layer=MET1_cond $X=3.295 $Y=1.37
+ $X2=2.905 $Y2=1.37
r130 41 43 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=3.347 $Y=0.755
+ $X2=3.347 $Y2=1.035
r131 36 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.37
+ $X2=5.175 $Y2=1.37
r132 33 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.44 $Y=1.34
+ $X2=3.44 $Y2=1.34
r133 33 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.44 $Y=1.34
+ $X2=3.44 $Y2=1.035
r134 27 29 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=3.34 $Y=2.79
+ $X2=3.34 $Y2=3.295
r135 25 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=2.705
+ $X2=3.34 $Y2=2.79
r136 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=2.705
+ $X2=2.845 $Y2=2.705
r137 23 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.76 $Y=1.37
+ $X2=2.76 $Y2=1.37
r138 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=2.62
+ $X2=2.845 $Y2=2.705
r139 21 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.76 $Y=2.62
+ $X2=2.76 $Y2=1.37
r140 17 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.37 $X2=5.175 $Y2=1.37
r141 17 19 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.175 $Y=1.37
+ $X2=5.38 $Y2=1.37
r142 12 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.535
+ $X2=5.38 $Y2=1.37
r143 12 14 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=5.38 $Y=1.535
+ $X2=5.38 $Y2=3.235
r144 9 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.205
+ $X2=5.38 $Y2=1.37
r145 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.38 $Y=1.205
+ $X2=5.38 $Y2=0.835
r146 3 29 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=3.115
+ $Y=2.605 $X2=3.34 $Y2=3.295
r147 1 41 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.575 $X2=3.34 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%ON 1 3 11 15 18 23 25 27 29 30 31 34 38
+ 41 43
c76 25 0 1.62658e-19 $X=6.115 $Y=2.195
c77 18 0 7.28655e-20 $X=6.7 $Y=2.015
r78 40 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.115 $Y=2.11
+ $X2=6.115 $Y2=2.11
r79 38 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.7 $Y=2.015 $X2=6.7
+ $Y2=1.745
r80 36 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.7 $Y=2.025 $X2=6.7
+ $Y2=2.015
r81 34 41 5.51377 $w=1.73e-07 $l=8.7e-08 $layer=LI1_cond $X=6.702 $Y=1.658
+ $X2=6.702 $Y2=1.745
r82 33 34 10.9642 $w=1.73e-07 $l=1.73e-07 $layer=LI1_cond $X=6.702 $Y=1.485
+ $X2=6.702 $Y2=1.658
r83 32 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=2.11 $X2=6.115
+ $Y2=2.11
r84 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=2.11
+ $X2=6.7 $Y2=2.025
r85 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=2.11
+ $X2=6.2 $Y2=2.11
r86 29 33 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=6.615 $Y=1.4
+ $X2=6.702 $Y2=1.485
r87 29 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=1.4
+ $X2=6.2 $Y2=1.4
r88 25 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=2.195
+ $X2=6.115 $Y2=2.11
r89 25 27 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=6.115 $Y=2.195
+ $X2=6.115 $Y2=3.615
r90 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=1.315
+ $X2=6.2 $Y2=1.4
r91 21 23 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.115 $Y=1.315
+ $X2=6.115 $Y2=0.74
r92 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=2.015 $X2=6.7 $Y2=2.015
r93 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.015
+ $X2=6.7 $Y2=2.18
r94 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.015
+ $X2=6.7 $Y2=1.85
r95 15 20 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=6.76 $Y=3.235
+ $X2=6.76 $Y2=2.18
r96 11 19 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=6.76 $Y=0.835
+ $X2=6.76 $Y2=1.85
r97 3 27 600 $w=1.7e-07 $l=1.07068e-06 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=2.605 $X2=6.115 $Y2=3.615
r98 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.575 $X2=6.115 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__DFF_1%Q 1 3 13 17 20 24 26 30 33
c24 33 0 1.34149e-19 $X=6.97 $Y=2.48
r25 28 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=1.07
+ $X2=7.09 $Y2=1.07
r26 26 27 18.6961 $w=1.73e-07 $l=2.95e-07 $layer=LI1_cond $X=6.972 $Y=2.88
+ $X2=6.972 $Y2=3.175
r27 22 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.97 $Y=2.48
+ $X2=6.97 $Y2=2.48
r28 22 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.97 $Y=2.48
+ $X2=7.09 $Y2=2.48
r29 20 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=2.395
+ $X2=7.09 $Y2=2.48
r30 19 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.155
+ $X2=7.09 $Y2=1.07
r31 19 20 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.09 $Y=1.155
+ $X2=7.09 $Y2=2.395
r32 17 27 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.975 $Y=3.615
+ $X2=6.975 $Y2=3.175
r33 11 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=0.985
+ $X2=6.975 $Y2=1.07
r34 11 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.975 $Y=0.985
+ $X2=6.975 $Y2=0.74
r35 9 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=2.565
+ $X2=6.97 $Y2=2.48
r36 9 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.97 $Y=2.565
+ $X2=6.97 $Y2=2.88
r37 3 17 600 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=6.835
+ $Y=2.605 $X2=6.975 $Y2=3.615
r38 1 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.575 $X2=6.975 $Y2=0.74
.ends

