* File: sky130_osu_sc_18T_ls__aoi21_l.spice
* Created: Thu Oct 29 17:34:19 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ls__aoi21_l.pex.spice"
.subckt sky130_osu_sc_18T_ls__aoi21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1002 A_110_115# N_A0_M1002_g N_GND_M1002_s N_GND_M1002_b NSHORT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.9 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_110_115# N_GND_M1002_b NSHORT L=0.15 W=1
+ AD=0.184195 AS=0.105 PD=1.54023 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667
+ SA=75000.5 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1004 N_GND_M1004_d N_B0_M1004_g N_Y_M1000_d N_GND_M1002_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.136305 PD=2.01 PS=1.13977 NRD=0 NRS=9.72 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VDD_M1001_d N_A0_M1001_g N_A_27_617#_M1001_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1005 N_A_27_617#_M1005_d N_A1_M1005_g N_VDD_M1001_d N_VDD_M1001_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1003 N_Y_M1003_d N_B0_M1003_g N_A_27_617#_M1005_d N_VDD_M1001_b PHIGHVT L=0.15
+ W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=7.277 P=11.43
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__aoi21_l.pxi.spice"
*
.ends
*
*
