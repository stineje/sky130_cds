* File: sky130_osu_sc_15T_ms__dlat_1.spice
* Created: Fri Nov 12 14:43:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__dlat_1.pex.spice"
.subckt sky130_osu_sc_15T_ms__dlat_1  GND VDD D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1001 A_115_115# N_D_M1001_g N_GND_M1001_s N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1014 N_D_M1014_d N_CK_M1014_g A_115_115# N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1665 AS=0.0777 PD=1.19 PS=0.95 NRD=13.776 NRS=8.1 M=1 R=4.93333
+ SA=75000.6 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 A_307_115# N_A_157_393#_M1009_g N_D_M1014_d N_GND_M1001_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1665 PD=0.95 PS=1.19 NRD=8.1 NRS=13.776 M=1 R=4.93333
+ SA=75001.1 SB=75001 A=0.111 P=1.78 MULT=1
MM1003 N_GND_M1003_d N_A_349_89#_M1003_g A_307_115# N_GND_M1001_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.0777 PD=1.02 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_157_393#_M1004_d N_CK_M1004_g N_GND_M1003_d N_GND_M1001_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_349_89#_M1005_d N_D_M1005_g N_GND_M1005_s N_GND_M1001_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_GND_M1006_d N_A_349_89#_M1006_g N_QN_M1006_s N_GND_M1001_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_Q_M1007_d N_QN_M1007_g N_GND_M1006_d N_GND_M1001_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 A_115_565# N_D_M1002_g N_VDD_M1002_s N_VDD_M1002_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75001.9 A=0.3 P=4.3 MULT=1
MM1000 N_D_M1000_d N_A_157_393#_M1000_g A_115_565# N_VDD_M1002_b PSHORT L=0.15
+ W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75000.5 SB=75001.6 A=0.3 P=4.3 MULT=1
MM1015 A_307_565# N_CK_M1015_g N_D_M1000_d N_VDD_M1002_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333 SA=75001.1
+ SB=75001 A=0.3 P=4.3 MULT=1
MM1008 N_VDD_M1008_d N_A_349_89#_M1008_g A_307_565# N_VDD_M1002_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001.5
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1010 N_A_157_393#_M1010_d N_CK_M1010_g N_VDD_M1008_d N_VDD_M1002_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75001.9 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1011 N_A_349_89#_M1011_d N_D_M1011_g N_VDD_M1011_s N_VDD_M1002_b PSHORT L=0.15
+ W=2 AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.2 A=0.3 P=4.3 MULT=1
MM1012 N_VDD_M1012_d N_A_349_89#_M1012_g N_QN_M1012_s N_VDD_M1002_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1013 N_Q_M1013_d N_QN_M1013_g N_VDD_M1012_d N_VDD_M1002_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX16_noxref N_GND_M1001_b N_VDD_M1002_b NWDIODE A=14.406 P=15.89
pX17_noxref noxref_13 D D PROBETYPE=1
pX18_noxref noxref_14 CK CK PROBETYPE=1
pX19_noxref noxref_15 QN QN PROBETYPE=1
pX20_noxref noxref_16 Q Q PROBETYPE=1
c_753 A_115_565# 0 1.57671e-19 $X=0.575 $Y=2.825
*
.include "sky130_osu_sc_15T_ms__dlat_1.pxi.spice"
*
.ends
*
*
