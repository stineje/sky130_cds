* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_18T_ms__addf_l
** N=25 EP=0 IP=0 FDC=35
M0 gnd A 15 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=575 $D=9
M1 15 B gnd gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=575 $D=9
M2 CON CI 15 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=575 $D=9
M3 16 B CON gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=575 $D=9
M4 gnd A 16 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2050 $Y=575 $D=9
M5 17 A gnd gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2480 $Y=575 $D=9
M6 gnd B 17 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2910 $Y=575 $D=9
M7 17 CI gnd gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3340 $Y=575 $D=9
M8 7 CON 17 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3770 $Y=575 $D=9
M9 18 B 7 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4200 $Y=575 $D=9
M10 19 CI 18 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4610 $Y=575 $D=8
M11 gnd A 19 gnd nshort L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5020 $Y=575 $D=9
M12 S 7 gnd gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=5510 $Y=575 $D=9
M13 CO CON gnd gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=6460 $Y=575 $D=9
M14 vdd A 8 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=400 $Y=3085 $D=79
M15 8 B vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=830 $Y=3085 $D=79
M16 CON CI 8 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=1260 $Y=3085 $D=79
M17 9 B CON vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=1690 $Y=3085 $D=79
M18 vdd A 9 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=2050 $Y=3085 $D=79
M19 10 A vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=2480 $Y=3085 $D=79
M20 vdd B 10 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=2910 $Y=3085 $D=79
M21 10 CI vdd vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=3340 $Y=3085 $D=79
M22 7 CON 10 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=3770 $Y=3085 $D=79
M23 11 B 7 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=4200 $Y=3085 $D=79
M24 12 CI 11 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=4610 $Y=3085 $D=78
M25 vdd A 12 vdd pshort L=0.15 W=3 m=1 r=20 a=0.45 p=6.3 mult=1 $X=5020 $Y=3085 $D=79
M26 S 7 vdd vdd pshort L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=5510 $Y=4085 $D=79
M27 CO CON vdd vdd pshort L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=6460 $Y=4085 $D=79
X28 gnd vdd Dpar a=27.436 p=22.04 m=1 $[nwdiode] $X=-45 $Y=2905 $D=185
X29 20 A Probe probetype=1 $[A] $X=483 $Y=1848 $D=289
X30 21 B Probe probetype=1 $[B] $X=643 $Y=2588 $D=289
X31 22 CI Probe probetype=1 $[CI] $X=1323 $Y=2218 $D=289
X32 23 S Probe probetype=1 $[S] $X=5798 $Y=3363 $D=289
X33 24 CON Probe probetype=1 $[CON] $X=6138 $Y=1478 $D=289
X34 25 CO Probe probetype=1 $[CO] $X=6748 $Y=2958 $D=289
.ENDS
***************************************
