* File: sky130_osu_sc_15T_hs__addh_1.pxi.spice
* Created: Fri Nov 12 14:26:25 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%GND N_GND_M1006_d N_GND_M1001_d N_GND_M1006_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_25_p N_GND_c_9_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_15T_HS__ADDH_1%GND
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%VDD N_VDD_M1009_d N_VDD_M1012_d N_VDD_M1003_d
+ N_VDD_M1009_b N_VDD_c_97_p N_VDD_c_98_p N_VDD_c_111_p N_VDD_c_119_p
+ N_VDD_c_101_p N_VDD_c_104_p N_VDD_c_106_p VDD N_VDD_c_99_p
+ PM_SKY130_OSU_SC_15T_HS__ADDH_1%VDD
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%CON N_CON_M1004_d N_CON_M1003_s N_CON_M1000_d
+ N_CON_M1006_g N_CON_M1009_g N_CON_c_157_n N_CON_c_158_n N_CON_c_160_n
+ N_CON_c_161_n N_CON_c_178_n N_CON_c_162_n N_CON_c_163_n N_CON_c_164_n
+ N_CON_c_165_n N_CON_c_183_n N_CON_c_166_n N_CON_c_167_n N_CON_c_169_n
+ N_CON_c_171_n CON PM_SKY130_OSU_SC_15T_HS__ADDH_1%CON
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%B N_B_M1007_g N_B_M1011_g N_B_M1004_g
+ N_B_M1013_g N_B_c_289_n N_B_c_291_n N_B_c_292_n N_B_c_294_n N_B_c_295_n
+ N_B_c_296_n B PM_SKY130_OSU_SC_15T_HS__ADDH_1%B
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%A N_A_M1008_g N_A_M1012_g N_A_M1000_g
+ N_A_M1005_g N_A_c_390_n N_A_c_391_n N_A_c_392_n N_A_c_393_n N_A_c_394_n A
+ N_A_c_396_n PM_SKY130_OSU_SC_15T_HS__ADDH_1%A
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%A_208_565# N_A_208_565#_M1008_d
+ N_A_208_565#_M1011_d N_A_208_565#_c_470_n N_A_208_565#_c_471_n
+ N_A_208_565#_M1002_g N_A_208_565#_c_473_n N_A_208_565#_c_474_n
+ N_A_208_565#_c_475_n N_A_208_565#_M1001_g N_A_208_565#_c_479_n
+ N_A_208_565#_c_481_n N_A_208_565#_M1010_g N_A_208_565#_M1003_g
+ N_A_208_565#_c_485_n N_A_208_565#_c_486_n N_A_208_565#_c_501_n
+ N_A_208_565#_c_504_n N_A_208_565#_c_507_n N_A_208_565#_c_487_n
+ N_A_208_565#_c_491_n N_A_208_565#_c_492_n
+ PM_SKY130_OSU_SC_15T_HS__ADDH_1%A_208_565#
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%S N_S_M1006_s N_S_M1009_s N_S_c_586_n
+ N_S_c_593_n S N_S_c_591_n N_S_c_598_n PM_SKY130_OSU_SC_15T_HS__ADDH_1%S
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%CO N_CO_M1001_s N_CO_M1002_d N_CO_c_617_n
+ N_CO_c_624_n N_CO_c_620_n N_CO_c_621_n N_CO_c_622_n CO
+ PM_SKY130_OSU_SC_15T_HS__ADDH_1%CO
x_PM_SKY130_OSU_SC_15T_HS__ADDH_1%A_570_115# N_A_570_115#_M1010_d
+ N_A_570_115#_M1005_d N_A_570_115#_c_673_n N_A_570_115#_c_668_n
+ N_A_570_115#_c_670_n PM_SKY130_OSU_SC_15T_HS__ADDH_1%A_570_115#
cc_1 N_GND_M1006_b N_CON_M1006_g 0.029545f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_CON_M1006_g 0.00606474f $X=0.665 $Y=0.152 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_CON_M1006_g 0.00882091f $X=0.75 $Y=0.885 $X2=0.475 $Y2=0.895
cc_4 N_GND_c_4_p N_CON_M1006_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.475 $Y2=0.895
cc_5 N_GND_M1006_b N_CON_M1009_g 0.060974f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.825
cc_6 N_GND_M1006_b N_CON_c_157_n 0.0413643f $X=-0.045 $Y=0 $X2=0.35 $Y2=1.59
cc_7 N_GND_M1006_b N_CON_c_158_n 0.00877401f $X=-0.045 $Y=0 $X2=0.635 $Y2=1.59
cc_8 N_GND_c_3_p N_CON_c_158_n 0.00255942f $X=0.75 $Y=0.885 $X2=0.635 $Y2=1.59
cc_9 N_GND_c_9_p N_CON_c_160_n 0.00470352f $X=2.56 $Y=0.74 $X2=2.62 $Y2=1.675
cc_10 N_GND_M1006_b N_CON_c_161_n 0.0155029f $X=-0.045 $Y=0 $X2=2.62 $Y2=2.605
cc_11 N_GND_M1006_b N_CON_c_162_n 0.0100275f $X=-0.045 $Y=0 $X2=3.335 $Y2=1.59
cc_12 N_GND_M1006_b N_CON_c_163_n 0.0112921f $X=-0.045 $Y=0 $X2=3.755 $Y2=2.69
cc_13 N_GND_M1006_b N_CON_c_164_n 0.00433753f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.505
cc_14 N_GND_M1006_b N_CON_c_165_n 0.00195909f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.065
cc_15 N_GND_M1006_b N_CON_c_166_n 2.79926e-19 $X=-0.045 $Y=0 $X2=2.62 $Y2=2.69
cc_16 N_GND_M1006_b N_CON_c_167_n 0.0196394f $X=-0.045 $Y=0 $X2=2.475 $Y2=1.59
cc_17 N_GND_c_3_p N_CON_c_167_n 0.00167316f $X=0.75 $Y=0.885 $X2=2.475 $Y2=1.59
cc_18 N_GND_M1006_b N_CON_c_169_n 0.0133709f $X=-0.045 $Y=0 $X2=0.78 $Y2=1.59
cc_19 N_GND_c_3_p N_CON_c_169_n 0.00391282f $X=0.75 $Y=0.885 $X2=0.78 $Y2=1.59
cc_20 N_GND_M1006_b N_CON_c_171_n 0.00474051f $X=-0.045 $Y=0 $X2=2.62 $Y2=1.59
cc_21 N_GND_c_9_p N_CON_c_171_n 0.00612077f $X=2.56 $Y=0.74 $X2=2.62 $Y2=1.59
cc_22 N_GND_M1006_b CON 0.00668459f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.59
cc_23 N_GND_M1006_b N_B_M1007_g 0.0399402f $X=-0.045 $Y=0 $X2=0.965 $Y2=0.895
cc_24 N_GND_c_3_p N_B_M1007_g 0.00482006f $X=0.75 $Y=0.885 $X2=0.965 $Y2=0.895
cc_25 N_GND_c_25_p N_B_M1007_g 0.00606474f $X=2.475 $Y=0.152 $X2=0.965 $Y2=0.895
cc_26 N_GND_c_4_p N_B_M1007_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.965 $Y2=0.895
cc_27 N_GND_M1006_b N_B_M1011_g 0.0282323f $X=-0.045 $Y=0 $X2=0.965 $Y2=3.825
cc_28 N_GND_M1006_b N_B_M1004_g 0.0334167f $X=-0.045 $Y=0 $X2=3.205 $Y2=0.995
cc_29 N_GND_c_4_p N_B_M1004_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.205 $Y2=0.995
cc_30 N_GND_M1006_b N_B_M1013_g 0.0272084f $X=-0.045 $Y=0 $X2=3.265 $Y2=3.825
cc_31 N_GND_M1006_b N_B_c_289_n 0.0278498f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.96
cc_32 N_GND_c_3_p N_B_c_289_n 0.00118809f $X=0.75 $Y=0.885 $X2=0.905 $Y2=1.96
cc_33 N_GND_M1006_b N_B_c_291_n 0.0299556f $X=-0.045 $Y=0 $X2=3.205 $Y2=1.96
cc_34 N_GND_M1006_b N_B_c_292_n 0.00405307f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.96
cc_35 N_GND_c_3_p N_B_c_292_n 0.00118993f $X=0.75 $Y=0.885 $X2=0.905 $Y2=1.96
cc_36 N_GND_M1006_b N_B_c_294_n 0.00365598f $X=-0.045 $Y=0 $X2=3.205 $Y2=1.96
cc_37 N_GND_M1006_b N_B_c_295_n 0.00204225f $X=-0.045 $Y=0 $X2=1.05 $Y2=1.96
cc_38 N_GND_M1006_b N_B_c_296_n 0.0175295f $X=-0.045 $Y=0 $X2=3.06 $Y2=1.96
cc_39 N_GND_M1006_b B 0.00164195f $X=-0.045 $Y=0 $X2=3.21 $Y2=1.96
cc_40 N_GND_M1006_b N_A_M1008_g 0.0611551f $X=-0.045 $Y=0 $X2=1.325 $Y2=0.895
cc_41 N_GND_c_25_p N_A_M1008_g 0.00606474f $X=2.475 $Y=0.152 $X2=1.325 $Y2=0.895
cc_42 N_GND_c_4_p N_A_M1008_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.325 $Y2=0.895
cc_43 N_GND_M1006_b N_A_M1012_g 0.00835457f $X=-0.045 $Y=0 $X2=1.395 $Y2=3.825
cc_44 N_GND_M1006_b N_A_M1000_g 0.0108664f $X=-0.045 $Y=0 $X2=3.625 $Y2=3.825
cc_45 N_GND_M1006_b N_A_M1005_g 0.0755267f $X=-0.045 $Y=0 $X2=3.635 $Y2=0.995
cc_46 N_GND_c_4_p N_A_M1005_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.635 $Y2=0.995
cc_47 N_GND_M1006_b N_A_c_390_n 0.0253796f $X=-0.045 $Y=0 $X2=1.385 $Y2=2.33
cc_48 N_GND_M1006_b N_A_c_391_n 0.034256f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.33
cc_49 N_GND_M1006_b N_A_c_392_n 9.49347e-19 $X=-0.045 $Y=0 $X2=1.385 $Y2=2.33
cc_50 N_GND_M1006_b N_A_c_393_n 0.00995238f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.33
cc_51 N_GND_M1006_b N_A_c_394_n 0.00430309f $X=-0.045 $Y=0 $X2=1.53 $Y2=2.33
cc_52 N_GND_M1006_b A 0.00380188f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.33
cc_53 N_GND_M1006_b N_A_c_396_n 0.0115252f $X=-0.045 $Y=0 $X2=3.54 $Y2=2.33
cc_54 N_GND_M1006_b N_A_208_565#_c_470_n 0.0382337f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=1.86
cc_55 N_GND_M1006_b N_A_208_565#_c_471_n 0.0270254f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=2.335
cc_56 N_GND_M1006_b N_A_208_565#_M1002_g 0.00928694f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=3.825
cc_57 N_GND_M1006_b N_A_208_565#_c_473_n 0.0168404f $X=-0.045 $Y=0 $X2=2.21
+ $Y2=1.565
cc_58 N_GND_M1006_b N_A_208_565#_c_474_n 0.0616052f $X=-0.045 $Y=0 $X2=2.76
+ $Y2=2.41
cc_59 N_GND_M1006_b N_A_208_565#_c_475_n 0.0189866f $X=-0.045 $Y=0 $X2=2.285
+ $Y2=1.49
cc_60 N_GND_c_25_p N_A_208_565#_c_475_n 0.00606474f $X=2.475 $Y=0.152 $X2=2.285
+ $Y2=1.49
cc_61 N_GND_c_9_p N_A_208_565#_c_475_n 0.00873252f $X=2.56 $Y=0.74 $X2=2.285
+ $Y2=1.49
cc_62 N_GND_c_4_p N_A_208_565#_c_475_n 0.00468827f $X=3.74 $Y=0.19 $X2=2.285
+ $Y2=1.49
cc_63 N_GND_M1006_b N_A_208_565#_c_479_n 0.0273212f $X=-0.045 $Y=0 $X2=2.7
+ $Y2=1.565
cc_64 N_GND_c_9_p N_A_208_565#_c_479_n 0.00319024f $X=2.56 $Y=0.74 $X2=2.7
+ $Y2=1.565
cc_65 N_GND_M1006_b N_A_208_565#_c_481_n 0.0209741f $X=-0.045 $Y=0 $X2=2.775
+ $Y2=1.49
cc_66 N_GND_c_9_p N_A_208_565#_c_481_n 0.00163921f $X=2.56 $Y=0.74 $X2=2.775
+ $Y2=1.49
cc_67 N_GND_c_4_p N_A_208_565#_c_481_n 0.00468827f $X=3.74 $Y=0.19 $X2=2.775
+ $Y2=1.49
cc_68 N_GND_M1006_b N_A_208_565#_M1003_g 0.00900107f $X=-0.045 $Y=0 $X2=2.835
+ $Y2=3.825
cc_69 N_GND_M1006_b N_A_208_565#_c_485_n 0.00492701f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=2.41
cc_70 N_GND_M1006_b N_A_208_565#_c_486_n 0.00608465f $X=-0.045 $Y=0 $X2=2.285
+ $Y2=1.565
cc_71 N_GND_M1006_b N_A_208_565#_c_487_n 0.00877765f $X=-0.045 $Y=0 $X2=1.54
+ $Y2=0.885
cc_72 N_GND_c_3_p N_A_208_565#_c_487_n 8.71428e-19 $X=0.75 $Y=0.885 $X2=1.54
+ $Y2=0.885
cc_73 N_GND_c_25_p N_A_208_565#_c_487_n 0.00741243f $X=2.475 $Y=0.152 $X2=1.54
+ $Y2=0.885
cc_74 N_GND_c_4_p N_A_208_565#_c_487_n 0.00476261f $X=3.74 $Y=0.19 $X2=1.54
+ $Y2=0.885
cc_75 N_GND_M1006_b N_A_208_565#_c_491_n 0.0137594f $X=-0.045 $Y=0 $X2=1.725
+ $Y2=2.665
cc_76 N_GND_M1006_b N_A_208_565#_c_492_n 0.00684174f $X=-0.045 $Y=0 $X2=1.725
+ $Y2=1.695
cc_77 N_GND_M1006_b N_S_c_586_n 0.00480895f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.885
cc_78 N_GND_c_2_p N_S_c_586_n 0.00736239f $X=0.665 $Y=0.152 $X2=0.26 $Y2=0.885
cc_79 N_GND_c_3_p N_S_c_586_n 0.0157284f $X=0.75 $Y=0.885 $X2=0.26 $Y2=0.885
cc_80 N_GND_c_4_p N_S_c_586_n 0.00476261f $X=3.74 $Y=0.19 $X2=0.26 $Y2=0.885
cc_81 N_GND_M1006_b S 0.063433f $X=-0.045 $Y=0 $X2=0.25 $Y2=2.125
cc_82 N_GND_M1006_b N_S_c_591_n 0.0121294f $X=-0.045 $Y=0 $X2=0.26 $Y2=1.215
cc_83 N_GND_c_3_p N_S_c_591_n 0.00348655f $X=0.75 $Y=0.885 $X2=0.26 $Y2=1.215
cc_84 N_GND_M1006_b N_CO_c_617_n 0.00155645f $X=-0.045 $Y=0 $X2=2.07 $Y2=0.74
cc_85 N_GND_c_25_p N_CO_c_617_n 0.00750025f $X=2.475 $Y=0.152 $X2=2.07 $Y2=0.74
cc_86 N_GND_c_4_p N_CO_c_617_n 0.00474053f $X=3.74 $Y=0.19 $X2=2.07 $Y2=0.74
cc_87 N_GND_c_9_p N_CO_c_620_n 0.00482015f $X=2.56 $Y=0.74 $X2=2.175 $Y2=1.25
cc_88 N_GND_M1006_b N_CO_c_621_n 0.00130468f $X=-0.045 $Y=0 $X2=2.175 $Y2=2.7
cc_89 N_GND_M1006_b N_CO_c_622_n 0.0146768f $X=-0.045 $Y=0 $X2=2.137 $Y2=2.615
cc_90 N_GND_M1006_b CO 0.00219851f $X=-0.045 $Y=0 $X2=2.175 $Y2=2.7
cc_91 N_GND_M1006_b N_A_570_115#_c_668_n 0.0652319f $X=-0.045 $Y=0 $X2=3.765
+ $Y2=0.56
cc_92 N_GND_c_4_p N_A_570_115#_c_668_n 0.024842f $X=3.74 $Y=0.19 $X2=3.765
+ $Y2=0.56
cc_93 N_GND_M1006_b N_A_570_115#_c_670_n 0.0145317f $X=-0.045 $Y=0 $X2=3.075
+ $Y2=0.56
cc_94 N_GND_c_9_p N_A_570_115#_c_670_n 0.0062002f $X=2.56 $Y=0.74 $X2=3.075
+ $Y2=0.56
cc_95 N_GND_c_4_p N_A_570_115#_c_670_n 0.00506617f $X=3.74 $Y=0.19 $X2=3.075
+ $Y2=0.56
cc_96 N_VDD_M1009_b N_CON_M1009_g 0.0278142f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_97 N_VDD_c_97_p N_CON_M1009_g 0.00496961f $X=0.665 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_98 N_VDD_c_98_p N_CON_M1009_g 0.0192185f $X=0.75 $Y=3.215 $X2=0.475 $Y2=3.825
cc_99 N_VDD_c_99_p N_CON_M1009_g 0.00429146f $X=3.74 $Y=5.36 $X2=0.475 $Y2=3.825
cc_100 N_VDD_M1009_b N_CON_c_178_n 0.00290115f $X=-0.045 $Y=2.645 $X2=2.62
+ $Y2=3.215
cc_101 N_VDD_c_101_p N_CON_c_178_n 0.00469914f $X=2.965 $Y=5.397 $X2=2.62
+ $Y2=3.215
cc_102 N_VDD_c_99_p N_CON_c_178_n 0.00435496f $X=3.74 $Y=5.36 $X2=2.62 $Y2=3.215
cc_103 N_VDD_M1009_b N_CON_c_163_n 0.0218832f $X=-0.045 $Y=2.645 $X2=3.755
+ $Y2=2.69
cc_104 N_VDD_c_104_p N_CON_c_163_n 0.0121906f $X=3.05 $Y=3.215 $X2=3.755
+ $Y2=2.69
cc_105 N_VDD_M1009_b N_CON_c_183_n 0.00419737f $X=-0.045 $Y=2.645 $X2=3.84
+ $Y2=3.215
cc_106 N_VDD_c_106_p N_CON_c_183_n 0.00452684f $X=3.74 $Y=5.33 $X2=3.84
+ $Y2=3.215
cc_107 N_VDD_c_99_p N_CON_c_183_n 0.00435496f $X=3.74 $Y=5.36 $X2=3.84 $Y2=3.215
cc_108 N_VDD_M1009_b N_CON_c_166_n 0.00108117f $X=-0.045 $Y=2.645 $X2=2.62
+ $Y2=2.69
cc_109 N_VDD_M1009_b N_B_M1011_g 0.0216302f $X=-0.045 $Y=2.645 $X2=0.965
+ $Y2=3.825
cc_110 N_VDD_c_98_p N_B_M1011_g 0.00373151f $X=0.75 $Y=3.215 $X2=0.965 $Y2=3.825
cc_111 N_VDD_c_111_p N_B_M1011_g 0.00496961f $X=1.525 $Y=5.397 $X2=0.965
+ $Y2=3.825
cc_112 N_VDD_c_99_p N_B_M1011_g 0.00429146f $X=3.74 $Y=5.36 $X2=0.965 $Y2=3.825
cc_113 N_VDD_M1009_b N_B_M1013_g 0.0185755f $X=-0.045 $Y=2.645 $X2=3.265
+ $Y2=3.825
cc_114 N_VDD_c_104_p N_B_M1013_g 0.00354579f $X=3.05 $Y=3.215 $X2=3.265
+ $Y2=3.825
cc_115 N_VDD_c_106_p N_B_M1013_g 0.00496961f $X=3.74 $Y=5.33 $X2=3.265 $Y2=3.825
cc_116 N_VDD_c_99_p N_B_M1013_g 0.00429146f $X=3.74 $Y=5.36 $X2=3.265 $Y2=3.825
cc_117 N_VDD_M1009_b N_A_M1012_g 0.0197771f $X=-0.045 $Y=2.645 $X2=1.395
+ $Y2=3.825
cc_118 N_VDD_c_111_p N_A_M1012_g 0.00496961f $X=1.525 $Y=5.397 $X2=1.395
+ $Y2=3.825
cc_119 N_VDD_c_119_p N_A_M1012_g 0.00373151f $X=1.61 $Y=3.555 $X2=1.395
+ $Y2=3.825
cc_120 N_VDD_c_99_p N_A_M1012_g 0.00429146f $X=3.74 $Y=5.36 $X2=1.395 $Y2=3.825
cc_121 N_VDD_M1009_b N_A_M1000_g 0.0243418f $X=-0.045 $Y=2.645 $X2=3.625
+ $Y2=3.825
cc_122 N_VDD_c_106_p N_A_M1000_g 0.00496961f $X=3.74 $Y=5.33 $X2=3.625 $Y2=3.825
cc_123 N_VDD_c_99_p N_A_M1000_g 0.00429146f $X=3.74 $Y=5.36 $X2=3.625 $Y2=3.825
cc_124 N_VDD_M1009_b N_A_208_565#_M1002_g 0.0247637f $X=-0.045 $Y=2.645
+ $X2=1.885 $Y2=3.825
cc_125 N_VDD_c_119_p N_A_208_565#_M1002_g 0.0162477f $X=1.61 $Y=3.555 $X2=1.885
+ $Y2=3.825
cc_126 N_VDD_c_101_p N_A_208_565#_M1002_g 0.00496961f $X=2.965 $Y=5.397
+ $X2=1.885 $Y2=3.825
cc_127 N_VDD_c_99_p N_A_208_565#_M1002_g 0.00429146f $X=3.74 $Y=5.36 $X2=1.885
+ $Y2=3.825
cc_128 N_VDD_M1009_b N_A_208_565#_M1003_g 0.0252169f $X=-0.045 $Y=2.645
+ $X2=2.835 $Y2=3.825
cc_129 N_VDD_c_101_p N_A_208_565#_M1003_g 0.00496961f $X=2.965 $Y=5.397
+ $X2=2.835 $Y2=3.825
cc_130 N_VDD_c_104_p N_A_208_565#_M1003_g 0.00354579f $X=3.05 $Y=3.215 $X2=2.835
+ $Y2=3.825
cc_131 N_VDD_c_99_p N_A_208_565#_M1003_g 0.00429146f $X=3.74 $Y=5.36 $X2=2.835
+ $Y2=3.825
cc_132 N_VDD_M1009_b N_A_208_565#_c_501_n 0.00198641f $X=-0.045 $Y=2.645
+ $X2=1.18 $Y2=3.555
cc_133 N_VDD_c_111_p N_A_208_565#_c_501_n 0.00456907f $X=1.525 $Y=5.397 $X2=1.18
+ $Y2=3.555
cc_134 N_VDD_c_99_p N_A_208_565#_c_501_n 0.00434939f $X=3.74 $Y=5.36 $X2=1.18
+ $Y2=3.555
cc_135 N_VDD_M1012_d N_A_208_565#_c_504_n 0.00566044f $X=1.47 $Y=2.825 $X2=1.64
+ $Y2=2.75
cc_136 N_VDD_M1009_b N_A_208_565#_c_504_n 0.00273697f $X=-0.045 $Y=2.645
+ $X2=1.64 $Y2=2.75
cc_137 N_VDD_c_119_p N_A_208_565#_c_504_n 0.00659105f $X=1.61 $Y=3.555 $X2=1.64
+ $Y2=2.75
cc_138 N_VDD_M1009_b N_A_208_565#_c_507_n 0.00518782f $X=-0.045 $Y=2.645
+ $X2=1.265 $Y2=2.75
cc_139 N_VDD_M1009_b N_A_208_565#_c_491_n 3.89739e-19 $X=-0.045 $Y=2.645
+ $X2=1.725 $Y2=2.665
cc_140 N_VDD_M1009_b N_S_c_593_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.07
cc_141 N_VDD_c_97_p N_S_c_593_n 0.00452684f $X=0.665 $Y=5.397 $X2=0.26 $Y2=3.07
cc_142 N_VDD_c_98_p N_S_c_593_n 0.0426358f $X=0.75 $Y=3.215 $X2=0.26 $Y2=3.07
cc_143 N_VDD_c_99_p N_S_c_593_n 0.00435496f $X=3.74 $Y=5.36 $X2=0.26 $Y2=3.07
cc_144 N_VDD_M1009_b S 0.0096041f $X=-0.045 $Y=2.645 $X2=0.25 $Y2=2.125
cc_145 N_VDD_M1009_b N_S_c_598_n 0.0102428f $X=-0.045 $Y=2.645 $X2=0.26 $Y2=3.07
cc_146 N_VDD_c_98_p N_S_c_598_n 0.00528993f $X=0.75 $Y=3.215 $X2=0.26 $Y2=3.07
cc_147 N_VDD_M1009_b N_CO_c_624_n 0.00274939f $X=-0.045 $Y=2.645 $X2=2.1
+ $Y2=3.215
cc_148 N_VDD_c_101_p N_CO_c_624_n 0.00475705f $X=2.965 $Y=5.397 $X2=2.1
+ $Y2=3.215
cc_149 N_VDD_c_99_p N_CO_c_624_n 0.00435496f $X=3.74 $Y=5.36 $X2=2.1 $Y2=3.215
cc_150 N_VDD_M1009_b N_CO_c_621_n 0.00360959f $X=-0.045 $Y=2.645 $X2=2.175
+ $Y2=2.7
cc_151 N_VDD_M1009_b CO 0.0105263f $X=-0.045 $Y=2.645 $X2=2.175 $Y2=2.7
cc_152 N_CON_M1006_g N_B_M1007_g 0.0378719f $X=0.475 $Y=0.895 $X2=0.965
+ $Y2=0.895
cc_153 N_CON_c_158_n N_B_M1007_g 0.00317949f $X=0.635 $Y=1.59 $X2=0.965
+ $Y2=0.895
cc_154 N_CON_c_167_n N_B_M1007_g 0.0103705f $X=2.475 $Y=1.59 $X2=0.965 $Y2=0.895
cc_155 N_CON_c_169_n N_B_M1007_g 9.80511e-19 $X=0.78 $Y=1.59 $X2=0.965 $Y2=0.895
cc_156 N_CON_M1009_g N_B_M1011_g 0.0620831f $X=0.475 $Y=3.825 $X2=0.965
+ $Y2=3.825
cc_157 N_CON_c_161_n N_B_M1004_g 0.00298059f $X=2.62 $Y=2.605 $X2=3.205
+ $Y2=0.995
cc_158 N_CON_c_162_n N_B_M1004_g 0.0120887f $X=3.335 $Y=1.59 $X2=3.205 $Y2=0.995
cc_159 N_CON_c_165_n N_B_M1004_g 0.00288927f $X=3.42 $Y=1.065 $X2=3.205
+ $Y2=0.995
cc_160 N_CON_c_171_n N_B_M1004_g 4.76806e-19 $X=2.62 $Y=1.59 $X2=3.205 $Y2=0.995
cc_161 CON N_B_M1004_g 0.00638136f $X=3.42 $Y=1.59 $X2=3.205 $Y2=0.995
cc_162 N_CON_c_161_n N_B_M1013_g 0.00509671f $X=2.62 $Y=2.605 $X2=3.265
+ $Y2=3.825
cc_163 N_CON_c_163_n N_B_M1013_g 0.0160357f $X=3.755 $Y=2.69 $X2=3.265 $Y2=3.825
cc_164 N_CON_M1009_g N_B_c_289_n 0.0198105f $X=0.475 $Y=3.825 $X2=0.905 $Y2=1.96
cc_165 N_CON_c_167_n N_B_c_289_n 0.0017113f $X=2.475 $Y=1.59 $X2=0.905 $Y2=1.96
cc_166 N_CON_c_161_n N_B_c_291_n 0.00527976f $X=2.62 $Y=2.605 $X2=3.205 $Y2=1.96
cc_167 N_CON_c_162_n N_B_c_291_n 0.00297725f $X=3.335 $Y=1.59 $X2=3.205 $Y2=1.96
cc_168 N_CON_c_163_n N_B_c_291_n 0.00235541f $X=3.755 $Y=2.69 $X2=3.205 $Y2=1.96
cc_169 CON N_B_c_291_n 0.00117979f $X=3.42 $Y=1.59 $X2=3.205 $Y2=1.96
cc_170 N_CON_M1009_g N_B_c_292_n 0.00376362f $X=0.475 $Y=3.825 $X2=0.905
+ $Y2=1.96
cc_171 N_CON_c_167_n N_B_c_292_n 0.00349538f $X=2.475 $Y=1.59 $X2=0.905 $Y2=1.96
cc_172 N_CON_c_169_n N_B_c_292_n 7.89715e-19 $X=0.78 $Y=1.59 $X2=0.905 $Y2=1.96
cc_173 N_CON_c_161_n N_B_c_294_n 0.00612449f $X=2.62 $Y=2.605 $X2=3.205 $Y2=1.96
cc_174 N_CON_c_162_n N_B_c_294_n 0.0159093f $X=3.335 $Y=1.59 $X2=3.205 $Y2=1.96
cc_175 N_CON_c_163_n N_B_c_294_n 0.00416532f $X=3.755 $Y=2.69 $X2=3.205 $Y2=1.96
cc_176 N_CON_c_164_n N_B_c_294_n 0.00205373f $X=3.42 $Y=1.505 $X2=3.205 $Y2=1.96
cc_177 CON N_B_c_294_n 9.81883e-19 $X=3.42 $Y=1.59 $X2=3.205 $Y2=1.96
cc_178 N_CON_M1009_g N_B_c_295_n 3.21736e-19 $X=0.475 $Y=3.825 $X2=1.05 $Y2=1.96
cc_179 N_CON_c_167_n N_B_c_295_n 0.024704f $X=2.475 $Y=1.59 $X2=1.05 $Y2=1.96
cc_180 N_CON_c_169_n N_B_c_295_n 0.00206194f $X=0.78 $Y=1.59 $X2=1.05 $Y2=1.96
cc_181 N_CON_c_161_n N_B_c_296_n 0.0139114f $X=2.62 $Y=2.605 $X2=3.06 $Y2=1.96
cc_182 N_CON_c_162_n N_B_c_296_n 0.0132985f $X=3.335 $Y=1.59 $X2=3.06 $Y2=1.96
cc_183 N_CON_c_167_n N_B_c_296_n 0.116608f $X=2.475 $Y=1.59 $X2=3.06 $Y2=1.96
cc_184 N_CON_c_171_n N_B_c_296_n 0.0254758f $X=2.62 $Y=1.59 $X2=3.06 $Y2=1.96
cc_185 N_CON_c_161_n B 0.00223952f $X=2.62 $Y=2.605 $X2=3.21 $Y2=1.96
cc_186 N_CON_c_162_n B 0.00321159f $X=3.335 $Y=1.59 $X2=3.21 $Y2=1.96
cc_187 CON B 0.0176994f $X=3.42 $Y=1.59 $X2=3.21 $Y2=1.96
cc_188 N_CON_c_167_n N_A_M1008_g 0.0102813f $X=2.475 $Y=1.59 $X2=1.325 $Y2=0.895
cc_189 N_CON_c_163_n N_A_M1000_g 0.015762f $X=3.755 $Y=2.69 $X2=3.625 $Y2=3.825
cc_190 N_CON_c_183_n N_A_M1000_g 0.00669003f $X=3.84 $Y=3.215 $X2=3.625
+ $Y2=3.825
cc_191 N_CON_c_164_n N_A_M1005_g 0.00402015f $X=3.42 $Y=1.505 $X2=3.635
+ $Y2=0.995
cc_192 N_CON_c_165_n N_A_M1005_g 0.00288927f $X=3.42 $Y=1.065 $X2=3.635
+ $Y2=0.995
cc_193 CON N_A_M1005_g 0.010636f $X=3.42 $Y=1.59 $X2=3.635 $Y2=0.995
cc_194 N_CON_c_163_n N_A_c_391_n 0.00303009f $X=3.755 $Y=2.69 $X2=3.685 $Y2=2.33
cc_195 N_CON_c_163_n N_A_c_393_n 0.0189273f $X=3.755 $Y=2.69 $X2=3.685 $Y2=2.33
cc_196 CON N_A_c_393_n 3.86961e-19 $X=3.42 $Y=1.59 $X2=3.685 $Y2=2.33
cc_197 N_CON_c_163_n A 0.00711502f $X=3.755 $Y=2.69 $X2=3.685 $Y2=2.33
cc_198 CON A 0.00132366f $X=3.42 $Y=1.59 $X2=3.685 $Y2=2.33
cc_199 N_CON_c_161_n N_A_c_396_n 0.0228953f $X=2.62 $Y=2.605 $X2=3.54 $Y2=2.33
cc_200 N_CON_c_163_n N_A_c_396_n 0.0305931f $X=3.755 $Y=2.69 $X2=3.54 $Y2=2.33
cc_201 N_CON_c_164_n N_A_c_396_n 8.38986e-19 $X=3.42 $Y=1.505 $X2=3.54 $Y2=2.33
cc_202 CON N_A_c_396_n 0.0098042f $X=3.42 $Y=1.59 $X2=3.54 $Y2=2.33
cc_203 N_CON_c_167_n N_A_208_565#_c_470_n 0.0103748f $X=2.475 $Y=1.59 $X2=1.885
+ $Y2=1.86
cc_204 N_CON_c_167_n N_A_208_565#_c_473_n 0.00225837f $X=2.475 $Y=1.59 $X2=2.21
+ $Y2=1.565
cc_205 N_CON_c_161_n N_A_208_565#_c_474_n 0.0141245f $X=2.62 $Y=2.605 $X2=2.76
+ $Y2=2.41
cc_206 N_CON_c_162_n N_A_208_565#_c_474_n 0.00257529f $X=3.335 $Y=1.59 $X2=2.76
+ $Y2=2.41
cc_207 N_CON_c_171_n N_A_208_565#_c_475_n 2.41495e-19 $X=2.62 $Y=1.59 $X2=2.285
+ $Y2=1.49
cc_208 N_CON_c_160_n N_A_208_565#_c_479_n 0.00929899f $X=2.62 $Y=1.675 $X2=2.7
+ $Y2=1.565
cc_209 N_CON_c_162_n N_A_208_565#_c_479_n 0.0101401f $X=3.335 $Y=1.59 $X2=2.7
+ $Y2=1.565
cc_210 N_CON_c_167_n N_A_208_565#_c_479_n 0.00553403f $X=2.475 $Y=1.59 $X2=2.7
+ $Y2=1.565
cc_211 N_CON_c_171_n N_A_208_565#_c_479_n 0.00162604f $X=2.62 $Y=1.59 $X2=2.7
+ $Y2=1.565
cc_212 N_CON_c_171_n N_A_208_565#_c_481_n 0.00294886f $X=2.62 $Y=1.59 $X2=2.775
+ $Y2=1.49
cc_213 N_CON_c_161_n N_A_208_565#_M1003_g 0.0046186f $X=2.62 $Y=2.605 $X2=2.835
+ $Y2=3.825
cc_214 N_CON_c_178_n N_A_208_565#_M1003_g 0.00669003f $X=2.62 $Y=3.215 $X2=2.835
+ $Y2=3.825
cc_215 N_CON_c_163_n N_A_208_565#_M1003_g 0.0162813f $X=3.755 $Y=2.69 $X2=2.835
+ $Y2=3.825
cc_216 N_CON_c_167_n N_A_208_565#_c_486_n 0.00467421f $X=2.475 $Y=1.59 $X2=2.285
+ $Y2=1.565
cc_217 N_CON_c_167_n N_A_208_565#_c_487_n 0.0108903f $X=2.475 $Y=1.59 $X2=1.54
+ $Y2=0.885
cc_218 N_CON_c_167_n N_A_208_565#_c_492_n 0.0233954f $X=2.475 $Y=1.59 $X2=1.725
+ $Y2=1.695
cc_219 N_CON_M1006_g N_S_c_586_n 0.00716144f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=0.885
cc_220 N_CON_c_157_n N_S_c_586_n 0.00243007f $X=0.35 $Y=1.59 $X2=0.26 $Y2=0.885
cc_221 N_CON_c_158_n N_S_c_586_n 0.00919709f $X=0.635 $Y=1.59 $X2=0.26 $Y2=0.885
cc_222 N_CON_M1009_g N_S_c_593_n 0.00485682f $X=0.475 $Y=3.825 $X2=0.26 $Y2=3.07
cc_223 N_CON_M1006_g S 0.00219688f $X=0.475 $Y=0.895 $X2=0.25 $Y2=2.125
cc_224 N_CON_M1009_g S 0.026126f $X=0.475 $Y=3.825 $X2=0.25 $Y2=2.125
cc_225 N_CON_c_157_n S 0.0074247f $X=0.35 $Y=1.59 $X2=0.25 $Y2=2.125
cc_226 N_CON_c_158_n S 0.0144314f $X=0.635 $Y=1.59 $X2=0.25 $Y2=2.125
cc_227 N_CON_c_169_n S 0.0220567f $X=0.78 $Y=1.59 $X2=0.25 $Y2=2.125
cc_228 N_CON_M1006_g N_S_c_591_n 0.00595114f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=1.215
cc_229 N_CON_c_157_n N_S_c_591_n 0.00148757f $X=0.35 $Y=1.59 $X2=0.26 $Y2=1.215
cc_230 N_CON_c_158_n N_S_c_591_n 0.00260285f $X=0.635 $Y=1.59 $X2=0.26 $Y2=1.215
cc_231 N_CON_M1009_g N_S_c_598_n 0.00321348f $X=0.475 $Y=3.825 $X2=0.26 $Y2=3.07
cc_232 N_CON_c_178_n N_CO_c_624_n 0.0867869f $X=2.62 $Y=3.215 $X2=2.1 $Y2=3.215
cc_233 N_CON_c_167_n N_CO_c_620_n 0.00532638f $X=2.475 $Y=1.59 $X2=2.175
+ $Y2=1.25
cc_234 N_CON_c_178_n N_CO_c_621_n 3.73019e-19 $X=2.62 $Y=3.215 $X2=2.175 $Y2=2.7
cc_235 N_CON_c_160_n N_CO_c_622_n 0.00670709f $X=2.62 $Y=1.675 $X2=2.137
+ $Y2=2.615
cc_236 N_CON_c_161_n N_CO_c_622_n 0.0448782f $X=2.62 $Y=2.605 $X2=2.137
+ $Y2=2.615
cc_237 N_CON_c_166_n N_CO_c_622_n 0.00730853f $X=2.62 $Y=2.69 $X2=2.137
+ $Y2=2.615
cc_238 N_CON_c_167_n N_CO_c_622_n 0.0120817f $X=2.475 $Y=1.59 $X2=2.137
+ $Y2=2.615
cc_239 N_CON_c_171_n N_CO_c_622_n 0.00207393f $X=2.62 $Y=1.59 $X2=2.137
+ $Y2=2.615
cc_240 N_CON_c_161_n CO 5.70376e-19 $X=2.62 $Y=2.605 $X2=2.175 $Y2=2.7
cc_241 N_CON_c_178_n CO 0.00122973f $X=2.62 $Y=3.215 $X2=2.175 $Y2=2.7
cc_242 N_CON_c_166_n CO 0.00605606f $X=2.62 $Y=2.69 $X2=2.175 $Y2=2.7
cc_243 N_CON_c_162_n N_A_570_115#_c_673_n 0.0101003f $X=3.335 $Y=1.59 $X2=2.99
+ $Y2=0.74
cc_244 N_CON_M1004_d N_A_570_115#_c_668_n 0.00176461f $X=3.28 $Y=0.575 $X2=3.765
+ $Y2=0.56
cc_245 N_CON_c_165_n N_A_570_115#_c_668_n 0.0130031f $X=3.42 $Y=1.065 $X2=3.765
+ $Y2=0.56
cc_246 N_B_M1007_g N_A_M1008_g 0.0639188f $X=0.965 $Y=0.895 $X2=1.325 $Y2=0.895
cc_247 N_B_c_292_n N_A_M1008_g 0.00121678f $X=0.905 $Y=1.96 $X2=1.325 $Y2=0.895
cc_248 N_B_c_295_n N_A_M1008_g 7.94897e-19 $X=1.05 $Y=1.96 $X2=1.325 $Y2=0.895
cc_249 N_B_c_296_n N_A_M1008_g 0.00595709f $X=3.06 $Y=1.96 $X2=1.325 $Y2=0.895
cc_250 N_B_M1011_g N_A_M1012_g 0.0405421f $X=0.965 $Y=3.825 $X2=1.395 $Y2=3.825
cc_251 N_B_M1004_g N_A_M1005_g 0.0414265f $X=3.205 $Y=0.995 $X2=3.635 $Y2=0.995
cc_252 N_B_c_291_n N_A_M1005_g 0.022402f $X=3.205 $Y=1.96 $X2=3.635 $Y2=0.995
cc_253 N_B_c_294_n N_A_M1005_g 0.00376362f $X=3.205 $Y=1.96 $X2=3.635 $Y2=0.995
cc_254 B N_A_M1005_g 9.23221e-19 $X=3.21 $Y=1.96 $X2=3.635 $Y2=0.995
cc_255 N_B_c_289_n N_A_c_390_n 0.0639188f $X=0.905 $Y=1.96 $X2=1.385 $Y2=2.33
cc_256 N_B_c_296_n N_A_c_390_n 7.99243e-19 $X=3.06 $Y=1.96 $X2=1.385 $Y2=2.33
cc_257 N_B_M1013_g N_A_c_391_n 0.168643f $X=3.265 $Y=3.825 $X2=3.685 $Y2=2.33
cc_258 N_B_M1011_g N_A_c_392_n 0.00286993f $X=0.965 $Y=3.825 $X2=1.385 $Y2=2.33
cc_259 N_B_c_296_n N_A_c_392_n 0.00428104f $X=3.06 $Y=1.96 $X2=1.385 $Y2=2.33
cc_260 N_B_M1013_g N_A_c_393_n 0.00278747f $X=3.265 $Y=3.825 $X2=3.685 $Y2=2.33
cc_261 N_B_M1011_g N_A_c_394_n 0.00405562f $X=0.965 $Y=3.825 $X2=1.53 $Y2=2.33
cc_262 N_B_c_296_n N_A_c_394_n 0.0263377f $X=3.06 $Y=1.96 $X2=1.53 $Y2=2.33
cc_263 N_B_M1013_g A 7.94897e-19 $X=3.265 $Y=3.825 $X2=3.685 $Y2=2.33
cc_264 N_B_M1013_g N_A_c_396_n 0.00633265f $X=3.265 $Y=3.825 $X2=3.54 $Y2=2.33
cc_265 N_B_c_291_n N_A_c_396_n 0.00210214f $X=3.205 $Y=1.96 $X2=3.54 $Y2=2.33
cc_266 N_B_c_294_n N_A_c_396_n 0.00225835f $X=3.205 $Y=1.96 $X2=3.54 $Y2=2.33
cc_267 N_B_c_296_n N_A_c_396_n 0.128931f $X=3.06 $Y=1.96 $X2=3.54 $Y2=2.33
cc_268 B N_A_c_396_n 0.0270107f $X=3.21 $Y=1.96 $X2=3.54 $Y2=2.33
cc_269 N_B_c_296_n N_A_208_565#_c_471_n 0.00725075f $X=3.06 $Y=1.96 $X2=1.885
+ $Y2=2.335
cc_270 N_B_c_296_n N_A_208_565#_c_473_n 0.00119779f $X=3.06 $Y=1.96 $X2=2.21
+ $Y2=1.565
cc_271 N_B_M1013_g N_A_208_565#_c_474_n 0.0381911f $X=3.265 $Y=3.825 $X2=2.76
+ $Y2=2.41
cc_272 N_B_c_296_n N_A_208_565#_c_474_n 0.00176131f $X=3.06 $Y=1.96 $X2=2.76
+ $Y2=2.41
cc_273 N_B_M1004_g N_A_208_565#_c_481_n 0.022187f $X=3.205 $Y=0.995 $X2=2.775
+ $Y2=1.49
cc_274 N_B_M1011_g N_A_208_565#_c_507_n 0.00507079f $X=0.965 $Y=3.825 $X2=1.265
+ $Y2=2.75
cc_275 N_B_c_296_n N_A_208_565#_c_507_n 0.0051538f $X=3.06 $Y=1.96 $X2=1.265
+ $Y2=2.75
cc_276 N_B_c_292_n N_A_208_565#_c_491_n 0.00316158f $X=0.905 $Y=1.96 $X2=1.725
+ $Y2=2.665
cc_277 N_B_c_295_n N_A_208_565#_c_491_n 0.00129846f $X=1.05 $Y=1.96 $X2=1.725
+ $Y2=2.665
cc_278 N_B_c_296_n N_A_208_565#_c_491_n 0.0153226f $X=3.06 $Y=1.96 $X2=1.725
+ $Y2=2.665
cc_279 N_B_c_295_n N_A_208_565#_c_492_n 5.15761e-19 $X=1.05 $Y=1.96 $X2=1.725
+ $Y2=1.695
cc_280 N_B_c_296_n N_A_208_565#_c_492_n 0.00890945f $X=3.06 $Y=1.96 $X2=1.725
+ $Y2=1.695
cc_281 N_B_M1007_g S 4.21151e-19 $X=0.965 $Y=0.895 $X2=0.25 $Y2=2.125
cc_282 N_B_c_292_n S 0.00429487f $X=0.905 $Y=1.96 $X2=0.25 $Y2=2.125
cc_283 N_B_c_295_n S 0.0134542f $X=1.05 $Y=1.96 $X2=0.25 $Y2=2.125
cc_284 N_B_M1007_g N_S_c_591_n 3.7658e-19 $X=0.965 $Y=0.895 $X2=0.26 $Y2=1.215
cc_285 N_B_c_296_n N_CO_c_622_n 0.0136433f $X=3.06 $Y=1.96 $X2=2.137 $Y2=2.615
cc_286 N_B_M1004_g N_A_570_115#_c_668_n 0.012637f $X=3.205 $Y=0.995 $X2=3.765
+ $Y2=0.56
cc_287 N_A_M1008_g N_A_208_565#_c_470_n 0.0166096f $X=1.325 $Y=0.895 $X2=1.885
+ $Y2=1.86
cc_288 N_A_M1008_g N_A_208_565#_c_471_n 0.00833244f $X=1.325 $Y=0.895 $X2=1.885
+ $Y2=2.335
cc_289 N_A_c_390_n N_A_208_565#_c_471_n 0.0147848f $X=1.385 $Y=2.33 $X2=1.885
+ $Y2=2.335
cc_290 N_A_c_396_n N_A_208_565#_c_471_n 0.00210973f $X=3.54 $Y=2.33 $X2=1.885
+ $Y2=2.335
cc_291 N_A_M1012_g N_A_208_565#_M1002_g 0.0513848f $X=1.395 $Y=3.825 $X2=1.885
+ $Y2=3.825
cc_292 N_A_c_396_n N_A_208_565#_c_474_n 0.0139241f $X=3.54 $Y=2.33 $X2=2.76
+ $Y2=2.41
cc_293 N_A_c_396_n N_A_208_565#_c_485_n 0.00700381f $X=3.54 $Y=2.33 $X2=1.885
+ $Y2=2.41
cc_294 N_A_M1012_g N_A_208_565#_c_504_n 0.0147914f $X=1.395 $Y=3.825 $X2=1.64
+ $Y2=2.75
cc_295 N_A_c_390_n N_A_208_565#_c_504_n 0.00348735f $X=1.385 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_296 N_A_c_392_n N_A_208_565#_c_504_n 0.0111584f $X=1.385 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_297 N_A_c_394_n N_A_208_565#_c_504_n 0.00509311f $X=1.53 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_298 N_A_c_396_n N_A_208_565#_c_504_n 0.00467069f $X=3.54 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_299 N_A_c_390_n N_A_208_565#_c_507_n 7.25782e-19 $X=1.385 $Y=2.33 $X2=1.265
+ $Y2=2.75
cc_300 N_A_c_394_n N_A_208_565#_c_507_n 0.00124978f $X=1.53 $Y=2.33 $X2=1.265
+ $Y2=2.75
cc_301 N_A_M1008_g N_A_208_565#_c_487_n 0.0155978f $X=1.325 $Y=0.895 $X2=1.54
+ $Y2=0.885
cc_302 N_A_M1008_g N_A_208_565#_c_491_n 0.00392362f $X=1.325 $Y=0.895 $X2=1.725
+ $Y2=2.665
cc_303 N_A_M1012_g N_A_208_565#_c_491_n 0.00360042f $X=1.395 $Y=3.825 $X2=1.725
+ $Y2=2.665
cc_304 N_A_c_390_n N_A_208_565#_c_491_n 0.00193142f $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_305 N_A_c_392_n N_A_208_565#_c_491_n 0.0224238f $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_306 N_A_c_394_n N_A_208_565#_c_491_n 0.00168305f $X=1.53 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_307 N_A_c_396_n N_A_208_565#_c_491_n 0.0185059f $X=3.54 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_308 N_A_M1008_g N_A_208_565#_c_492_n 0.00736605f $X=1.325 $Y=0.895 $X2=1.725
+ $Y2=1.695
cc_309 N_A_c_390_n N_A_208_565#_c_492_n 0.00175929f $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=1.695
cc_310 N_A_c_392_n N_A_208_565#_c_492_n 2.52704e-19 $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=1.695
cc_311 N_A_c_396_n N_CO_c_621_n 0.00105312f $X=3.54 $Y=2.33 $X2=2.175 $Y2=2.7
cc_312 N_A_c_396_n N_CO_c_622_n 0.0133702f $X=3.54 $Y=2.33 $X2=2.137 $Y2=2.615
cc_313 N_A_c_396_n CO 0.0346374f $X=3.54 $Y=2.33 $X2=2.175 $Y2=2.7
cc_314 N_A_M1005_g N_A_570_115#_c_668_n 0.0135957f $X=3.635 $Y=0.995 $X2=3.765
+ $Y2=0.56
cc_315 N_A_208_565#_c_487_n N_CO_c_617_n 0.0246852f $X=1.54 $Y=0.885 $X2=2.07
+ $Y2=0.74
cc_316 N_A_208_565#_c_473_n N_CO_c_620_n 0.00430718f $X=2.21 $Y=1.565 $X2=2.175
+ $Y2=1.25
cc_317 N_A_208_565#_c_475_n N_CO_c_620_n 0.00630936f $X=2.285 $Y=1.49 $X2=2.175
+ $Y2=1.25
cc_318 N_A_208_565#_c_481_n N_CO_c_620_n 3.96157e-19 $X=2.775 $Y=1.49 $X2=2.175
+ $Y2=1.25
cc_319 N_A_208_565#_c_487_n N_CO_c_620_n 0.00748803f $X=1.54 $Y=0.885 $X2=2.175
+ $Y2=1.25
cc_320 N_A_208_565#_M1002_g N_CO_c_621_n 0.00954321f $X=1.885 $Y=3.825 $X2=2.175
+ $Y2=2.7
cc_321 N_A_208_565#_c_474_n N_CO_c_621_n 0.00140819f $X=2.76 $Y=2.41 $X2=2.175
+ $Y2=2.7
cc_322 N_A_208_565#_c_504_n N_CO_c_621_n 0.0104146f $X=1.64 $Y=2.75 $X2=2.175
+ $Y2=2.7
cc_323 N_A_208_565#_c_491_n N_CO_c_621_n 0.00298908f $X=1.725 $Y=2.665 $X2=2.175
+ $Y2=2.7
cc_324 N_A_208_565#_c_470_n N_CO_c_622_n 0.0106736f $X=1.885 $Y=1.86 $X2=2.137
+ $Y2=2.615
cc_325 N_A_208_565#_M1002_g N_CO_c_622_n 0.00273706f $X=1.885 $Y=3.825 $X2=2.137
+ $Y2=2.615
cc_326 N_A_208_565#_c_473_n N_CO_c_622_n 0.00779052f $X=2.21 $Y=1.565 $X2=2.137
+ $Y2=2.615
cc_327 N_A_208_565#_c_474_n N_CO_c_622_n 0.0137108f $X=2.76 $Y=2.41 $X2=2.137
+ $Y2=2.615
cc_328 N_A_208_565#_c_475_n N_CO_c_622_n 0.00543017f $X=2.285 $Y=1.49 $X2=2.137
+ $Y2=2.615
cc_329 N_A_208_565#_c_481_n N_CO_c_622_n 7.59428e-19 $X=2.775 $Y=1.49 $X2=2.137
+ $Y2=2.615
cc_330 N_A_208_565#_M1003_g N_CO_c_622_n 8.14457e-19 $X=2.835 $Y=3.825 $X2=2.137
+ $Y2=2.615
cc_331 N_A_208_565#_c_486_n N_CO_c_622_n 0.0035441f $X=2.285 $Y=1.565 $X2=2.137
+ $Y2=2.615
cc_332 N_A_208_565#_c_487_n N_CO_c_622_n 0.00671312f $X=1.54 $Y=0.885 $X2=2.137
+ $Y2=2.615
cc_333 N_A_208_565#_c_491_n N_CO_c_622_n 0.0354244f $X=1.725 $Y=2.665 $X2=2.137
+ $Y2=2.615
cc_334 N_A_208_565#_c_492_n N_CO_c_622_n 0.0222011f $X=1.725 $Y=1.695 $X2=2.137
+ $Y2=2.615
cc_335 N_A_208_565#_M1002_g CO 7.58429e-19 $X=1.885 $Y=3.825 $X2=2.175 $Y2=2.7
cc_336 N_A_208_565#_c_474_n CO 0.0027071f $X=2.76 $Y=2.41 $X2=2.175 $Y2=2.7
cc_337 N_A_208_565#_c_504_n CO 0.00111652f $X=1.64 $Y=2.75 $X2=2.175 $Y2=2.7
cc_338 N_A_208_565#_c_491_n CO 0.0012063f $X=1.725 $Y=2.665 $X2=2.175 $Y2=2.7
cc_339 N_A_208_565#_c_481_n N_A_570_115#_c_670_n 9.82882e-19 $X=2.775 $Y=1.49
+ $X2=3.075 $Y2=0.56
