* File: sky130_osu_sc_18T_hs__dffs_l.pex.spice
* Created: Thu Oct 29 17:07:45 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%GND 1 2 3 4 5 6 67 71 77 79 89 91 101
+ 103 113 115 122 126 142 144
c192 101 0 1.67294e-19 $X=5.14 $Y=0.825
c193 77 0 3.07193e-19 $X=1.64 $Y=0.825
c194 67 0 1.27355e-19 $X=-0.05 $Y=0
r195 142 144 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=7.815 $Y2=0.152
r196 120 122 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.825
r197 116 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=0.152
+ $X2=6.88 $Y2=0.152
r198 111 137 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.152
r199 111 113 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.825
r200 103 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=0.152
+ $X2=6.88 $Y2=0.152
r201 99 101 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.14 $Y=0.305
+ $X2=5.14 $Y2=0.825
r202 92 133 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.152
+ $X2=3.39 $Y2=0.152
r203 87 133 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.152
r204 87 89 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.825
r205 79 133 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.152
+ $X2=3.39 $Y2=0.152
r206 75 77 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.64 $Y=0.305
+ $X2=1.64 $Y2=0.825
r207 73 74 15.8697 $w=3.03e-07 $l=4.2e-07 $layer=LI1_cond $X=1.555 $Y=0.152
+ $X2=1.135 $Y2=0.152
r208 69 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r209 67 120 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r210 67 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r211 67 126 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=0.335 $Y=0.152
+ $X2=0.965 $Y2=0.152
r212 67 144 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=0.17
+ $X2=7.815 $Y2=0.17
r213 67 142 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=0.17
+ $X2=0.335 $Y2=0.17
r214 67 99 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.14 $Y2=0.305
r215 67 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.055 $Y2=0.152
r216 67 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.225 $Y2=0.152
r217 67 75 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.64 $Y2=0.305
r218 67 73 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.555 $Y2=0.152
r219 67 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.725 $Y2=0.152
r220 67 69 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r221 67 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r222 67 74 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r223 67 115 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r224 67 116 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.965 $Y2=0.152
r225 67 103 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.795 $Y2=0.152
r226 67 104 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=5.225 $Y2=0.152
r227 67 91 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=5.055 $Y2=0.152
r228 67 92 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.475 $Y2=0.152
r229 67 79 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=3.305 $Y2=0.152
r230 67 80 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=1.725 $Y2=0.152
r231 6 122 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.825
r232 5 113 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.575 $X2=6.88 $Y2=0.825
r233 4 101 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5
+ $Y=0.575 $X2=5.14 $Y2=0.825
r234 3 89 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.575 $X2=3.39 $Y2=0.825
r235 2 77 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.575 $X2=1.64 $Y2=0.825
r236 1 71 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%VDD 1 2 3 4 5 6 7 8 61 65 69 75 83 87 95
+ 99 107 111 117 121 127 131 137 152 157 158
r105 157 158 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=6.49
+ $X2=7.815 $Y2=6.49
r106 152 157 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=6.507
+ $X2=7.815 $Y2=6.507
r107 152 155 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=6.49
+ $X2=0.335 $Y2=6.49
r108 137 140 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.9 $Y=4.475
+ $X2=7.9 $Y2=5.835
r109 135 158 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=6.507
r110 135 140 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=5.835
r111 132 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.035 $Y=6.507
+ $X2=6.95 $Y2=6.507
r112 132 134 3.7785 $w=3.03e-07 $l=1e-07 $layer=LI1_cond $X=7.035 $Y=6.507
+ $X2=7.135 $Y2=6.507
r113 131 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.9 $Y2=6.507
r114 131 134 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.135 $Y2=6.507
r115 127 130 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.95 $Y=4.815
+ $X2=6.95 $Y2=5.835
r116 125 150 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.95 $Y=6.355
+ $X2=6.95 $Y2=6.507
r117 125 130 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.95 $Y=6.355
+ $X2=6.95 $Y2=5.835
r118 122 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.09 $Y2=6.507
r119 122 124 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.455 $Y2=6.507
r120 121 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=6.507
+ $X2=6.95 $Y2=6.507
r121 121 124 15.4919 $w=3.03e-07 $l=4.1e-07 $layer=LI1_cond $X=6.865 $Y=6.507
+ $X2=6.455 $Y2=6.507
r122 117 120 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.09 $Y=4.815
+ $X2=6.09 $Y2=5.835
r123 115 149 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=6.507
r124 115 120 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=5.835
r125 112 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.14 $Y2=6.507
r126 112 114 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.775 $Y2=6.507
r127 111 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=6.09 $Y2=6.507
r128 111 114 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=5.775 $Y2=6.507
r129 107 110 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.14 $Y=3.455
+ $X2=5.14 $Y2=5.835
r130 105 148 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.14 $Y=6.355
+ $X2=5.14 $Y2=6.507
r131 105 110 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.14 $Y=6.355
+ $X2=5.14 $Y2=5.835
r132 102 104 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=6.507
+ $X2=4.415 $Y2=6.507
r133 100 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=6.507
+ $X2=3.39 $Y2=6.507
r134 100 102 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.475 $Y=6.507
+ $X2=3.735 $Y2=6.507
r135 99 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=6.507
+ $X2=5.14 $Y2=6.507
r136 99 104 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=5.055 $Y=6.507
+ $X2=4.415 $Y2=6.507
r137 95 98 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=3.39 $Y=3.795
+ $X2=3.39 $Y2=5.835
r138 93 146 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.39 $Y=6.355
+ $X2=3.39 $Y2=6.507
r139 93 98 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=6.355
+ $X2=3.39 $Y2=5.835
r140 90 92 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.375 $Y=6.507
+ $X2=3.055 $Y2=6.507
r141 88 145 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=6.507
+ $X2=1.64 $Y2=6.507
r142 88 90 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=1.725 $Y=6.507
+ $X2=2.375 $Y2=6.507
r143 87 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=6.507
+ $X2=3.39 $Y2=6.507
r144 87 92 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.305 $Y=6.507
+ $X2=3.055 $Y2=6.507
r145 83 86 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.64 $Y=3.795
+ $X2=1.64 $Y2=5.835
r146 81 145 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.64 $Y=6.355
+ $X2=1.64 $Y2=6.507
r147 81 86 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.64 $Y=6.355
+ $X2=1.64 $Y2=5.835
r148 80 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r149 79 145 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=6.507
+ $X2=1.64 $Y2=6.507
r150 79 80 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=1.555 $Y=6.507
+ $X2=1.205 $Y2=6.507
r151 75 78 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=4.815
+ $X2=1.12 $Y2=5.835
r152 73 143 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r153 73 78 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r154 70 155 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r155 70 72 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.015 $Y2=6.507
r156 69 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r157 69 72 0.7557 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.015 $Y2=6.507
r158 65 68 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=4.815
+ $X2=0.26 $Y2=5.835
r159 63 155 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r160 63 68 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r161 61 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=6.355 $X2=7.815 $Y2=6.44
r162 61 155 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=6.355 $X2=0.335 $Y2=6.44
r163 61 148 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=6.355 $X2=5.095 $Y2=6.44
r164 61 145 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=6.355 $X2=1.695 $Y2=6.44
r165 61 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=6.355 $X2=7.135 $Y2=6.44
r166 61 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=6.355 $X2=6.455 $Y2=6.44
r167 61 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=6.355 $X2=5.775 $Y2=6.44
r168 61 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=6.355 $X2=4.415 $Y2=6.44
r169 61 102 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=6.355 $X2=3.735 $Y2=6.44
r170 61 92 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=6.355 $X2=3.055 $Y2=6.44
r171 61 90 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=6.355 $X2=2.375 $Y2=6.44
r172 61 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=6.355 $X2=1.015 $Y2=6.44
r173 8 140 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=4.085 $X2=7.9 $Y2=5.835
r174 8 137 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=4.085 $X2=7.9 $Y2=4.475
r175 7 130 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=4.085 $X2=6.95 $Y2=5.835
r176 7 127 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=4.085 $X2=6.95 $Y2=4.815
r177 6 120 300 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=5.965
+ $Y=4.085 $X2=6.09 $Y2=5.835
r178 6 117 300 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=2 $X=5.965
+ $Y=4.085 $X2=6.09 $Y2=4.815
r179 5 110 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5
+ $Y=3.085 $X2=5.14 $Y2=5.835
r180 5 107 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5
+ $Y=3.085 $X2=5.14 $Y2=3.455
r181 4 98 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.25
+ $Y=3.085 $X2=3.39 $Y2=5.835
r182 4 95 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=3.25
+ $Y=3.085 $X2=3.39 $Y2=3.795
r183 3 86 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=1.515 $Y=3.085 $X2=1.64 $Y2=5.835
r184 3 83 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=1.515 $Y=3.085 $X2=1.64 $Y2=3.795
r185 2 78 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=5.835
r186 2 75 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=4.815
r187 1 68 300 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=5.835
r188 1 65 300 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=4.815
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%SN 3 7 9 11 14 16 17 19 22 25 26 30 34
r130 34 37 19.0665 $w=3.16e-07 $l=1.25e-07 $layer=POLY_cond $X=6.735 $Y=1.59
+ $X2=6.86 $Y2=1.59
r131 33 34 10.6772 $w=3.16e-07 $l=7e-08 $layer=POLY_cond $X=6.665 $Y=1.59
+ $X2=6.735 $Y2=1.59
r132 30 32 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.85
+ $X2=0.367 $Y2=2.015
r133 30 31 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.85
+ $X2=0.367 $Y2=1.685
r134 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.85 $X2=0.32 $Y2=1.85
r135 26 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.59 $X2=6.86 $Y2=1.59
r136 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.86 $Y=1.48
+ $X2=6.86 $Y2=1.48
r137 22 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.48
+ $X2=0.32 $Y2=1.85
r138 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=1.48
+ $X2=0.32 $Y2=1.48
r139 17 19 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.465 $Y=1.48
+ $X2=0.32 $Y2=1.48
r140 16 25 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.715 $Y=1.48
+ $X2=6.86 $Y2=1.48
r141 16 17 6.01801 $w=1.7e-07 $l=6.25e-06 $layer=MET1_cond $X=6.715 $Y=1.48
+ $X2=0.465 $Y2=1.48
r142 12 34 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.755
+ $X2=6.735 $Y2=1.59
r143 12 14 1707.51 $w=1.5e-07 $l=3.33e-06 $layer=POLY_cond $X=6.735 $Y=1.755
+ $X2=6.735 $Y2=5.085
r144 9 33 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.665 $Y=1.425
+ $X2=6.665 $Y2=1.59
r145 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.665 $Y=1.425
+ $X2=6.665 $Y2=0.945
r146 7 32 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=0.475 $Y=5.085
+ $X2=0.475 $Y2=2.015
r147 3 31 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=1.685
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%A_152_89# 1 2 9 13 18 19 20 21 22 23 25
+ 28 32 37
c86 37 0 1.71621e-19 $X=2.507 $Y=1.415
c87 20 0 1.29912e-19 $X=2.33 $Y=1.765
r88 38 40 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.835 $Y=2.305
+ $X2=0.905 $Y2=2.305
r89 36 37 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.507 $Y=1.245
+ $X2=2.507 $Y2=1.415
r90 32 34 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=2.515 $Y=3.455
+ $X2=2.515 $Y2=5.835
r91 30 32 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=2.515 $Y=3.27
+ $X2=2.515 $Y2=3.455
r92 28 36 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=2.515 $Y=0.825
+ $X2=2.515 $Y2=1.245
r93 25 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.415 $Y=1.68
+ $X2=2.415 $Y2=1.415
r94 22 30 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.345 $Y=3.185
+ $X2=2.515 $Y2=3.27
r95 22 23 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.345 $Y=3.185
+ $X2=1.115 $Y2=3.185
r96 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=1.765
+ $X2=2.415 $Y2=1.68
r97 20 21 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.33 $Y=1.765
+ $X2=1.115 $Y2=1.765
r98 19 40 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.03 $Y=2.305
+ $X2=0.905 $Y2=2.305
r99 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=2.305 $X2=1.03 $Y2=2.305
r100 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=3.1
+ $X2=1.115 $Y2=3.185
r101 16 18 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.03 $Y=3.1
+ $X2=1.03 $Y2=2.305
r102 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=1.85
+ $X2=1.115 $Y2=1.765
r103 15 18 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.03 $Y=1.85
+ $X2=1.03 $Y2=2.305
r104 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.47
+ $X2=0.905 $Y2=2.305
r105 11 13 1340.88 $w=1.5e-07 $l=2.615e-06 $layer=POLY_cond $X=0.905 $Y=2.47
+ $X2=0.905 $Y2=5.085
r106 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=2.14
+ $X2=0.835 $Y2=2.305
r107 7 9 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.835 $Y=2.14
+ $X2=0.835 $Y2=0.945
r108 2 34 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=2.29
+ $Y=3.085 $X2=2.515 $Y2=5.835
r109 2 32 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=2.29
+ $Y=3.085 $X2=2.515 $Y2=3.455
r110 1 28 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.575 $X2=2.515 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%D 3 7 10 12 16
c41 16 0 1.12321e-19 $X=1.915 $Y=2.22
c42 10 0 1.41836e-19 $X=1.915 $Y=2.22
r43 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=2.22
+ $X2=1.915 $Y2=2.385
r44 16 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=2.22
+ $X2=1.915 $Y2=2.055
r45 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=2.22 $X2=1.915 $Y2=2.22
r46 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.915 $Y=2.22
+ $X2=1.915 $Y2=2.22
r47 7 18 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=1.855 $Y=4.585
+ $X2=1.855 $Y2=2.385
r48 3 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.855 $Y=1.075
+ $X2=1.855 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%CK 3 7 10 13 17 18 20 23 24 25 26 30 31
+ 35 36 38 39 40 41 42 43 46 50 52 54 59 63 66 70
c218 63 0 1.29912e-19 $X=2.755 $Y=1.685
c219 59 0 1.41836e-19 $X=2.275 $Y=2.765
c220 39 0 6.79641e-20 $X=4.11 $Y=2.59
c221 30 0 1.98654e-19 $X=2.755 $Y=1.85
c222 26 0 1.86602e-19 $X=2.67 $Y=2.59
r223 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=2.765 $X2=5.5 $Y2=2.765
r224 70 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=2.765
+ $X2=4.505 $Y2=2.93
r225 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=2.765 $X2=4.505 $Y2=2.765
r226 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=2.765
+ $X2=2.275 $Y2=2.93
r227 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=2.765 $X2=2.275 $Y2=2.765
r228 54 74 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.5 $Y=2.59
+ $X2=5.5 $Y2=2.765
r229 52 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.5 $Y=2.59 $X2=5.5
+ $Y2=2.59
r230 50 69 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.505 $Y=2.59
+ $X2=4.505 $Y2=2.765
r231 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.505 $Y=2.59
+ $X2=4.505 $Y2=2.59
r232 46 58 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.275 $Y=2.59
+ $X2=2.275 $Y2=2.765
r233 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.275 $Y=2.59
+ $X2=2.275 $Y2=2.59
r234 43 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.65 $Y=2.59
+ $X2=4.505 $Y2=2.59
r235 42 52 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.355 $Y=2.59
+ $X2=5.5 $Y2=2.59
r236 42 43 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=5.355 $Y=2.59
+ $X2=4.65 $Y2=2.59
r237 41 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.42 $Y=2.59
+ $X2=2.275 $Y2=2.59
r238 40 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.36 $Y=2.59
+ $X2=4.505 $Y2=2.59
r239 40 41 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=4.36 $Y=2.59
+ $X2=2.42 $Y2=2.59
r240 38 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.59
+ $X2=4.505 $Y2=2.59
r241 38 39 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.42 $Y=2.59
+ $X2=4.11 $Y2=2.59
r242 36 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.85
+ $X2=4.025 $Y2=1.685
r243 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.85 $X2=4.025 $Y2=1.85
r244 33 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=2.505
+ $X2=4.11 $Y2=2.59
r245 33 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.025 $Y=2.505
+ $X2=4.025 $Y2=1.85
r246 31 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.85
+ $X2=2.755 $Y2=1.685
r247 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.85 $X2=2.755 $Y2=1.85
r248 28 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.755 $Y=2.505
+ $X2=2.755 $Y2=1.85
r249 27 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.59
+ $X2=2.275 $Y2=2.59
r250 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.67 $Y=2.59
+ $X2=2.755 $Y2=2.505
r251 26 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.67 $Y=2.59
+ $X2=2.36 $Y2=2.59
r252 24 25 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=5.382 $Y=1.685
+ $X2=5.382 $Y2=1.835
r253 23 75 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=5.41 $Y=2.6
+ $X2=5.457 $Y2=2.765
r254 23 25 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=5.41 $Y=2.6
+ $X2=5.41 $Y2=1.835
r255 18 75 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=5.355 $Y=2.93
+ $X2=5.457 $Y2=2.765
r256 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.355 $Y=2.93
+ $X2=5.355 $Y2=4.585
r257 17 24 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.355 $Y=1.075
+ $X2=5.355 $Y2=1.685
r258 13 72 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=4.565 $Y=4.585
+ $X2=4.565 $Y2=2.93
r259 10 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.965 $Y=1.075
+ $X2=3.965 $Y2=1.685
r260 7 63 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.815 $Y=1.075
+ $X2=2.815 $Y2=1.685
r261 3 61 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.215 $Y=4.585
+ $X2=2.215 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%A_27_115# 1 2 9 13 17 21 23 24 25 26 29
+ 31 32 35 39 40 43 46 47
c127 39 0 1.35571e-19 $X=3.11 $Y=1.85
c128 35 0 1.5821e-19 $X=3.345 $Y=2.765
c129 26 0 6.79641e-20 $X=3.53 $Y=2.765
c130 24 0 1.86602e-19 $X=3.25 $Y=2.765
c131 21 0 6.36774e-20 $X=3.605 $Y=4.585
c132 13 0 6.36774e-20 $X=3.175 $Y=4.585
r133 55 57 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=4.815
+ $X2=0.69 $Y2=5.835
r134 47 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.85 $X2=3.345 $Y2=1.85
r135 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.255 $Y=1.85
+ $X2=3.255 $Y2=1.85
r136 43 55 193.439 $w=1.68e-07 $l=2.965e-06 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=4.815
r137 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=1.85
r138 40 42 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.85
+ $X2=0.69 $Y2=1.85
r139 39 46 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.11 $Y=1.85
+ $X2=3.255 $Y2=1.85
r140 39 40 2.19056 $w=1.7e-07 $l=2.275e-06 $layer=MET1_cond $X=3.11 $Y=1.85
+ $X2=0.835 $Y2=1.85
r141 38 43 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.69 $Y=1.165
+ $X2=0.69 $Y2=1.85
r142 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=2.765 $X2=3.345 $Y2=2.765
r143 33 47 2.3025 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=3.345 $Y=1.935
+ $X2=3.255 $Y2=1.81
r144 33 35 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.345 $Y=1.935
+ $X2=3.345 $Y2=2.765
r145 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.08
+ $X2=0.69 $Y2=1.165
r146 31 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.08
+ $X2=0.345 $Y2=1.08
r147 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.995
+ $X2=0.345 $Y2=1.08
r148 27 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.26 $Y=0.995
+ $X2=0.26 $Y2=0.825
r149 26 36 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=2.765
+ $X2=3.345 $Y2=2.765
r150 25 51 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=1.85
+ $X2=3.345 $Y2=1.85
r151 24 36 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=2.765
+ $X2=3.345 $Y2=2.765
r152 23 51 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=1.85
+ $X2=3.345 $Y2=1.85
r153 19 26 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.605 $Y=2.9
+ $X2=3.53 $Y2=2.765
r154 19 21 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=3.605 $Y=2.9
+ $X2=3.605 $Y2=4.585
r155 15 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.605 $Y=1.715
+ $X2=3.53 $Y2=1.85
r156 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.605 $Y=1.715
+ $X2=3.605 $Y2=1.075
r157 11 24 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=2.9
+ $X2=3.25 $Y2=2.765
r158 11 13 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=3.175 $Y=2.9
+ $X2=3.175 $Y2=4.585
r159 7 23 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=1.715
+ $X2=3.25 $Y2=1.85
r160 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.175 $Y=1.715
+ $X2=3.175 $Y2=1.075
r161 2 57 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=5.835
r162 2 55 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=4.815
r163 1 29 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%A_428_89# 1 2 7 9 11 12 13 16 18 22 24
+ 27 30 33 35 36 37 40 44 47 50 55 56 59 63 66
c188 33 0 1.98654e-19 $X=2.335 $Y=1.76
c189 16 0 1.12321e-19 $X=2.815 $Y=4.585
r190 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=3.185
+ $X2=5.845 $Y2=3.185
r191 57 59 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=2.25
+ $X2=5.845 $Y2=2.25
r192 55 63 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=3.1
+ $X2=5.845 $Y2=3.185
r193 54 59 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.335
+ $X2=5.845 $Y2=2.25
r194 54 55 47.1364 $w=1.78e-07 $l=7.65e-07 $layer=LI1_cond $X=5.845 $Y=2.335
+ $X2=5.845 $Y2=3.1
r195 50 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.57 $Y=3.455
+ $X2=5.57 $Y2=5.835
r196 48 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=3.27
+ $X2=5.57 $Y2=3.185
r197 48 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.57 $Y=3.27
+ $X2=5.57 $Y2=3.455
r198 47 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=2.165
+ $X2=5.57 $Y2=2.25
r199 46 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.935
+ $X2=5.57 $Y2=1.85
r200 46 47 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.57 $Y=1.935
+ $X2=5.57 $Y2=2.165
r201 42 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.765
+ $X2=5.57 $Y2=1.85
r202 42 44 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.57 $Y=1.765
+ $X2=5.57 $Y2=0.825
r203 40 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.85
+ $X2=4.505 $Y2=2.015
r204 40 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.85
+ $X2=4.505 $Y2=1.685
r205 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=1.85 $X2=4.505 $Y2=1.85
r206 37 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=1.85
+ $X2=5.57 $Y2=1.85
r207 37 39 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.485 $Y=1.85
+ $X2=4.505 $Y2=1.85
r208 31 33 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.215 $Y=1.76
+ $X2=2.335 $Y2=1.76
r209 30 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.565 $Y=1.075
+ $X2=4.565 $Y2=1.685
r210 27 67 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.445 $Y=2.225
+ $X2=4.445 $Y2=2.015
r211 25 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=2.3
+ $X2=3.965 $Y2=2.3
r212 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.37 $Y=2.3
+ $X2=4.445 $Y2=2.225
r213 24 25 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.37 $Y=2.3
+ $X2=4.04 $Y2=2.3
r214 20 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.965 $Y=2.375
+ $X2=3.965 $Y2=2.3
r215 20 22 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=3.965 $Y=2.375
+ $X2=3.965 $Y2=4.585
r216 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.89 $Y=2.3
+ $X2=2.815 $Y2=2.3
r217 18 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.89 $Y=2.3
+ $X2=3.965 $Y2=2.3
r218 18 19 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.89 $Y=2.3 $X2=2.89
+ $Y2=2.3
r219 14 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.815 $Y=2.375
+ $X2=2.815 $Y2=2.3
r220 14 16 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=2.815 $Y=2.375
+ $X2=2.815 $Y2=4.585
r221 12 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.74 $Y=2.3
+ $X2=2.815 $Y2=2.3
r222 12 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.74 $Y=2.3
+ $X2=2.41 $Y2=2.3
r223 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.335 $Y=2.225
+ $X2=2.41 $Y2=2.3
r224 10 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.335 $Y=1.835
+ $X2=2.335 $Y2=1.76
r225 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.335 $Y=1.835
+ $X2=2.335 $Y2=2.225
r226 7 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.215 $Y=1.685
+ $X2=2.215 $Y2=1.76
r227 7 9 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.215 $Y=1.685
+ $X2=2.215 $Y2=1.075
r228 2 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5.43
+ $Y=3.085 $X2=5.57 $Y2=5.835
r229 2 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5.43
+ $Y=3.085 $X2=5.57 $Y2=3.455
r230 1 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.43
+ $Y=0.575 $X2=5.57 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%A_970_89# 1 2 9 13 21 25 28 29 30 33 35
+ 36 38 41 46 47 48 51 54 55 59 64 65
c166 64 0 2.20654e-19 $X=7.57 $Y=2.19
c167 29 0 8.77106e-20 $X=7.66 $Y=2.855
r168 64 66 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=2.19
+ $X2=7.572 $Y2=2.355
r169 64 65 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=2.19
+ $X2=7.572 $Y2=2.025
r170 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=2.19
+ $X2=4.985 $Y2=2.355
r171 59 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=2.19
+ $X2=4.985 $Y2=2.025
r172 55 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=2.19 $X2=7.57 $Y2=2.19
r173 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.57 $Y=2.19
+ $X2=7.57 $Y2=2.19
r174 51 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=2.19 $X2=4.985 $Y2=2.19
r175 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.985 $Y=2.19
+ $X2=4.985 $Y2=2.19
r176 48 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.13 $Y=2.19
+ $X2=4.985 $Y2=2.19
r177 47 54 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.425 $Y=2.19
+ $X2=7.57 $Y2=2.19
r178 47 48 2.20982 $w=1.7e-07 $l=2.295e-06 $layer=MET1_cond $X=7.425 $Y=2.19
+ $X2=5.13 $Y2=2.19
r179 45 55 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=6.605 $Y=2.19
+ $X2=7.57 $Y2=2.19
r180 45 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=2.19
+ $X2=6.52 $Y2=2.19
r181 41 43 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.52 $Y=4.815
+ $X2=6.52 $Y2=5.835
r182 39 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.275
+ $X2=6.52 $Y2=2.19
r183 39 41 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=6.52 $Y=2.275
+ $X2=6.52 $Y2=4.815
r184 38 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.105
+ $X2=6.52 $Y2=2.19
r185 37 38 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.52 $Y=1.165
+ $X2=6.52 $Y2=2.105
r186 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.435 $Y=1.08
+ $X2=6.52 $Y2=1.165
r187 35 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.435 $Y=1.08
+ $X2=6.175 $Y2=1.08
r188 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.09 $Y=0.995
+ $X2=6.175 $Y2=1.08
r189 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.09 $Y=0.995
+ $X2=6.09 $Y2=0.825
r190 29 30 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=2.855
+ $X2=7.66 $Y2=3.005
r191 29 66 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.635 $Y=2.855
+ $X2=7.635 $Y2=2.355
r192 28 65 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.635 $Y=1.8
+ $X2=7.635 $Y2=2.025
r193 27 28 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=1.65 $X2=7.66
+ $Y2=1.8
r194 25 30 1066.55 $w=1.5e-07 $l=2.08e-06 $layer=POLY_cond $X=7.685 $Y=5.085
+ $X2=7.685 $Y2=3.005
r195 21 27 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=7.685 $Y=0.945
+ $X2=7.685 $Y2=1.65
r196 13 61 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=4.925 $Y=4.585
+ $X2=4.925 $Y2=2.355
r197 9 60 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.925 $Y=1.075
+ $X2=4.925 $Y2=2.025
r198 2 43 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=4.085 $X2=6.52 $Y2=5.835
r199 2 41 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=4.085 $X2=6.52 $Y2=4.815
r200 1 33 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=5.965
+ $Y=0.575 $X2=6.09 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%A_808_115# 1 2 9 13 15 16 17 18 21 25 31
+ 32 35 38 39 45
c128 35 0 1.57671e-19 $X=3.685 $Y=1.85
c129 32 0 1.5821e-19 $X=3.83 $Y=1.85
c130 15 0 1.67294e-19 $X=4.095 $Y=1.43
r131 43 45 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.1 $Y=1.85
+ $X2=6.305 $Y2=1.85
r132 39 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.1
+ $Y=1.85 $X2=6.1 $Y2=1.85
r133 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.1 $Y=1.85 $X2=6.1
+ $Y2=1.85
r134 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=1.85
+ $X2=3.685 $Y2=1.85
r135 32 34 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.83 $Y=1.85
+ $X2=3.685 $Y2=1.85
r136 31 38 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.955 $Y=1.85
+ $X2=6.1 $Y2=1.85
r137 31 32 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=5.955 $Y=1.85
+ $X2=3.83 $Y2=1.85
r138 30 35 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.685 $Y=3.1
+ $X2=3.685 $Y2=1.85
r139 29 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.685 $Y=1.515
+ $X2=3.685 $Y2=1.85
r140 25 27 69.1466 $w=3.38e-07 $l=2.04e-06 $layer=LI1_cond $X=4.265 $Y=3.795
+ $X2=4.265 $Y2=5.835
r141 23 25 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=4.265 $Y=3.27
+ $X2=4.265 $Y2=3.795
r142 19 21 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=4.265 $Y=1.345
+ $X2=4.265 $Y2=0.825
r143 18 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.77 $Y=3.185
+ $X2=3.685 $Y2=3.1
r144 17 23 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=3.185
+ $X2=4.265 $Y2=3.27
r145 17 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=3.185
+ $X2=3.77 $Y2=3.185
r146 16 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.77 $Y=1.43
+ $X2=3.685 $Y2=1.515
r147 15 19 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=1.43
+ $X2=4.265 $Y2=1.345
r148 15 16 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=1.43
+ $X2=3.77 $Y2=1.43
r149 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=2.015
+ $X2=6.305 $Y2=1.85
r150 11 13 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=6.305 $Y=2.015
+ $X2=6.305 $Y2=5.085
r151 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.685
+ $X2=6.305 $Y2=1.85
r152 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.305 $Y=1.685
+ $X2=6.305 $Y2=0.945
r153 2 27 171.429 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=3 $X=4.04
+ $Y=3.085 $X2=4.265 $Y2=5.835
r154 2 25 171.429 $w=1.7e-07 $l=8.1477e-07 $layer=licon1_PDIFF $count=3 $X=4.04
+ $Y=3.085 $X2=4.265 $Y2=3.795
r155 1 21 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=4.04
+ $Y=0.575 $X2=4.265 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%QN 1 2 9 13 17 19 20 21 22 26 27 31 32
c83 32 0 8.77106e-20 $X=7.475 $Y=2.96
c84 21 0 9.99996e-20 $X=7.97 $Y=2.765
c85 19 0 1.20654e-19 $X=7.97 $Y=1.85
r86 39 41 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.47 $Y=4.475
+ $X2=7.47 $Y2=5.835
r87 31 39 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=7.47 $Y=2.96
+ $X2=7.47 $Y2=4.475
r88 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.47 $Y=2.96
+ $X2=7.47 $Y2=2.96
r89 28 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.47 $Y=2.85
+ $X2=7.47 $Y2=2.96
r90 27 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.395
+ $X2=8.055 $Y2=2.56
r91 27 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.395
+ $X2=8.055 $Y2=2.23
r92 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=2.395 $X2=8.055 $Y2=2.395
r93 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.055 $Y=2.68
+ $X2=8.055 $Y2=2.395
r94 23 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.055 $Y=1.935
+ $X2=8.055 $Y2=2.395
r95 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=2.765
+ $X2=7.47 $Y2=2.85
r96 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=2.765
+ $X2=8.055 $Y2=2.68
r97 21 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=2.765
+ $X2=7.555 $Y2=2.765
r98 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=1.85
+ $X2=8.055 $Y2=1.935
r99 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=1.85
+ $X2=7.555 $Y2=1.85
r100 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=1.765
+ $X2=7.555 $Y2=1.85
r101 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=7.47 $Y=1.765
+ $X2=7.47 $Y2=0.825
r102 13 36 1294.73 $w=1.5e-07 $l=2.525e-06 $layer=POLY_cond $X=8.115 $Y=5.085
+ $X2=8.115 $Y2=2.56
r103 9 35 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=8.115 $Y=0.945
+ $X2=8.115 $Y2=2.23
r104 2 41 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=4.085 $X2=7.47 $Y2=5.835
r105 2 39 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=4.085 $X2=7.47 $Y2=4.475
r106 1 17 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFS_L%Q 1 2 9 13 18 21 24 26
r22 26 29 6.68493 $w=2.19e-07 $l=1.2e-07 $layer=LI1_cond $X=8.325 $Y=3.287
+ $X2=8.445 $Y2=3.287
r23 24 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.325 $Y=3.33
+ $X2=8.325 $Y2=3.33
r24 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=1.515
+ $X2=8.445 $Y2=1.515
r25 18 29 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.445 $Y=3.16
+ $X2=8.445 $Y2=3.287
r26 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=1.6
+ $X2=8.445 $Y2=1.515
r27 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=8.445 $Y=1.6
+ $X2=8.445 $Y2=3.16
r28 13 15 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=8.33 $Y=4.475
+ $X2=8.33 $Y2=5.835
r29 11 26 2.22295 $w=1.7e-07 $l=1.30476e-07 $layer=LI1_cond $X=8.33 $Y=3.415
+ $X2=8.325 $Y2=3.287
r30 11 13 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=8.33 $Y=3.415
+ $X2=8.33 $Y2=4.475
r31 7 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=1.43 $X2=8.33
+ $Y2=1.515
r32 7 9 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.33 $Y=1.43 $X2=8.33
+ $Y2=0.825
r33 2 15 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=4.085 $X2=8.33 $Y2=5.835
r34 2 13 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=4.085 $X2=8.33 $Y2=4.475
r35 1 9 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.575 $X2=8.33 $Y2=0.825
.ends

