* File: sky130_osu_sc_12T_ls__tnbufi_1.pex.spice
* Created: Fri Nov 12 15:40:49 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_1%GND 1 17 19 26 35 38
r34 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r35 28 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r36 24 33 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r37 24 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r38 19 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r39 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r40 17 28 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=0.775
+ $Y2=0.152
r41 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r42 1 26 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_1%VDD 1 13 15 21 25 29 32
r19 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r20 25 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r21 23 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r22 23 25 9.8 $w=3.05e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287 $X2=1.02
+ $Y2=4.287
r23 19 27 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r24 19 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=3.295
r25 15 27 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r26 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r27 13 25 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r28 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r29 1 21 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_1%A_27_115# 1 3 11 16 20 24 28 30 33
r44 29 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.695
+ $X2=0.26 $Y2=1.695
r45 28 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=1.695
+ $X2=0.69 $Y2=1.695
r46 28 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.695
+ $X2=0.345 $Y2=1.695
r47 24 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r48 22 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.78 $X2=0.26
+ $Y2=1.695
r49 22 24 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=0.26 $Y=1.78
+ $X2=0.26 $Y2=2.955
r50 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.61 $X2=0.26
+ $Y2=1.695
r51 18 20 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.26 $Y=1.61
+ $X2=0.26 $Y2=0.755
r52 14 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.695 $X2=0.69 $Y2=1.695
r53 14 16 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=1.695
+ $X2=0.905 $Y2=1.695
r54 9 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.53
+ $X2=0.905 $Y2=1.695
r55 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.905 $Y=1.53
+ $X2=0.905 $Y2=0.835
r56 3 26 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r57 3 24 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r58 1 20 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_1%OE 3 5 6 8 11 14 19 25
r42 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r43 19 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.69 $Y=2.285
+ $X2=0.69 $Y2=2.48
r44 17 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=2.285 $X2=0.69 $Y2=2.285
r45 12 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.245
+ $X2=0.475 $Y2=1.245
r46 6 17 49.2914 $w=4.58e-07 $l=4.23124e-07 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.587 $Y2=2.285
r47 6 11 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=3.235
r48 6 8 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=2.53
+ $X2=0.475 $Y2=3.235
r49 3 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.17
+ $X2=0.475 $Y2=1.245
r50 3 5 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=1.17
+ $X2=0.475 $Y2=0.835
r51 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=1.32 $X2=0.27
+ $Y2=1.245
r52 1 6 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.27 $Y=1.32 $X2=0.27
+ $Y2=2.38
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_1%A 3 7 10 15 20 23
r47 17 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.61
+ $X2=1.325 $Y2=1.61
r48 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=2.85
+ $X2=1.14 $Y2=2.85
r49 13 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.695
+ $X2=1.14 $Y2=1.61
r50 13 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.14 $Y=1.695
+ $X2=1.14 $Y2=2.85
r51 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.61 $X2=1.325 $Y2=1.61
r52 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.61
+ $X2=1.325 $Y2=1.775
r53 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.61
+ $X2=1.325 $Y2=1.445
r54 7 12 748.638 $w=1.5e-07 $l=1.46e-06 $layer=POLY_cond $X=1.265 $Y=3.235
+ $X2=1.265 $Y2=1.775
r55 3 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.265 $Y=0.835
+ $X2=1.265 $Y2=1.445
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__TNBUFI_1%Y 1 3 10 16 26 29 32
r32 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.995
+ $X2=1.48 $Y2=2.11
r33 24 26 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.48 $Y=1.995
+ $X2=1.48 $Y2=1.34
r34 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.48 $Y=1.115
+ $X2=1.48 $Y2=1
r35 23 26 0.216649 $w=1.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.48 $Y=1.115
+ $X2=1.48 $Y2=1.34
r36 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.48 $Y=2.955
+ $X2=1.48 $Y2=3.635
r37 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=2.11
+ $X2=1.48 $Y2=2.11
r38 16 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.48 $Y=2.11
+ $X2=1.48 $Y2=2.955
r39 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.48 $Y=1 $X2=1.48
+ $Y2=1
r40 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.48 $Y=0.755
+ $X2=1.48 $Y2=1
r41 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.48 $Y2=3.635
r42 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.48 $Y2=2.955
r43 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.34 $Y=0.575
+ $X2=1.48 $Y2=0.755
.ends

