* File: sky130_osu_sc_18T_hs__buf_4.pex.spice
* Created: Fri Nov 12 13:48:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__BUF_4%GND 1 2 3 31 35 39 41 42 49 63 65
r57 63 65 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r58 47 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.825
r59 41 47 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.325 $Y=0.152
+ $X2=2.41 $Y2=0.305
r60 37 42 3.38889 $w=3.06e-07 $l=8.6487e-08 $layer=LI1_cond $X=1.55 $Y=0.155
+ $X2=1.635 $Y2=0.152
r61 37 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.825
r62 33 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r63 31 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r64 31 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r65 31 37 21.1307 $w=3.06e-07 $l=5.3e-07 $layer=LI1_cond $X=1.02 $Y=0.155
+ $X2=1.55 $Y2=0.155
r66 31 33 13.1569 $w=3.06e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=0.155
+ $X2=0.69 $Y2=0.155
r67 31 33 13.9542 $w=3.06e-07 $l=3.5e-07 $layer=LI1_cond $X=0.34 $Y=0.155
+ $X2=0.69 $Y2=0.155
r68 31 41 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r69 31 42 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r70 3 49 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r71 2 39 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r72 1 35 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_4%VDD 1 2 3 25 27 34 38 44 48 55 62 66
r44 62 66 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r45 55 58 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r46 53 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=5.835
r47 51 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.47 $X2=1.7
+ $Y2=6.47
r48 49 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.55 $Y2=6.507
r49 49 51 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.7 $Y2=6.507
r50 48 53 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=2.41 $Y2=6.355
r51 48 51 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=1.7 $Y2=6.507
r52 44 47 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r53 42 60 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=6.507
r54 42 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=5.835
r55 39 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r56 39 41 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r57 38 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.55 $Y2=6.507
r58 38 41 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.02 $Y2=6.507
r59 34 37 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r60 32 59 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r61 32 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r62 29 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r63 27 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r64 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r65 25 51 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r66 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r67 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r68 3 58 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r69 3 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r70 2 47 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r71 2 44 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r72 1 37 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r73 1 34 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_4%A 3 7 10 14 20
r39 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=3.33
r40 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2.48
+ $X2=0.635 $Y2=3.33
r41 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.48 $X2=0.635 $Y2=2.48
r42 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.645
r43 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.315
r44 7 12 994.766 $w=1.5e-07 $l=1.94e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.645
r45 3 11 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.315
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_4%A_27_115# 1 3 11 13 15 17 20 22 24 25 26
+ 27 28 31 33 35 36 38 42 44 46 56 57 60 64 68 70 73
c118 33 0 1.33323e-19 $X=1.765 $Y=3.01
c119 31 0 1.33323e-19 $X=1.765 $Y=1.075
c120 22 0 1.33323e-19 $X=1.335 $Y=3.01
c121 20 0 1.33323e-19 $X=1.335 $Y=1.075
r122 69 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.935
+ $X2=0.26 $Y2=1.935
r123 68 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.965 $Y2=1.935
r124 68 69 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.345 $Y2=1.935
r125 64 66 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r126 62 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=1.935
r127 62 64 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=3.455
r128 58 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=1.935
r129 58 60 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r130 53 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.935 $X2=0.965 $Y2=1.935
r131 53 54 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=1.18 $Y2=1.935
r132 51 53 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.935
+ $X2=0.965 $Y2=1.935
r133 49 50 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.935
+ $X2=1.335 $Y2=2.935
r134 47 49 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.935
+ $X2=1.18 $Y2=2.935
r135 44 46 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=4.585
r136 40 42 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r137 39 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.935
+ $X2=1.765 $Y2=2.935
r138 38 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=2.195 $Y2=3.01
r139 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=1.84 $Y2=2.935
r140 37 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.765 $Y2=1.845
r141 36 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.77
r142 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r143 33 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=2.935
r144 33 35 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=4.585
r145 29 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.845
r146 29 31 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r147 28 50 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.935
+ $X2=1.335 $Y2=2.935
r148 27 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.765 $Y2=2.935
r149 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.41 $Y2=2.935
r150 25 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.765 $Y2=1.845
r151 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.41 $Y2=1.845
r152 22 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=2.935
r153 22 24 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=4.585
r154 18 26 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.41 $Y2=1.845
r155 18 54 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.18 $Y2=1.935
r156 18 20 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r157 17 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.86
+ $X2=1.18 $Y2=2.935
r158 16 54 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=1.935
r159 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=2.86
r160 13 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=2.935
r161 13 15 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=4.585
r162 9 51 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.935
r163 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.075
r164 3 66 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r165 3 64 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r166 1 60 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__BUF_4%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c80 55 0 1.33323e-19 $X=1.98 $Y=2.845
c81 54 0 1.33323e-19 $X=1.98 $Y=1.595
c82 46 0 1.33323e-19 $X=1.12 $Y=2.845
c83 45 0 1.33323e-19 $X=1.12 $Y=1.595
r84 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.845
+ $X2=1.98 $Y2=2.96
r85 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=1.48
r86 54 55 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=2.845
r87 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.96
+ $X2=1.12 $Y2=2.96
r88 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.98 $Y2=2.96
r89 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.265 $Y2=2.96
r90 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1.48
+ $X2=1.12 $Y2=1.48
r91 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.98 $Y2=1.48
r92 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.265 $Y2=1.48
r93 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.96
r94 46 48 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.27
r95 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=1.48
r96 45 48 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=2.27
r97 41 43 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r98 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=2.96
r99 38 41 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=3.455
r100 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=1.48
r101 32 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.98 $Y=0.825
+ $X2=1.98 $Y2=1.48
r102 27 29 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r103 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=2.96
r104 24 27 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=3.455
r105 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=1.48
r106 18 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.12 $Y=0.825
+ $X2=1.12 $Y2=1.48
r107 6 43 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r108 6 41 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r109 5 29 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r110 5 27 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r111 2 32 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r112 1 18 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
.ends

