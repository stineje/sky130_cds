* File: sky130_osu_sc_15T_hs__and2_8.pex.spice
* Created: Fri Nov 12 14:27:15 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__AND2_8%GND 1 2 3 4 5 63 65 73 75 82 84 91 93
+ 100 102 110 123 125
r141 123 125 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=4.42 $Y2=0.152
r142 108 110 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.56 $Y=0.305
+ $X2=4.56 $Y2=0.9
r143 102 108 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.475
+ $Y=0.152 $X2=4.56 $Y2=0.305
r144 98 100 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.9
r145 94 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r146 89 116 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r147 89 91 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.9
r148 85 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r149 84 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r150 80 115 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r151 80 82 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.9
r152 75 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r153 71 73 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.9
r154 63 125 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r155 63 123 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r156 63 98 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.7 $Y2=0.305
r157 63 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.615 $Y2=0.152
r158 63 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.152
+ $X2=3.785 $Y2=0.152
r159 63 71 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r160 63 65 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r161 63 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r162 63 102 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.475 $Y2=0.152
r163 63 103 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=3.785 $Y2=0.152
r164 63 93 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r165 63 94 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r166 63 84 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r167 63 85 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r168 63 75 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r169 63 76 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r170 63 65 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r171 5 110 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.575 $X2=4.56 $Y2=0.9
r172 4 100 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.9
r173 3 91 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.9
r174 2 82 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.9
r175 1 73 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.9
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__AND2_8%VDD 1 2 3 4 5 6 53 57 61 67 71 77 81 87
+ 91 97 101 108 121 125
r87 121 125 1.90014 $w=3.05e-07 $l=4.08e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=4.42 $Y2=5.397
r88 113 121 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r89 108 111 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.56 $Y=3.215
+ $X2=4.56 $Y2=4.575
r90 106 111 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.56 $Y=5.245
+ $X2=4.56 $Y2=4.575
r91 104 125 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.42 $Y=5.36
+ $X2=4.42 $Y2=5.36
r92 102 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=5.397
+ $X2=3.7 $Y2=5.397
r93 102 104 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=5.397
+ $X2=4.42 $Y2=5.397
r94 101 106 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.475 $Y=5.397
+ $X2=4.56 $Y2=5.245
r95 101 104 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=4.475 $Y=5.397
+ $X2=4.42 $Y2=5.397
r96 97 100 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.7 $Y=3.215
+ $X2=3.7 $Y2=4.575
r97 95 119 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.7 $Y=5.245
+ $X2=3.7 $Y2=5.397
r98 95 100 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.7 $Y=5.245
+ $X2=3.7 $Y2=4.575
r99 92 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=2.84 $Y2=5.397
r100 92 94 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=3.06 $Y2=5.397
r101 91 119 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.7 $Y2=5.397
r102 91 94 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.06 $Y2=5.397
r103 87 90 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.215
+ $X2=2.84 $Y2=4.575
r104 85 117 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=5.397
r105 85 90 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.575
r106 82 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r107 82 84 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r108 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.397
r109 81 84 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r110 77 80 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.215
+ $X2=1.98 $Y2=4.575
r111 75 116 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r112 75 80 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.575
r113 72 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r114 72 74 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r115 71 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r116 71 74 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r117 67 70 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=3.555
+ $X2=1.12 $Y2=4.575
r118 65 115 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r119 65 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.575
r120 62 113 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r121 62 64 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r122 61 115 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r123 61 64 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r124 57 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.895
+ $X2=0.26 $Y2=4.575
r125 55 113 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r126 55 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.575
r127 53 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=5.245 $X2=4.42 $Y2=5.33
r128 53 119 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r129 53 94 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r130 53 84 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r131 53 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r132 53 64 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r133 53 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r134 6 111 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.825 $X2=4.56 $Y2=4.575
r135 6 108 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.825 $X2=4.56 $Y2=3.215
r136 5 100 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=4.575
r137 5 97 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=3.215
r138 4 90 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.575
r139 4 87 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.215
r140 3 80 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.575
r141 3 77 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.215
r142 2 70 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r143 2 67 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.555
r144 1 60 400 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r145 1 57 400 $w=1.7e-07 $l=1.13077e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__AND2_8%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=3.07
+ $X2=0.275 $Y2=3.07
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.07
+ $X2=0.27 $Y2=3.07
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.505
+ $X2=0.27 $Y2=3.07
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.505 $X2=0.27 $Y2=2.505
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.505
+ $X2=0.475 $Y2=2.505
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=2.505
r38 5 7 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=3.825
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=2.505
r40 1 3 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=0.895
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__AND2_8%B 3 7 10 14 22
c41 7 0 1.37149e-19 $X=0.905 $Y=3.825
r42 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.7
+ $X2=0.955 $Y2=2.7
r43 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.7 $X2=0.95
+ $Y2=2.7
r44 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.165
+ $X2=0.95 $Y2=2.7
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.165 $X2=0.95 $Y2=2.165
r46 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2.33
r47 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2
r48 7 12 766.585 $w=1.5e-07 $l=1.495e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.33
r49 3 11 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=0.835 $Y=0.895
+ $X2=0.835 $Y2=2
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__AND2_8%A_27_115# 1 3 11 13 15 17 18 22 24 26 27
+ 28 29 33 35 37 38 40 44 46 48 49 51 55 58 59 61 62 64 68 70 72 73 75 79 81 83
+ 84 86 90 92 94 95 101 102 103 104 105 106 107 108 109 110 111 114 116 117 122
+ 128 130 131 132
c243 79 0 1.77221e-19 $X=3.915 $Y=0.895
c244 68 0 1.33323e-19 $X=3.485 $Y=0.895
c245 55 0 1.33323e-19 $X=3.055 $Y=0.895
c246 44 0 1.33323e-19 $X=2.625 $Y=0.895
c247 33 0 1.33323e-19 $X=2.195 $Y=0.895
c248 22 0 1.33323e-19 $X=1.765 $Y=0.895
r249 131 132 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.305
+ $X2=0.65 $Y2=3.475
r250 126 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=0.61 $Y2=1.675
r251 126 128 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=1.43 $Y2=1.675
r252 122 124 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=3.555
+ $X2=0.69 $Y2=4.575
r253 122 132 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.555
+ $X2=0.69 $Y2=3.475
r254 118 130 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=1.675
r255 118 131 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=3.305
r256 116 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.61 $Y2=1.675
r257 116 117 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.345 $Y2=1.675
r258 112 117 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.345 $Y2=1.675
r259 112 114 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.9
r260 99 128 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.675 $X2=1.43 $Y2=1.675
r261 97 99 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.675
+ $X2=1.43 $Y2=1.675
r262 96 97 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.37 $Y2=1.675
r263 92 94 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=4.345 $Y=2.7
+ $X2=4.345 $Y2=3.825
r264 88 90 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.345 $Y=1.51
+ $X2=4.345 $Y2=0.895
r265 87 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=2.625
+ $X2=3.915 $Y2=2.625
r266 86 92 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=2.625
+ $X2=4.345 $Y2=2.7
r267 86 87 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=2.625
+ $X2=3.99 $Y2=2.625
r268 85 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.585
+ $X2=3.915 $Y2=1.585
r269 84 88 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.27 $Y=1.585
+ $X2=4.345 $Y2=1.51
r270 84 85 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.585
+ $X2=3.99 $Y2=1.585
r271 81 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=2.7
+ $X2=3.915 $Y2=2.625
r272 81 83 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.915 $Y=2.7
+ $X2=3.915 $Y2=3.825
r273 77 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=1.51
+ $X2=3.915 $Y2=1.585
r274 77 79 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.915 $Y=1.51
+ $X2=3.915 $Y2=0.895
r275 76 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.625
+ $X2=3.485 $Y2=2.625
r276 75 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.625
+ $X2=3.915 $Y2=2.625
r277 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.625
+ $X2=3.56 $Y2=2.625
r278 74 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.585
+ $X2=3.485 $Y2=1.585
r279 73 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.585
+ $X2=3.915 $Y2=1.585
r280 73 74 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.585
+ $X2=3.56 $Y2=1.585
r281 70 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=2.625
r282 70 72 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=3.825
r283 66 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.51
+ $X2=3.485 $Y2=1.585
r284 66 68 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.485 $Y=1.51
+ $X2=3.485 $Y2=0.895
r285 65 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.625
+ $X2=3.055 $Y2=2.625
r286 64 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.485 $Y2=2.625
r287 64 65 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.13 $Y2=2.625
r288 63 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.585
+ $X2=3.055 $Y2=1.585
r289 62 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.585
+ $X2=3.485 $Y2=1.585
r290 62 63 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.585
+ $X2=3.13 $Y2=1.585
r291 59 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=2.625
r292 59 61 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=3.825
r293 58 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.55
+ $X2=3.055 $Y2=2.625
r294 57 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.66
+ $X2=3.055 $Y2=1.585
r295 57 58 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.055 $Y=1.66
+ $X2=3.055 $Y2=2.55
r296 53 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.51
+ $X2=3.055 $Y2=1.585
r297 53 55 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.055 $Y=1.51
+ $X2=3.055 $Y2=0.895
r298 52 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.625
+ $X2=2.625 $Y2=2.625
r299 51 107 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=3.055 $Y2=2.625
r300 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=2.7 $Y2=2.625
r301 50 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.585
+ $X2=2.625 $Y2=1.585
r302 49 106 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.585
+ $X2=3.055 $Y2=1.585
r303 49 50 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.585
+ $X2=2.7 $Y2=1.585
r304 46 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=2.625
r305 46 48 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r306 42 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.625 $Y2=1.585
r307 42 44 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.625 $Y2=0.895
r308 41 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r309 40 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.625
r310 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r311 39 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.585
+ $X2=2.195 $Y2=1.585
r312 38 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.625 $Y2=1.585
r313 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.27 $Y2=1.585
r314 35 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=2.625
r315 35 37 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r316 31 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=1.585
r317 31 33 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=0.895
r318 30 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r319 29 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r320 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r321 27 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=2.195 $Y2=1.585
r322 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=1.84 $Y2=1.585
r323 24 101 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r324 24 26 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r325 20 28 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.84 $Y2=1.585
r326 20 99 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.43 $Y2=1.675
r327 20 22 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=0.895
r328 19 95 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.625
+ $X2=1.352 $Y2=2.625
r329 18 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r330 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.445 $Y2=2.625
r331 17 95 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.55
+ $X2=1.352 $Y2=2.625
r332 16 97 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=1.675
r333 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=2.55
r334 13 95 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.352 $Y2=2.625
r335 13 15 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r336 9 96 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=1.675
r337 9 11 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.895
r338 3 124 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.575
r339 3 122 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.555
r340 1 114 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.9
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__AND2_8%Y 1 2 3 4 9 10 11 12 34 40 48 54 62 68
+ 76 82 89 90 92 94 96 99 100 101 102 103 104 105 106 107 110 111 125
c164 110 0 1.33323e-19 $X=4.13 $Y=1.335
c165 104 0 3.10545e-19 $X=3.27 $Y=1.335
c166 101 0 2.66647e-19 $X=2.555 $Y=1.22
c167 89 0 1.33323e-19 $X=1.55 $Y=1.335
c168 40 0 1.37149e-19 $X=1.55 $Y=2.33
r169 111 127 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=2.215
+ $X2=4.13 $Y2=2.33
r170 110 125 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=4.13 $Y=1.335
+ $X2=4.13 $Y2=1.22
r171 110 111 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=4.13 $Y=1.335
+ $X2=4.13 $Y2=2.215
r172 107 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.415 $Y=2.33
+ $X2=3.27 $Y2=2.33
r173 106 127 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.985 $Y=2.33
+ $X2=4.13 $Y2=2.33
r174 106 107 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.985 $Y=2.33
+ $X2=3.415 $Y2=2.33
r175 105 123 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.215
+ $X2=3.27 $Y2=2.33
r176 104 121 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=1.22
r177 104 105 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=2.215
r178 103 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.33
+ $X2=2.41 $Y2=2.33
r179 102 123 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.33
+ $X2=3.27 $Y2=2.33
r180 102 103 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.33
+ $X2=2.555 $Y2=2.33
r181 101 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.22
+ $X2=2.41 $Y2=1.22
r182 100 121 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=3.27 $Y2=1.22
r183 100 101 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=2.555 $Y2=1.22
r184 99 119 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.215
+ $X2=2.41 $Y2=2.33
r185 98 117 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r186 98 99 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.215
r187 97 115 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.33
+ $X2=1.55 $Y2=2.33
r188 96 119 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=2.41 $Y2=2.33
r189 96 97 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=1.695 $Y2=2.33
r190 95 113 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r191 94 117 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r192 94 95 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r193 90 115 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r194 90 92 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r195 89 113 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r196 89 92 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r197 85 87 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.13 $Y=3.215
+ $X2=4.13 $Y2=4.575
r198 82 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=2.33
+ $X2=4.13 $Y2=2.33
r199 82 85 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.13 $Y=2.33
+ $X2=4.13 $Y2=3.215
r200 79 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.13 $Y=1.22
+ $X2=4.13 $Y2=1.22
r201 76 79 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.13 $Y=0.9 $X2=4.13
+ $Y2=1.22
r202 71 73 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.27 $Y=3.215
+ $X2=3.27 $Y2=4.575
r203 68 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.33
+ $X2=3.27 $Y2=2.33
r204 68 71 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.27 $Y=2.33
+ $X2=3.27 $Y2=3.215
r205 65 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.22
+ $X2=3.27 $Y2=1.22
r206 62 65 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.27 $Y=0.9 $X2=3.27
+ $Y2=1.22
r207 57 59 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.215
+ $X2=2.41 $Y2=4.575
r208 54 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=2.33
r209 54 57 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=3.215
r210 51 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r211 48 51 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.41 $Y=0.9 $X2=2.41
+ $Y2=1.22
r212 43 45 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.215
+ $X2=1.55 $Y2=4.575
r213 40 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r214 40 43 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=3.215
r215 37 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r216 34 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.55 $Y=0.9 $X2=1.55
+ $Y2=1.22
r217 12 87 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.825 $X2=4.13 $Y2=4.575
r218 12 85 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.825 $X2=4.13 $Y2=3.215
r219 11 73 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=4.575
r220 11 71 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=3.215
r221 10 59 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.575
r222 10 57 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.215
r223 9 45 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.575
r224 9 43 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.215
r225 4 76 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.9
r226 3 62 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.9
r227 2 48 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.9
r228 1 34 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.9
.ends

