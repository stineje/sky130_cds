* File: sky130_osu_sc_12T_hs__addf_1.pxi.spice
* Created: Fri Nov 12 15:06:11 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%GND N_GND_M1013_d N_GND_M1027_d N_GND_M1024_d
+ N_GND_M1004_d N_GND_M1023_s N_GND_M1013_b N_GND_c_2_p N_GND_c_3_p N_GND_c_7_p
+ N_GND_c_8_p N_GND_c_19_p N_GND_c_54_p N_GND_c_28_p N_GND_c_26_p N_GND_c_131_p
+ N_GND_c_108_p N_GND_c_55_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_HS__ADDF_1%GND
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%VDD N_VDD_M1000_d N_VDD_M1016_d N_VDD_M1011_d
+ N_VDD_M1021_d N_VDD_M1010_s N_VDD_M1000_b N_VDD_c_177_p N_VDD_c_178_p
+ N_VDD_c_181_p N_VDD_c_182_p N_VDD_c_189_p N_VDD_c_208_p N_VDD_c_192_p
+ N_VDD_c_193_p N_VDD_c_257_p N_VDD_c_243_p N_VDD_c_244_p VDD N_VDD_c_179_p
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%VDD
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%A N_A_M1013_g N_A_M1000_g N_A_c_305_n
+ N_A_M1027_g N_A_c_347_n N_A_M1016_g N_A_c_309_n N_A_c_311_n N_A_c_312_n
+ N_A_c_313_n N_A_c_314_n N_A_c_315_n N_A_c_316_n N_A_M1022_g N_A_c_354_n
+ N_A_M1009_g N_A_M1004_g N_A_M1021_g N_A_c_320_n N_A_c_321_n N_A_c_322_n
+ N_A_c_323_n N_A_c_324_n N_A_c_326_n N_A_c_330_n N_A_c_331_n N_A_c_332_n
+ N_A_c_333_n N_A_c_335_n N_A_c_336_n N_A_c_338_n N_A_c_339_n N_A_c_340_n
+ N_A_c_341_n A N_A_c_342_n PM_SKY130_OSU_SC_12T_HS__ADDF_1%A
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%B N_B_M1001_g N_B_M1019_g N_B_M1025_g
+ N_B_M1012_g N_B_M1024_g N_B_M1011_g N_B_M1017_g N_B_M1006_g N_B_c_551_n
+ N_B_c_552_n N_B_c_553_n N_B_c_554_n N_B_c_555_n N_B_c_556_n N_B_c_584_n
+ N_B_c_585_n N_B_c_557_n N_B_c_558_n N_B_c_559_n N_B_c_560_n N_B_c_561_n
+ N_B_c_562_n B N_B_c_563_n N_B_c_593_n N_B_c_564_n N_B_c_565_n N_B_c_566_n
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%B
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%CI N_CI_M1003_g N_CI_M1020_g N_CI_M1014_g
+ N_CI_M1002_g N_CI_M1008_g N_CI_M1026_g N_CI_c_819_n N_CI_c_820_n N_CI_c_821_n
+ N_CI_c_822_n N_CI_c_823_n N_CI_c_824_n N_CI_c_825_n N_CI_c_826_n N_CI_c_827_n
+ N_CI_c_828_n CI N_CI_c_829_n PM_SKY130_OSU_SC_12T_HS__ADDF_1%CI
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%CON N_CON_M1003_d N_CON_M1020_d N_CON_M1015_g
+ N_CON_M1005_g N_CON_M1023_g N_CON_M1010_g N_CON_c_992_n N_CON_c_993_n
+ N_CON_c_994_n N_CON_c_1020_n N_CON_c_997_n N_CON_c_998_n N_CON_c_999_n
+ N_CON_c_1026_n N_CON_c_1000_n N_CON_c_1001_n N_CON_c_1003_n N_CON_c_1005_n
+ N_CON_c_1006_n N_CON_c_1008_n CON PM_SKY130_OSU_SC_12T_HS__ADDF_1%CON
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_784_115# N_A_784_115#_M1015_d
+ N_A_784_115#_M1005_d N_A_784_115#_M1018_g N_A_784_115#_M1007_g
+ N_A_784_115#_c_1161_n N_A_784_115#_c_1162_n N_A_784_115#_c_1163_n
+ N_A_784_115#_c_1164_n N_A_784_115#_c_1177_n N_A_784_115#_c_1178_n
+ N_A_784_115#_c_1181_n N_A_784_115#_c_1165_n N_A_784_115#_c_1183_n
+ N_A_784_115#_c_1166_n N_A_784_115#_c_1169_n
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_784_115#
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_27_521# N_A_27_521#_M1000_s
+ N_A_27_521#_M1019_d N_A_27_521#_c_1285_n N_A_27_521#_c_1288_n
+ N_A_27_521#_c_1290_n PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_27_521#
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_526_521# N_A_526_521#_M1009_d
+ N_A_526_521#_M1002_d N_A_526_521#_c_1300_n N_A_526_521#_c_1302_n
+ N_A_526_521#_c_1305_n PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_526_521#
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%S N_S_M1018_d N_S_M1007_d N_S_c_1317_n
+ N_S_c_1323_n N_S_c_1321_n N_S_c_1322_n N_S_c_1328_n S
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%S
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%CO N_CO_M1023_d N_CO_M1010_d N_CO_c_1368_n CO
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%CO
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_27_115# N_A_27_115#_M1013_s
+ N_A_27_115#_M1001_d N_A_27_115#_c_1384_n N_A_27_115#_c_1387_n
+ N_A_27_115#_c_1390_n N_A_27_115#_c_1394_n
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_27_115#
x_PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_526_115# N_A_526_115#_M1022_d
+ N_A_526_115#_M1014_d N_A_526_115#_c_1410_n N_A_526_115#_c_1415_n
+ N_A_526_115#_c_1418_n N_A_526_115#_c_1419_n
+ PM_SKY130_OSU_SC_12T_HS__ADDF_1%A_526_115#
cc_1 N_GND_M1013_b N_A_M1013_g 0.0516715f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_A_M1013_g 0.00640094f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_A_M1013_g 0.00411218f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.85
cc_4 N_GND_c_4_p N_A_M1013_g 0.0048006f $X=6.46 $Y=0.19 $X2=0.475 $Y2=0.85
cc_5 N_GND_M1013_b N_A_M1000_g 0.0395507f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_6 N_GND_M1013_b N_A_c_305_n 0.0158117f $X=-0.045 $Y=0 $X2=2.125 $Y2=1.205
cc_7 N_GND_c_7_p N_A_c_305_n 0.0063578f $X=2.255 $Y=0.152 $X2=2.125 $Y2=1.205
cc_8 N_GND_c_8_p N_A_c_305_n 0.00387281f $X=2.34 $Y=0.755 $X2=2.125 $Y2=1.205
cc_9 N_GND_c_4_p N_A_c_305_n 0.00478641f $X=6.46 $Y=0.19 $X2=2.125 $Y2=1.205
cc_10 N_GND_M1013_b N_A_c_309_n 0.00951622f $X=-0.045 $Y=0 $X2=2.36 $Y2=1.28
cc_11 N_GND_c_8_p N_A_c_309_n 0.00304403f $X=2.34 $Y=0.755 $X2=2.36 $Y2=1.28
cc_12 N_GND_M1013_b N_A_c_311_n 0.00808138f $X=-0.045 $Y=0 $X2=2.2 $Y2=1.28
cc_13 N_GND_M1013_b N_A_c_312_n 0.00726068f $X=-0.045 $Y=0 $X2=2.36 $Y2=2.405
cc_14 N_GND_M1013_b N_A_c_313_n 0.00580819f $X=-0.045 $Y=0 $X2=2.2 $Y2=2.405
cc_15 N_GND_M1013_b N_A_c_314_n 0.0192889f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.65
cc_16 N_GND_M1013_b N_A_c_315_n 0.0260893f $X=-0.045 $Y=0 $X2=2.435 $Y2=2.33
cc_17 N_GND_M1013_b N_A_c_316_n 0.0164635f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.205
cc_18 N_GND_c_8_p N_A_c_316_n 0.00385579f $X=2.34 $Y=0.755 $X2=2.555 $Y2=1.205
cc_19 N_GND_c_19_p N_A_c_316_n 0.0063578f $X=3.115 $Y=0.152 $X2=2.555 $Y2=1.205
cc_20 N_GND_c_4_p N_A_c_316_n 0.00478641f $X=6.46 $Y=0.19 $X2=2.555 $Y2=1.205
cc_21 N_GND_M1013_b N_A_c_320_n 0.0323293f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.74
cc_22 N_GND_M1013_b N_A_c_321_n 0.00769664f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.28
cc_23 N_GND_M1013_b N_A_c_322_n 0.0103282f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.815
cc_24 N_GND_M1013_b N_A_c_323_n 0.00749597f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.405
cc_25 N_GND_M1013_b N_A_c_324_n 0.0278882f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.4
cc_26 N_GND_c_26_p N_A_c_324_n 0.00148435f $X=5.31 $Y=0.755 $X2=5.155 $Y2=1.4
cc_27 N_GND_M1013_b N_A_c_326_n 0.0189719f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.235
cc_28 N_GND_c_28_p N_A_c_326_n 0.0063578f $X=5.225 $Y=0.152 $X2=5.155 $Y2=1.235
cc_29 N_GND_c_26_p N_A_c_326_n 0.00404581f $X=5.31 $Y=0.755 $X2=5.155 $Y2=1.235
cc_30 N_GND_c_4_p N_A_c_326_n 0.00478641f $X=6.46 $Y=0.19 $X2=5.155 $Y2=1.235
cc_31 N_GND_M1013_b N_A_c_330_n 0.0355583f $X=-0.045 $Y=0 $X2=5.13 $Y2=2.295
cc_32 N_GND_M1013_b N_A_c_331_n 0.010282f $X=-0.045 $Y=0 $X2=5.13 $Y2=2.445
cc_33 N_GND_M1013_b N_A_c_332_n 0.0092608f $X=-0.045 $Y=0 $X2=0.485 $Y2=1.74
cc_34 N_GND_M1013_b N_A_c_333_n 0.0044243f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.485
cc_35 N_GND_c_26_p N_A_c_333_n 0.00269796f $X=5.31 $Y=0.755 $X2=5.155 $Y2=1.485
cc_36 N_GND_M1013_b N_A_c_335_n 0.00242935f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.74
cc_37 N_GND_M1013_b N_A_c_336_n 0.0048047f $X=-0.045 $Y=0 $X2=2.495 $Y2=1.65
cc_38 N_GND_c_8_p N_A_c_336_n 0.00110181f $X=2.34 $Y=0.755 $X2=2.495 $Y2=1.65
cc_39 N_GND_M1013_b N_A_c_338_n 0.0177352f $X=-0.045 $Y=0 $X2=2.35 $Y2=1.74
cc_40 N_GND_M1013_b N_A_c_339_n 0.003389f $X=-0.045 $Y=0 $X2=0.63 $Y2=1.74
cc_41 N_GND_M1013_b N_A_c_340_n 0.0213556f $X=-0.045 $Y=0 $X2=5.01 $Y2=1.74
cc_42 N_GND_M1013_b N_A_c_341_n 0.00137541f $X=-0.045 $Y=0 $X2=2.64 $Y2=1.74
cc_43 N_GND_M1013_b N_A_c_342_n 0.00715594f $X=-0.045 $Y=0 $X2=5.155 $Y2=1.74
cc_44 N_GND_M1013_b N_B_M1001_g 0.0610991f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.85
cc_45 N_GND_c_3_p N_B_M1001_g 0.00385579f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.85
cc_46 N_GND_c_7_p N_B_M1001_g 0.0063578f $X=2.255 $Y=0.152 $X2=0.905 $Y2=0.85
cc_47 N_GND_c_4_p N_B_M1001_g 0.00478641f $X=6.46 $Y=0.19 $X2=0.905 $Y2=0.85
cc_48 N_GND_M1013_b N_B_M1025_g 0.0458794f $X=-0.045 $Y=0 $X2=1.765 $Y2=0.85
cc_49 N_GND_c_7_p N_B_M1025_g 0.0063578f $X=2.255 $Y=0.152 $X2=1.765 $Y2=0.85
cc_50 N_GND_c_4_p N_B_M1025_g 0.00478641f $X=6.46 $Y=0.19 $X2=1.765 $Y2=0.85
cc_51 N_GND_M1013_b N_B_M1012_g 0.0152061f $X=-0.045 $Y=0 $X2=1.765 $Y2=3.235
cc_52 N_GND_M1013_b N_B_M1024_g 0.0297212f $X=-0.045 $Y=0 $X2=2.985 $Y2=0.85
cc_53 N_GND_c_19_p N_B_M1024_g 0.00605374f $X=3.115 $Y=0.152 $X2=2.985 $Y2=0.85
cc_54 N_GND_c_54_p N_B_M1024_g 0.00385579f $X=3.2 $Y=0.615 $X2=2.985 $Y2=0.85
cc_55 N_GND_c_55_p N_B_M1024_g 0.00244503f $X=3.2 $Y=0.7 $X2=2.985 $Y2=0.85
cc_56 N_GND_c_4_p N_B_M1024_g 0.00478641f $X=6.46 $Y=0.19 $X2=2.985 $Y2=0.85
cc_57 N_GND_M1013_b N_B_M1011_g 0.0291906f $X=-0.045 $Y=0 $X2=2.985 $Y2=3.235
cc_58 N_GND_M1013_b N_B_M1017_g 0.0502292f $X=-0.045 $Y=0 $X2=4.275 $Y2=0.85
cc_59 N_GND_c_28_p N_B_M1017_g 0.00470332f $X=5.225 $Y=0.152 $X2=4.275 $Y2=0.85
cc_60 N_GND_c_4_p N_B_M1017_g 0.00478641f $X=6.46 $Y=0.19 $X2=4.275 $Y2=0.85
cc_61 N_GND_M1013_b N_B_M1006_g 0.00556194f $X=-0.045 $Y=0 $X2=4.275 $Y2=3.235
cc_62 N_GND_M1013_b N_B_c_551_n 0.0213189f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.28
cc_63 N_GND_M1013_b N_B_c_552_n 0.040936f $X=-0.045 $Y=0 $X2=2.015 $Y2=1.95
cc_64 N_GND_M1013_b N_B_c_553_n 0.0259722f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.655
cc_65 N_GND_M1013_b N_B_c_554_n 0.0243323f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.135
cc_66 N_GND_M1013_b N_B_c_555_n 0.00674304f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.28
cc_67 N_GND_M1013_b N_B_c_556_n 0.00820793f $X=-0.045 $Y=0 $X2=2.015 $Y2=1.95
cc_68 N_GND_M1013_b N_B_c_557_n 0.00696391f $X=-0.045 $Y=0 $X2=2.975 $Y2=1.655
cc_69 N_GND_M1013_b N_B_c_558_n 7.38055e-19 $X=-0.045 $Y=0 $X2=4.265 $Y2=2.48
cc_70 N_GND_M1013_b N_B_c_559_n 0.00123225f $X=-0.045 $Y=0 $X2=0.485 $Y2=2.28
cc_71 N_GND_M1013_b N_B_c_560_n 0.00256466f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.135
cc_72 N_GND_M1013_b N_B_c_561_n 0.00771729f $X=-0.045 $Y=0 $X2=2.16 $Y2=2.48
cc_73 N_GND_M1013_b N_B_c_562_n 0.00353565f $X=-0.045 $Y=0 $X2=0.63 $Y2=2.48
cc_74 N_GND_M1013_b N_B_c_563_n 0.00166561f $X=-0.045 $Y=0 $X2=2.83 $Y2=2.48
cc_75 N_GND_M1013_b N_B_c_564_n 0.00426493f $X=-0.045 $Y=0 $X2=4.12 $Y2=2.48
cc_76 N_GND_M1013_b N_B_c_565_n 0.00143905f $X=-0.045 $Y=0 $X2=3.12 $Y2=2.48
cc_77 N_GND_M1013_b N_B_c_566_n 0.00169392f $X=-0.045 $Y=0 $X2=4.265 $Y2=2.48
cc_78 N_GND_M1013_b N_CI_M1003_g 0.036914f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.85
cc_79 N_GND_c_7_p N_CI_M1003_g 0.0063578f $X=2.255 $Y=0.152 $X2=1.335 $Y2=0.85
cc_80 N_GND_c_4_p N_CI_M1003_g 0.00478641f $X=6.46 $Y=0.19 $X2=1.335 $Y2=0.85
cc_81 N_GND_M1013_b N_CI_M1020_g 0.0240147f $X=-0.045 $Y=0 $X2=1.335 $Y2=3.235
cc_82 N_GND_M1013_b N_CI_M1014_g 0.0510446f $X=-0.045 $Y=0 $X2=3.415 $Y2=0.85
cc_83 N_GND_c_54_p N_CI_M1014_g 0.00385579f $X=3.2 $Y=0.615 $X2=3.415 $Y2=0.85
cc_84 N_GND_c_28_p N_CI_M1014_g 0.00605374f $X=5.225 $Y=0.152 $X2=3.415 $Y2=0.85
cc_85 N_GND_c_55_p N_CI_M1014_g 0.00244503f $X=3.2 $Y=0.7 $X2=3.415 $Y2=0.85
cc_86 N_GND_c_4_p N_CI_M1014_g 0.00478641f $X=6.46 $Y=0.19 $X2=3.415 $Y2=0.85
cc_87 N_GND_M1013_b N_CI_M1002_g 0.00772364f $X=-0.045 $Y=0 $X2=3.415 $Y2=3.235
cc_88 N_GND_M1013_b N_CI_M1008_g 0.043155f $X=-0.045 $Y=0 $X2=4.685 $Y2=0.85
cc_89 N_GND_c_28_p N_CI_M1008_g 0.0063578f $X=5.225 $Y=0.152 $X2=4.685 $Y2=0.85
cc_90 N_GND_c_4_p N_CI_M1008_g 0.00478641f $X=6.46 $Y=0.19 $X2=4.685 $Y2=0.85
cc_91 N_GND_M1013_b N_CI_M1026_g 0.0163976f $X=-0.045 $Y=0 $X2=4.685 $Y2=3.235
cc_92 N_GND_M1013_b N_CI_c_819_n 0.0281941f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.74
cc_93 N_GND_M1013_b N_CI_c_820_n 0.0264026f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.11
cc_94 N_GND_M1013_b N_CI_c_821_n 0.0264213f $X=-0.045 $Y=0 $X2=4.745 $Y2=1.92
cc_95 N_GND_M1013_b N_CI_c_822_n 0.00449824f $X=-0.045 $Y=0 $X2=1.325 $Y2=1.74
cc_96 N_GND_M1013_b N_CI_c_823_n 0.00277243f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.11
cc_97 N_GND_M1013_b N_CI_c_824_n 0.00259325f $X=-0.045 $Y=0 $X2=4.745 $Y2=1.92
cc_98 N_GND_M1013_b N_CI_c_825_n 0.0134752f $X=-0.045 $Y=0 $X2=3.25 $Y2=2.11
cc_99 N_GND_M1013_b N_CI_c_826_n 0.00577278f $X=-0.045 $Y=0 $X2=1.48 $Y2=2.11
cc_100 N_GND_M1013_b N_CI_c_827_n 0.00807096f $X=-0.045 $Y=0 $X2=4.6 $Y2=2.11
cc_101 N_GND_M1013_b N_CI_c_828_n 0.00194451f $X=-0.045 $Y=0 $X2=3.585 $Y2=2.11
cc_102 N_GND_M1013_b N_CI_c_829_n 0.00568214f $X=-0.045 $Y=0 $X2=4.745 $Y2=2.11
cc_103 N_GND_M1013_b N_CON_M1015_g 0.0212849f $X=-0.045 $Y=0 $X2=3.845 $Y2=0.85
cc_104 N_GND_c_28_p N_CON_M1015_g 0.0063578f $X=5.225 $Y=0.152 $X2=3.845
+ $Y2=0.85
cc_105 N_GND_c_4_p N_CON_M1015_g 0.00478641f $X=6.46 $Y=0.19 $X2=3.845 $Y2=0.85
cc_106 N_GND_M1013_b N_CON_M1005_g 0.0327504f $X=-0.045 $Y=0 $X2=3.845 $Y2=3.235
cc_107 N_GND_M1013_b N_CON_M1023_g 0.088861f $X=-0.045 $Y=0 $X2=6.535 $Y2=0.85
cc_108 N_GND_c_108_p N_CON_M1023_g 0.0067724f $X=6.32 $Y=0.74 $X2=6.535 $Y2=0.85
cc_109 N_GND_c_4_p N_CON_M1023_g 0.00481485f $X=6.46 $Y=0.19 $X2=6.535 $Y2=0.85
cc_110 N_GND_M1013_b N_CON_c_992_n 0.024727f $X=-0.045 $Y=0 $X2=3.845 $Y2=1.455
cc_111 N_GND_M1013_b N_CON_c_993_n 0.0347581f $X=-0.045 $Y=0 $X2=6.41 $Y2=2.26
cc_112 N_GND_M1013_b N_CON_c_994_n 0.00157985f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_113 N_GND_c_7_p N_CON_c_994_n 0.00766062f $X=2.255 $Y=0.152 $X2=1.55
+ $Y2=0.755
cc_114 N_GND_c_4_p N_CON_c_994_n 0.00474629f $X=6.46 $Y=0.19 $X2=1.55 $Y2=0.755
cc_115 N_GND_M1013_b N_CON_c_997_n 0.00832872f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.37
cc_116 N_GND_M1013_b N_CON_c_998_n 0.00668618f $X=-0.045 $Y=0 $X2=6.41 $Y2=2.26
cc_117 N_GND_M1013_b N_CON_c_999_n 0.00296804f $X=-0.045 $Y=0 $X2=1.665 $Y2=1.2
cc_118 N_GND_M1013_b N_CON_c_1000_n 0.00512091f $X=-0.045 $Y=0 $X2=3.845
+ $Y2=1.455
cc_119 N_GND_M1013_b N_CON_c_1001_n 0.0119069f $X=-0.045 $Y=0 $X2=6.41 $Y2=1.37
cc_120 N_GND_c_108_p N_CON_c_1001_n 0.00701922f $X=6.32 $Y=0.74 $X2=6.41
+ $Y2=1.37
cc_121 N_GND_M1013_b N_CON_c_1003_n 0.0249658f $X=-0.045 $Y=0 $X2=3.855 $Y2=1.37
cc_122 N_GND_c_8_p N_CON_c_1003_n 0.00531517f $X=2.34 $Y=0.755 $X2=3.855
+ $Y2=1.37
cc_123 N_GND_M1013_b N_CON_c_1005_n 0.00362533f $X=-0.045 $Y=0 $X2=1.81 $Y2=1.37
cc_124 N_GND_M1013_b N_CON_c_1006_n 0.0424907f $X=-0.045 $Y=0 $X2=5.995 $Y2=1.37
cc_125 N_GND_c_26_p N_CON_c_1006_n 0.00544802f $X=5.31 $Y=0.755 $X2=5.995
+ $Y2=1.37
cc_126 N_GND_M1013_b N_CON_c_1008_n 0.00371124f $X=-0.045 $Y=0 $X2=4.1 $Y2=1.37
cc_127 N_GND_M1013_b CON 0.0204437f $X=-0.045 $Y=0 $X2=6.14 $Y2=1.37
cc_128 N_GND_c_108_p CON 0.00129067f $X=6.32 $Y=0.74 $X2=6.14 $Y2=1.37
cc_129 N_GND_M1013_b N_A_784_115#_M1018_g 0.0715819f $X=-0.045 $Y=0 $X2=5.585
+ $Y2=0.85
cc_130 N_GND_c_26_p N_A_784_115#_M1018_g 0.00727449f $X=5.31 $Y=0.755 $X2=5.585
+ $Y2=0.85
cc_131 N_GND_c_131_p N_A_784_115#_M1018_g 0.00644441f $X=6.235 $Y=0.152
+ $X2=5.585 $Y2=0.85
cc_132 N_GND_c_108_p N_A_784_115#_M1018_g 0.00460621f $X=6.32 $Y=0.74 $X2=5.585
+ $Y2=0.85
cc_133 N_GND_c_4_p N_A_784_115#_M1018_g 0.00481485f $X=6.46 $Y=0.19 $X2=5.585
+ $Y2=0.85
cc_134 N_GND_M1013_b N_A_784_115#_c_1161_n 0.0268825f $X=-0.045 $Y=0 $X2=5.585
+ $Y2=2.275
cc_135 N_GND_M1013_b N_A_784_115#_c_1162_n 0.0078334f $X=-0.045 $Y=0 $X2=3.845
+ $Y2=2.55
cc_136 N_GND_M1013_b N_A_784_115#_c_1163_n 0.00598918f $X=-0.045 $Y=0 $X2=4.225
+ $Y2=1.795
cc_137 N_GND_M1013_b N_A_784_115#_c_1164_n 0.00222689f $X=-0.045 $Y=0 $X2=3.93
+ $Y2=1.795
cc_138 N_GND_M1013_b N_A_784_115#_c_1165_n 0.00566268f $X=-0.045 $Y=0 $X2=4.31
+ $Y2=1.71
cc_139 N_GND_M1013_b N_A_784_115#_c_1166_n 0.00158825f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=0.74
cc_140 N_GND_c_28_p N_A_784_115#_c_1166_n 0.0120982f $X=5.225 $Y=0.152 $X2=4.06
+ $Y2=0.74
cc_141 N_GND_c_4_p N_A_784_115#_c_1166_n 0.0107468f $X=6.46 $Y=0.19 $X2=4.06
+ $Y2=0.74
cc_142 N_GND_M1013_b N_A_784_115#_c_1169_n 0.00781412f $X=-0.045 $Y=0 $X2=5.415
+ $Y2=2.275
cc_143 N_GND_M1013_b N_S_c_1317_n 0.0142036f $X=-0.045 $Y=0 $X2=5.8 $Y2=0.755
cc_144 N_GND_c_131_p N_S_c_1317_n 0.00736239f $X=6.235 $Y=0.152 $X2=5.8
+ $Y2=0.755
cc_145 N_GND_c_108_p N_S_c_1317_n 0.0140971f $X=6.32 $Y=0.74 $X2=5.8 $Y2=0.755
cc_146 N_GND_c_4_p N_S_c_1317_n 0.00476261f $X=6.46 $Y=0.19 $X2=5.8 $Y2=0.755
cc_147 N_GND_M1013_b N_S_c_1321_n 0.0133222f $X=-0.045 $Y=0 $X2=5.925 $Y2=2.685
cc_148 N_GND_M1013_b N_S_c_1322_n 0.0110471f $X=-0.045 $Y=0 $X2=5.925 $Y2=1.74
cc_149 N_GND_M1013_b N_CO_c_1368_n 0.0677803f $X=-0.045 $Y=0 $X2=6.75 $Y2=0.755
cc_150 N_GND_c_4_p N_CO_c_1368_n 0.00476261f $X=6.46 $Y=0.19 $X2=6.75 $Y2=0.755
cc_151 N_GND_M1013_b CO 0.00667411f $X=-0.045 $Y=0 $X2=6.75 $Y2=2.48
cc_152 N_GND_M1013_b N_A_27_115#_c_1384_n 0.0015601f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_153 N_GND_c_2_p N_A_27_115#_c_1384_n 0.00735421f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_154 N_GND_c_4_p N_A_27_115#_c_1384_n 0.00476028f $X=6.46 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_155 N_GND_M1013_d N_A_27_115#_c_1387_n 0.00176461f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.16
cc_156 N_GND_M1013_b N_A_27_115#_c_1387_n 0.00866634f $X=-0.045 $Y=0 $X2=1.035
+ $Y2=1.16
cc_157 N_GND_c_3_p N_A_27_115#_c_1387_n 0.0135055f $X=0.69 $Y=0.74 $X2=1.035
+ $Y2=1.16
cc_158 N_GND_M1013_b N_A_27_115#_c_1390_n 0.00158594f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.755
cc_159 N_GND_c_3_p N_A_27_115#_c_1390_n 2.23682e-19 $X=0.69 $Y=0.74 $X2=1.12
+ $Y2=0.755
cc_160 N_GND_c_7_p N_A_27_115#_c_1390_n 0.00775164f $X=2.255 $Y=0.152 $X2=1.12
+ $Y2=0.755
cc_161 N_GND_c_4_p N_A_27_115#_c_1390_n 0.00477923f $X=6.46 $Y=0.19 $X2=1.12
+ $Y2=0.755
cc_162 N_GND_M1013_b N_A_27_115#_c_1394_n 0.0107358f $X=-0.045 $Y=0 $X2=0.262
+ $Y2=1.16
cc_163 N_GND_M1013_b N_A_526_115#_c_1410_n 0.00158398f $X=-0.045 $Y=0 $X2=2.77
+ $Y2=0.755
cc_164 N_GND_c_8_p N_A_526_115#_c_1410_n 2.23682e-19 $X=2.34 $Y=0.755 $X2=2.77
+ $Y2=0.755
cc_165 N_GND_c_19_p N_A_526_115#_c_1410_n 0.00792421f $X=3.115 $Y=0.152 $X2=2.77
+ $Y2=0.755
cc_166 N_GND_c_54_p N_A_526_115#_c_1410_n 2.23682e-19 $X=3.2 $Y=0.615 $X2=2.77
+ $Y2=0.755
cc_167 N_GND_c_4_p N_A_526_115#_c_1410_n 0.00476846f $X=6.46 $Y=0.19 $X2=2.77
+ $Y2=0.755
cc_168 N_GND_M1024_d N_A_526_115#_c_1415_n 0.00207687f $X=3.06 $Y=0.575
+ $X2=3.545 $Y2=1.115
cc_169 N_GND_M1013_b N_A_526_115#_c_1415_n 0.00587809f $X=-0.045 $Y=0 $X2=3.545
+ $Y2=1.115
cc_170 N_GND_c_55_p N_A_526_115#_c_1415_n 0.0115859f $X=3.2 $Y=0.7 $X2=3.545
+ $Y2=1.115
cc_171 N_GND_M1013_b N_A_526_115#_c_1418_n 0.00283355f $X=-0.045 $Y=0 $X2=2.855
+ $Y2=1.115
cc_172 N_GND_M1013_b N_A_526_115#_c_1419_n 0.00158398f $X=-0.045 $Y=0 $X2=3.63
+ $Y2=0.755
cc_173 N_GND_c_54_p N_A_526_115#_c_1419_n 2.23682e-19 $X=3.2 $Y=0.615 $X2=3.63
+ $Y2=0.755
cc_174 N_GND_c_28_p N_A_526_115#_c_1419_n 0.00770991f $X=5.225 $Y=0.152 $X2=3.63
+ $Y2=0.755
cc_175 N_GND_c_4_p N_A_526_115#_c_1419_n 0.00476846f $X=6.46 $Y=0.19 $X2=3.63
+ $Y2=0.755
cc_176 N_VDD_M1000_b N_A_M1000_g 0.0259953f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_177 N_VDD_c_177_p N_A_M1000_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_178 N_VDD_c_178_p N_A_M1000_g 0.00337744f $X=0.69 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_179 N_VDD_c_179_p N_A_M1000_g 0.00468827f $X=6.46 $Y=4.25 $X2=0.475 $Y2=3.235
cc_180 N_VDD_M1000_b N_A_c_347_n 0.0154424f $X=-0.045 $Y=2.425 $X2=2.125
+ $Y2=2.48
cc_181 N_VDD_c_181_p N_A_c_347_n 0.00606474f $X=2.255 $Y=4.287 $X2=2.125
+ $Y2=2.48
cc_182 N_VDD_c_182_p N_A_c_347_n 0.00337744f $X=2.34 $Y=3.295 $X2=2.125 $Y2=2.48
cc_183 N_VDD_c_179_p N_A_c_347_n 0.00468827f $X=6.46 $Y=4.25 $X2=2.125 $Y2=2.48
cc_184 N_VDD_M1000_b N_A_c_312_n 0.00289837f $X=-0.045 $Y=2.425 $X2=2.36
+ $Y2=2.405
cc_185 N_VDD_c_182_p N_A_c_312_n 5.81807e-19 $X=2.34 $Y=3.295 $X2=2.36 $Y2=2.405
cc_186 N_VDD_M1000_b N_A_c_313_n 0.00143424f $X=-0.045 $Y=2.425 $X2=2.2
+ $Y2=2.405
cc_187 N_VDD_M1000_b N_A_c_354_n 0.0163636f $X=-0.045 $Y=2.425 $X2=2.555
+ $Y2=2.48
cc_188 N_VDD_c_182_p N_A_c_354_n 0.00337744f $X=2.34 $Y=3.295 $X2=2.555 $Y2=2.48
cc_189 N_VDD_c_189_p N_A_c_354_n 0.00606474f $X=3.115 $Y=4.287 $X2=2.555
+ $Y2=2.48
cc_190 N_VDD_c_179_p N_A_c_354_n 0.00468827f $X=6.46 $Y=4.25 $X2=2.555 $Y2=2.48
cc_191 N_VDD_M1000_b N_A_M1021_g 0.0203595f $X=-0.045 $Y=2.425 $X2=5.095
+ $Y2=3.235
cc_192 N_VDD_c_192_p N_A_M1021_g 0.0061469f $X=5.225 $Y=4.287 $X2=5.095
+ $Y2=3.235
cc_193 N_VDD_c_193_p N_A_M1021_g 0.0037786f $X=5.31 $Y=3.635 $X2=5.095 $Y2=3.235
cc_194 N_VDD_c_179_p N_A_M1021_g 0.00471609f $X=6.46 $Y=4.25 $X2=5.095 $Y2=3.235
cc_195 N_VDD_M1000_b N_A_c_323_n 0.00319137f $X=-0.045 $Y=2.425 $X2=2.555
+ $Y2=2.405
cc_196 N_VDD_M1000_b N_A_c_331_n 0.0032153f $X=-0.045 $Y=2.425 $X2=5.13
+ $Y2=2.445
cc_197 N_VDD_M1000_b N_B_M1019_g 0.0182122f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_198 N_VDD_c_178_p N_B_M1019_g 0.00337744f $X=0.69 $Y=3.635 $X2=0.905
+ $Y2=3.235
cc_199 N_VDD_c_181_p N_B_M1019_g 0.00606474f $X=2.255 $Y=4.287 $X2=0.905
+ $Y2=3.235
cc_200 N_VDD_c_179_p N_B_M1019_g 0.00468827f $X=6.46 $Y=4.25 $X2=0.905 $Y2=3.235
cc_201 N_VDD_M1000_b N_B_M1012_g 0.018554f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=3.235
cc_202 N_VDD_c_181_p N_B_M1012_g 0.0061469f $X=2.255 $Y=4.287 $X2=1.765
+ $Y2=3.235
cc_203 N_VDD_c_182_p N_B_M1012_g 0.00177739f $X=2.34 $Y=3.295 $X2=1.765
+ $Y2=3.235
cc_204 N_VDD_c_179_p N_B_M1012_g 0.00471609f $X=6.46 $Y=4.25 $X2=1.765 $Y2=3.235
cc_205 N_VDD_M1000_b N_B_M1011_g 0.0193458f $X=-0.045 $Y=2.425 $X2=2.985
+ $Y2=3.235
cc_206 N_VDD_c_182_p N_B_M1011_g 4.9048e-19 $X=2.34 $Y=3.295 $X2=2.985 $Y2=3.235
cc_207 N_VDD_c_189_p N_B_M1011_g 0.0061469f $X=3.115 $Y=4.287 $X2=2.985
+ $Y2=3.235
cc_208 N_VDD_c_208_p N_B_M1011_g 0.00332149f $X=3.2 $Y=3.7 $X2=2.985 $Y2=3.235
cc_209 N_VDD_c_179_p N_B_M1011_g 0.00471609f $X=6.46 $Y=4.25 $X2=2.985 $Y2=3.235
cc_210 N_VDD_M1000_b N_B_M1006_g 0.0190171f $X=-0.045 $Y=2.425 $X2=4.275
+ $Y2=3.235
cc_211 N_VDD_c_192_p N_B_M1006_g 0.0061469f $X=5.225 $Y=4.287 $X2=4.275
+ $Y2=3.235
cc_212 N_VDD_c_179_p N_B_M1006_g 0.00471609f $X=6.46 $Y=4.25 $X2=4.275 $Y2=3.235
cc_213 N_VDD_M1000_b N_B_c_551_n 0.00509255f $X=-0.045 $Y=2.425 $X2=0.895
+ $Y2=2.28
cc_214 N_VDD_M1000_b N_B_c_584_n 0.00204928f $X=-0.045 $Y=2.425 $X2=2.1 $Y2=2.48
cc_215 N_VDD_M1000_b N_B_c_585_n 0.00243177f $X=-0.045 $Y=2.425 $X2=2.305
+ $Y2=2.48
cc_216 N_VDD_c_182_p N_B_c_585_n 0.00305822f $X=2.34 $Y=3.295 $X2=2.305 $Y2=2.48
cc_217 N_VDD_M1000_b N_B_c_557_n 0.00125334f $X=-0.045 $Y=2.425 $X2=2.975
+ $Y2=1.655
cc_218 N_VDD_M1000_b N_B_c_558_n 7.43789e-19 $X=-0.045 $Y=2.425 $X2=4.265
+ $Y2=2.48
cc_219 N_VDD_M1000_b N_B_c_559_n 0.00190563f $X=-0.045 $Y=2.425 $X2=0.485
+ $Y2=2.28
cc_220 N_VDD_M1000_b N_B_c_561_n 0.0151656f $X=-0.045 $Y=2.425 $X2=2.16 $Y2=2.48
cc_221 N_VDD_M1000_b N_B_c_562_n 0.00845167f $X=-0.045 $Y=2.425 $X2=0.63
+ $Y2=2.48
cc_222 N_VDD_M1000_b N_B_c_563_n 0.00454131f $X=-0.045 $Y=2.425 $X2=2.83
+ $Y2=2.48
cc_223 N_VDD_M1000_b N_B_c_593_n 0.00497303f $X=-0.045 $Y=2.425 $X2=2.45
+ $Y2=2.48
cc_224 N_VDD_c_182_p N_B_c_593_n 0.00464167f $X=2.34 $Y=3.295 $X2=2.45 $Y2=2.48
cc_225 N_VDD_M1000_b N_B_c_564_n 0.00819904f $X=-0.045 $Y=2.425 $X2=4.12
+ $Y2=2.48
cc_226 N_VDD_M1000_b N_B_c_565_n 0.00220137f $X=-0.045 $Y=2.425 $X2=3.12
+ $Y2=2.48
cc_227 N_VDD_M1000_b N_B_c_566_n 0.00404898f $X=-0.045 $Y=2.425 $X2=4.265
+ $Y2=2.48
cc_228 N_VDD_M1000_b N_CI_M1020_g 0.0197242f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=3.235
cc_229 N_VDD_c_178_p N_CI_M1020_g 4.9048e-19 $X=0.69 $Y=3.635 $X2=1.335
+ $Y2=3.235
cc_230 N_VDD_c_181_p N_CI_M1020_g 0.0061469f $X=2.255 $Y=4.287 $X2=1.335
+ $Y2=3.235
cc_231 N_VDD_c_179_p N_CI_M1020_g 0.00471609f $X=6.46 $Y=4.25 $X2=1.335
+ $Y2=3.235
cc_232 N_VDD_M1000_b N_CI_M1002_g 0.0196567f $X=-0.045 $Y=2.425 $X2=3.415
+ $Y2=3.235
cc_233 N_VDD_c_208_p N_CI_M1002_g 0.00332149f $X=3.2 $Y=3.7 $X2=3.415 $Y2=3.235
cc_234 N_VDD_c_192_p N_CI_M1002_g 0.0061469f $X=5.225 $Y=4.287 $X2=3.415
+ $Y2=3.235
cc_235 N_VDD_c_179_p N_CI_M1002_g 0.00471609f $X=6.46 $Y=4.25 $X2=3.415
+ $Y2=3.235
cc_236 N_VDD_M1000_b N_CI_M1026_g 0.0206788f $X=-0.045 $Y=2.425 $X2=4.685
+ $Y2=3.235
cc_237 N_VDD_c_192_p N_CI_M1026_g 0.0061469f $X=5.225 $Y=4.287 $X2=4.685
+ $Y2=3.235
cc_238 N_VDD_c_179_p N_CI_M1026_g 0.00471609f $X=6.46 $Y=4.25 $X2=4.685
+ $Y2=3.235
cc_239 N_VDD_M1000_b N_CON_M1005_g 0.0189866f $X=-0.045 $Y=2.425 $X2=3.845
+ $Y2=3.235
cc_240 N_VDD_c_192_p N_CON_M1005_g 0.0061469f $X=5.225 $Y=4.287 $X2=3.845
+ $Y2=3.235
cc_241 N_VDD_c_179_p N_CON_M1005_g 0.00471609f $X=6.46 $Y=4.25 $X2=3.845
+ $Y2=3.235
cc_242 N_VDD_M1000_b N_CON_M1010_g 0.0292927f $X=-0.045 $Y=2.425 $X2=6.535
+ $Y2=3.235
cc_243 N_VDD_c_243_p N_CON_M1010_g 0.00675484f $X=6.32 $Y=2.955 $X2=6.535
+ $Y2=3.235
cc_244 N_VDD_c_244_p N_CON_M1010_g 0.0061469f $X=6.46 $Y=4.22 $X2=6.535
+ $Y2=3.235
cc_245 N_VDD_c_179_p N_CON_M1010_g 0.00471609f $X=6.46 $Y=4.25 $X2=6.535
+ $Y2=3.235
cc_246 N_VDD_M1000_b N_CON_c_993_n 0.00517554f $X=-0.045 $Y=2.425 $X2=6.41
+ $Y2=2.26
cc_247 N_VDD_c_243_p N_CON_c_993_n 0.00254427f $X=6.32 $Y=2.955 $X2=6.41
+ $Y2=2.26
cc_248 N_VDD_M1000_b N_CON_c_1020_n 0.00155118f $X=-0.045 $Y=2.425 $X2=1.55
+ $Y2=3.295
cc_249 N_VDD_c_181_p N_CON_c_1020_n 0.00737727f $X=2.255 $Y=4.287 $X2=1.55
+ $Y2=3.295
cc_250 N_VDD_c_179_p N_CON_c_1020_n 0.00475776f $X=6.46 $Y=4.25 $X2=1.55
+ $Y2=3.295
cc_251 N_VDD_M1000_b N_CON_c_997_n 0.0015365f $X=-0.045 $Y=2.425 $X2=1.665
+ $Y2=1.37
cc_252 N_VDD_M1000_b N_CON_c_998_n 0.00319259f $X=-0.045 $Y=2.425 $X2=6.41
+ $Y2=2.26
cc_253 N_VDD_c_243_p N_CON_c_998_n 0.00436457f $X=6.32 $Y=2.955 $X2=6.41
+ $Y2=2.26
cc_254 N_VDD_M1000_b N_CON_c_1026_n 0.00220635f $X=-0.045 $Y=2.425 $X2=1.665
+ $Y2=2.637
cc_255 N_VDD_M1000_b N_A_784_115#_M1007_g 0.0227865f $X=-0.045 $Y=2.425
+ $X2=5.585 $Y2=3.235
cc_256 N_VDD_c_193_p N_A_784_115#_M1007_g 0.00721426f $X=5.31 $Y=3.635 $X2=5.585
+ $Y2=3.235
cc_257 N_VDD_c_257_p N_A_784_115#_M1007_g 0.0061469f $X=6.235 $Y=4.287 $X2=5.585
+ $Y2=3.235
cc_258 N_VDD_c_243_p N_A_784_115#_M1007_g 0.00540522f $X=6.32 $Y=2.955 $X2=5.585
+ $Y2=3.235
cc_259 N_VDD_c_179_p N_A_784_115#_M1007_g 0.00471609f $X=6.46 $Y=4.25 $X2=5.585
+ $Y2=3.235
cc_260 N_VDD_M1000_b N_A_784_115#_c_1161_n 0.0046837f $X=-0.045 $Y=2.425
+ $X2=5.585 $Y2=2.275
cc_261 N_VDD_M1000_b N_A_784_115#_c_1162_n 0.0021798f $X=-0.045 $Y=2.425
+ $X2=3.845 $Y2=2.55
cc_262 N_VDD_M1000_b N_A_784_115#_c_1177_n 8.33439e-19 $X=-0.045 $Y=2.425
+ $X2=4.06 $Y2=2.94
cc_263 N_VDD_M1000_b N_A_784_115#_c_1178_n 0.00155118f $X=-0.045 $Y=2.425
+ $X2=4.06 $Y2=3.295
cc_264 N_VDD_c_192_p N_A_784_115#_c_1178_n 0.0075556f $X=5.225 $Y=4.287 $X2=4.06
+ $Y2=3.295
cc_265 N_VDD_c_179_p N_A_784_115#_c_1178_n 0.00475776f $X=6.46 $Y=4.25 $X2=4.06
+ $Y2=3.295
cc_266 N_VDD_M1021_d N_A_784_115#_c_1181_n 0.0101125f $X=5.17 $Y=2.605 $X2=5.33
+ $Y2=2.855
cc_267 N_VDD_c_193_p N_A_784_115#_c_1181_n 0.00666443f $X=5.31 $Y=3.635 $X2=5.33
+ $Y2=2.855
cc_268 N_VDD_M1021_d N_A_784_115#_c_1183_n 0.00273928f $X=5.17 $Y=2.605
+ $X2=5.415 $Y2=2.77
cc_269 N_VDD_M1000_b N_A_784_115#_c_1183_n 0.00271341f $X=-0.045 $Y=2.425
+ $X2=5.415 $Y2=2.77
cc_270 N_VDD_M1000_b N_A_784_115#_c_1169_n 6.60644e-19 $X=-0.045 $Y=2.425
+ $X2=5.415 $Y2=2.275
cc_271 N_VDD_M1000_b N_A_27_521#_c_1285_n 0.00156053f $X=-0.045 $Y=2.425
+ $X2=0.26 $Y2=3.295
cc_272 N_VDD_c_177_p N_A_27_521#_c_1285_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=3.295
cc_273 N_VDD_c_179_p N_A_27_521#_c_1285_n 0.00476261f $X=6.46 $Y=4.25 $X2=0.26
+ $Y2=3.295
cc_274 N_VDD_M1000_d N_A_27_521#_c_1288_n 0.005183f $X=0.55 $Y=2.605 $X2=1.035
+ $Y2=2.98
cc_275 N_VDD_c_178_p N_A_27_521#_c_1288_n 0.00809661f $X=0.69 $Y=3.635 $X2=1.035
+ $Y2=2.98
cc_276 N_VDD_M1000_b N_A_27_521#_c_1290_n 0.00155118f $X=-0.045 $Y=2.425
+ $X2=1.12 $Y2=3.295
cc_277 N_VDD_c_181_p N_A_27_521#_c_1290_n 0.00734006f $X=2.255 $Y=4.287 $X2=1.12
+ $Y2=3.295
cc_278 N_VDD_c_179_p N_A_27_521#_c_1290_n 0.00475776f $X=6.46 $Y=4.25 $X2=1.12
+ $Y2=3.295
cc_279 N_VDD_M1011_d N_A_526_521#_c_1300_n 0.0052102f $X=3.06 $Y=2.605 $X2=3.545
+ $Y2=3.23
cc_280 N_VDD_c_208_p N_A_526_521#_c_1300_n 0.0111505f $X=3.2 $Y=3.7 $X2=3.545
+ $Y2=3.23
cc_281 N_VDD_M1000_b N_A_526_521#_c_1302_n 0.00155282f $X=-0.045 $Y=2.425
+ $X2=3.63 $Y2=3.55
cc_282 N_VDD_c_192_p N_A_526_521#_c_1302_n 0.00737161f $X=5.225 $Y=4.287
+ $X2=3.63 $Y2=3.55
cc_283 N_VDD_c_179_p N_A_526_521#_c_1302_n 0.00476677f $X=6.46 $Y=4.25 $X2=3.63
+ $Y2=3.55
cc_284 N_VDD_M1000_b N_A_526_521#_c_1305_n 0.00155118f $X=-0.045 $Y=2.425
+ $X2=2.77 $Y2=3.295
cc_285 N_VDD_c_189_p N_A_526_521#_c_1305_n 0.0075556f $X=3.115 $Y=4.287 $X2=2.77
+ $Y2=3.295
cc_286 N_VDD_c_179_p N_A_526_521#_c_1305_n 0.00475776f $X=6.46 $Y=4.25 $X2=2.77
+ $Y2=3.295
cc_287 N_VDD_M1000_b N_S_c_1323_n 0.00156053f $X=-0.045 $Y=2.425 $X2=5.8
+ $Y2=3.295
cc_288 N_VDD_c_257_p N_S_c_1323_n 0.00736239f $X=6.235 $Y=4.287 $X2=5.8
+ $Y2=3.295
cc_289 N_VDD_c_243_p N_S_c_1323_n 0.0415754f $X=6.32 $Y=2.955 $X2=5.8 $Y2=3.295
cc_290 N_VDD_c_179_p N_S_c_1323_n 0.00476261f $X=6.46 $Y=4.25 $X2=5.8 $Y2=3.295
cc_291 N_VDD_M1000_b N_S_c_1321_n 0.00566411f $X=-0.045 $Y=2.425 $X2=5.925
+ $Y2=2.685
cc_292 N_VDD_M1000_b N_S_c_1328_n 0.0046764f $X=-0.045 $Y=2.425 $X2=5.925
+ $Y2=2.77
cc_293 N_VDD_c_243_p N_S_c_1328_n 0.00741835f $X=6.32 $Y=2.955 $X2=5.925
+ $Y2=2.77
cc_294 N_VDD_M1000_b S 0.00175337f $X=-0.045 $Y=2.425 $X2=5.8 $Y2=2.855
cc_295 N_VDD_c_243_p S 0.00402101f $X=6.32 $Y=2.955 $X2=5.8 $Y2=2.855
cc_296 N_VDD_M1000_b N_CO_c_1368_n 0.00679494f $X=-0.045 $Y=2.425 $X2=6.75
+ $Y2=0.755
cc_297 N_VDD_c_244_p N_CO_c_1368_n 0.00757793f $X=6.46 $Y=4.22 $X2=6.75
+ $Y2=0.755
cc_298 N_VDD_c_179_p N_CO_c_1368_n 0.00476261f $X=6.46 $Y=4.25 $X2=6.75
+ $Y2=0.755
cc_299 N_VDD_M1000_b CO 0.0109934f $X=-0.045 $Y=2.425 $X2=6.75 $Y2=2.48
cc_300 N_A_M1013_g N_B_M1001_g 0.0360289f $X=0.475 $Y=0.85 $X2=0.905 $Y2=0.85
cc_301 N_A_M1000_g N_B_M1001_g 0.0100215f $X=0.475 $Y=3.235 $X2=0.905 $Y2=0.85
cc_302 N_A_c_320_n N_B_M1001_g 0.0220665f $X=0.485 $Y=1.74 $X2=0.905 $Y2=0.85
cc_303 N_A_c_332_n N_B_M1001_g 0.00124108f $X=0.485 $Y=1.74 $X2=0.905 $Y2=0.85
cc_304 N_A_c_338_n N_B_M1001_g 0.00637076f $X=2.35 $Y=1.74 $X2=0.905 $Y2=0.85
cc_305 N_A_c_339_n N_B_M1001_g 8.6716e-19 $X=0.63 $Y=1.74 $X2=0.905 $Y2=0.85
cc_306 N_A_M1000_g N_B_M1019_g 0.0512896f $X=0.475 $Y=3.235 $X2=0.905 $Y2=3.235
cc_307 N_A_c_305_n N_B_M1025_g 0.058151f $X=2.125 $Y=1.205 $X2=1.765 $Y2=0.85
cc_308 N_A_c_314_n N_B_M1025_g 0.00743119f $X=2.495 $Y=1.65 $X2=1.765 $Y2=0.85
cc_309 N_A_c_336_n N_B_M1025_g 0.00118981f $X=2.495 $Y=1.65 $X2=1.765 $Y2=0.85
cc_310 N_A_c_338_n N_B_M1025_g 0.00215929f $X=2.35 $Y=1.74 $X2=1.765 $Y2=0.85
cc_311 N_A_c_313_n N_B_M1012_g 0.100647f $X=2.2 $Y=2.405 $X2=1.765 $Y2=3.235
cc_312 N_A_c_315_n N_B_M1012_g 0.00253344f $X=2.435 $Y=2.33 $X2=1.765 $Y2=3.235
cc_313 N_A_c_316_n N_B_M1024_g 0.0317886f $X=2.555 $Y=1.205 $X2=2.985 $Y2=0.85
cc_314 N_A_c_315_n N_B_M1011_g 0.0144389f $X=2.435 $Y=2.33 $X2=2.985 $Y2=3.235
cc_315 N_A_c_323_n N_B_M1011_g 0.0443538f $X=2.555 $Y=2.405 $X2=2.985 $Y2=3.235
cc_316 N_A_c_340_n N_B_M1017_g 6.15167e-19 $X=5.01 $Y=1.74 $X2=4.275 $Y2=0.85
cc_317 N_A_M1000_g N_B_c_551_n 0.0215713f $X=0.475 $Y=3.235 $X2=0.895 $Y2=2.28
cc_318 N_A_c_338_n N_B_c_551_n 0.00277106f $X=2.35 $Y=1.74 $X2=0.895 $Y2=2.28
cc_319 N_A_c_311_n N_B_c_552_n 0.00301833f $X=2.2 $Y=1.28 $X2=2.015 $Y2=1.95
cc_320 N_A_c_313_n N_B_c_552_n 0.00685208f $X=2.2 $Y=2.405 $X2=2.015 $Y2=1.95
cc_321 N_A_c_322_n N_B_c_552_n 0.0226249f $X=2.495 $Y=1.815 $X2=2.015 $Y2=1.95
cc_322 N_A_c_338_n N_B_c_552_n 0.00491533f $X=2.35 $Y=1.74 $X2=2.015 $Y2=1.95
cc_323 N_A_c_341_n N_B_c_552_n 4.52938e-19 $X=2.64 $Y=1.74 $X2=2.015 $Y2=1.95
cc_324 N_A_c_314_n N_B_c_553_n 0.0215223f $X=2.495 $Y=1.65 $X2=2.975 $Y2=1.655
cc_325 N_A_c_336_n N_B_c_553_n 0.0012108f $X=2.495 $Y=1.65 $X2=2.975 $Y2=1.655
cc_326 N_A_c_340_n N_B_c_553_n 0.00295199f $X=5.01 $Y=1.74 $X2=2.975 $Y2=1.655
cc_327 N_A_M1000_g N_B_c_555_n 4.31787e-19 $X=0.475 $Y=3.235 $X2=0.895 $Y2=2.28
cc_328 N_A_c_320_n N_B_c_555_n 0.00106522f $X=0.485 $Y=1.74 $X2=0.895 $Y2=2.28
cc_329 N_A_c_332_n N_B_c_555_n 0.00221967f $X=0.485 $Y=1.74 $X2=0.895 $Y2=2.28
cc_330 N_A_c_338_n N_B_c_555_n 0.0145415f $X=2.35 $Y=1.74 $X2=0.895 $Y2=2.28
cc_331 N_A_c_339_n N_B_c_555_n 5.69327e-19 $X=0.63 $Y=1.74 $X2=0.895 $Y2=2.28
cc_332 N_A_c_311_n N_B_c_556_n 4.3541e-19 $X=2.2 $Y=1.28 $X2=2.015 $Y2=1.95
cc_333 N_A_c_313_n N_B_c_556_n 0.00293439f $X=2.2 $Y=2.405 $X2=2.015 $Y2=1.95
cc_334 N_A_c_315_n N_B_c_556_n 0.00214417f $X=2.435 $Y=2.33 $X2=2.015 $Y2=1.95
cc_335 N_A_c_322_n N_B_c_556_n 0.00214621f $X=2.495 $Y=1.815 $X2=2.015 $Y2=1.95
cc_336 N_A_c_336_n N_B_c_556_n 0.00130269f $X=2.495 $Y=1.65 $X2=2.015 $Y2=1.95
cc_337 N_A_c_338_n N_B_c_556_n 0.00702452f $X=2.35 $Y=1.74 $X2=2.015 $Y2=1.95
cc_338 N_A_c_341_n N_B_c_556_n 0.00124164f $X=2.64 $Y=1.74 $X2=2.015 $Y2=1.95
cc_339 N_A_c_347_n N_B_c_584_n 0.00199314f $X=2.125 $Y=2.48 $X2=2.1 $Y2=2.48
cc_340 N_A_c_313_n N_B_c_584_n 8.16151e-19 $X=2.2 $Y=2.405 $X2=2.1 $Y2=2.48
cc_341 N_A_c_347_n N_B_c_585_n 0.0038234f $X=2.125 $Y=2.48 $X2=2.305 $Y2=2.48
cc_342 N_A_c_312_n N_B_c_585_n 0.00501184f $X=2.36 $Y=2.405 $X2=2.305 $Y2=2.48
cc_343 N_A_c_313_n N_B_c_585_n 0.00255742f $X=2.2 $Y=2.405 $X2=2.305 $Y2=2.48
cc_344 N_A_c_354_n N_B_c_585_n 7.94851e-19 $X=2.555 $Y=2.48 $X2=2.305 $Y2=2.48
cc_345 N_A_c_323_n N_B_c_585_n 0.00240608f $X=2.555 $Y=2.405 $X2=2.305 $Y2=2.48
cc_346 N_A_c_336_n N_B_c_585_n 6.12315e-19 $X=2.495 $Y=1.65 $X2=2.305 $Y2=2.48
cc_347 N_A_c_314_n N_B_c_557_n 7.07742e-19 $X=2.495 $Y=1.65 $X2=2.975 $Y2=1.655
cc_348 N_A_c_315_n N_B_c_557_n 0.00776148f $X=2.435 $Y=2.33 $X2=2.975 $Y2=1.655
cc_349 N_A_c_322_n N_B_c_557_n 2.63486e-19 $X=2.495 $Y=1.815 $X2=2.975 $Y2=1.655
cc_350 N_A_c_323_n N_B_c_557_n 0.00215473f $X=2.555 $Y=2.405 $X2=2.975 $Y2=1.655
cc_351 N_A_c_336_n N_B_c_557_n 0.0122325f $X=2.495 $Y=1.65 $X2=2.975 $Y2=1.655
cc_352 N_A_c_340_n N_B_c_557_n 0.0144678f $X=5.01 $Y=1.74 $X2=2.975 $Y2=1.655
cc_353 N_A_c_341_n N_B_c_557_n 0.00154249f $X=2.64 $Y=1.74 $X2=2.975 $Y2=1.655
cc_354 N_A_M1000_g N_B_c_559_n 0.0206879f $X=0.475 $Y=3.235 $X2=0.485 $Y2=2.28
cc_355 N_A_c_320_n N_B_c_559_n 4.18273e-19 $X=0.485 $Y=1.74 $X2=0.485 $Y2=2.28
cc_356 N_A_c_332_n N_B_c_559_n 0.00433553f $X=0.485 $Y=1.74 $X2=0.485 $Y2=2.28
cc_357 N_A_c_339_n N_B_c_559_n 0.001558f $X=0.63 $Y=1.74 $X2=0.485 $Y2=2.28
cc_358 N_A_c_340_n N_B_c_560_n 8.54952e-19 $X=5.01 $Y=1.74 $X2=4.265 $Y2=2.135
cc_359 N_A_c_347_n N_B_c_561_n 0.00455994f $X=2.125 $Y=2.48 $X2=2.16 $Y2=2.48
cc_360 N_A_c_313_n N_B_c_561_n 2.67951e-19 $X=2.2 $Y=2.405 $X2=2.16 $Y2=2.48
cc_361 N_A_M1000_g N_B_c_562_n 0.00373503f $X=0.475 $Y=3.235 $X2=0.63 $Y2=2.48
cc_362 N_A_c_320_n N_B_c_562_n 7.28634e-19 $X=0.485 $Y=1.74 $X2=0.63 $Y2=2.48
cc_363 N_A_c_332_n N_B_c_562_n 0.0010849f $X=0.485 $Y=1.74 $X2=0.63 $Y2=2.48
cc_364 N_A_c_339_n N_B_c_562_n 0.0141286f $X=0.63 $Y=1.74 $X2=0.63 $Y2=2.48
cc_365 N_A_c_354_n N_B_c_563_n 0.0078404f $X=2.555 $Y=2.48 $X2=2.83 $Y2=2.48
cc_366 N_A_c_323_n N_B_c_563_n 0.00206361f $X=2.555 $Y=2.405 $X2=2.83 $Y2=2.48
cc_367 N_A_c_347_n N_B_c_593_n 0.00213958f $X=2.125 $Y=2.48 $X2=2.45 $Y2=2.48
cc_368 N_A_c_312_n N_B_c_593_n 6.80224e-19 $X=2.36 $Y=2.405 $X2=2.45 $Y2=2.48
cc_369 N_A_c_313_n N_B_c_593_n 3.98925e-19 $X=2.2 $Y=2.405 $X2=2.45 $Y2=2.48
cc_370 N_A_c_354_n N_B_c_593_n 2.0394e-19 $X=2.555 $Y=2.48 $X2=2.45 $Y2=2.48
cc_371 N_A_c_323_n N_B_c_593_n 9.60339e-19 $X=2.555 $Y=2.405 $X2=2.45 $Y2=2.48
cc_372 N_A_c_340_n N_CI_M1014_g 0.00513502f $X=5.01 $Y=1.74 $X2=3.415 $Y2=0.85
cc_373 N_A_c_326_n N_CI_M1008_g 0.0579501f $X=5.155 $Y=1.235 $X2=4.685 $Y2=0.85
cc_374 N_A_c_330_n N_CI_M1008_g 0.00689222f $X=5.13 $Y=2.295 $X2=4.685 $Y2=0.85
cc_375 N_A_c_333_n N_CI_M1008_g 0.00127753f $X=5.155 $Y=1.485 $X2=4.685 $Y2=0.85
cc_376 N_A_c_335_n N_CI_M1008_g 0.00162427f $X=5.155 $Y=1.74 $X2=4.685 $Y2=0.85
cc_377 N_A_c_340_n N_CI_M1008_g 0.00280998f $X=5.01 $Y=1.74 $X2=4.685 $Y2=0.85
cc_378 N_A_c_342_n N_CI_M1008_g 4.41129e-19 $X=5.155 $Y=1.74 $X2=4.685 $Y2=0.85
cc_379 N_A_c_330_n N_CI_M1026_g 0.0075473f $X=5.13 $Y=2.295 $X2=4.685 $Y2=3.235
cc_380 N_A_c_331_n N_CI_M1026_g 0.0872519f $X=5.13 $Y=2.445 $X2=4.685 $Y2=3.235
cc_381 N_A_c_338_n N_CI_c_819_n 0.00549051f $X=2.35 $Y=1.74 $X2=1.325 $Y2=1.74
cc_382 N_A_c_340_n N_CI_c_820_n 0.00186852f $X=5.01 $Y=1.74 $X2=3.415 $Y2=2.11
cc_383 N_A_c_330_n N_CI_c_821_n 0.0213433f $X=5.13 $Y=2.295 $X2=4.745 $Y2=1.92
cc_384 N_A_c_335_n N_CI_c_821_n 3.03194e-19 $X=5.155 $Y=1.74 $X2=4.745 $Y2=1.92
cc_385 N_A_c_340_n N_CI_c_821_n 0.00289458f $X=5.01 $Y=1.74 $X2=4.745 $Y2=1.92
cc_386 N_A_c_342_n N_CI_c_821_n 4.65422e-19 $X=5.155 $Y=1.74 $X2=4.745 $Y2=1.92
cc_387 N_A_c_332_n N_CI_c_822_n 0.00245253f $X=0.485 $Y=1.74 $X2=1.325 $Y2=1.74
cc_388 N_A_c_338_n N_CI_c_822_n 0.0182763f $X=2.35 $Y=1.74 $X2=1.325 $Y2=1.74
cc_389 N_A_c_339_n N_CI_c_822_n 0.00173513f $X=0.63 $Y=1.74 $X2=1.325 $Y2=1.74
cc_390 N_A_c_340_n N_CI_c_823_n 0.00421142f $X=5.01 $Y=1.74 $X2=3.415 $Y2=2.11
cc_391 N_A_c_330_n N_CI_c_824_n 0.00303989f $X=5.13 $Y=2.295 $X2=4.745 $Y2=1.92
cc_392 N_A_c_335_n N_CI_c_824_n 0.00330605f $X=5.155 $Y=1.74 $X2=4.745 $Y2=1.92
cc_393 N_A_c_340_n N_CI_c_824_n 0.00807394f $X=5.01 $Y=1.74 $X2=4.745 $Y2=1.92
cc_394 N_A_c_342_n N_CI_c_824_n 0.00133759f $X=5.155 $Y=1.74 $X2=4.745 $Y2=1.92
cc_395 N_A_c_313_n N_CI_c_825_n 0.00376374f $X=2.2 $Y=2.405 $X2=3.25 $Y2=2.11
cc_396 N_A_c_315_n N_CI_c_825_n 0.00603893f $X=2.435 $Y=2.33 $X2=3.25 $Y2=2.11
cc_397 N_A_c_323_n N_CI_c_825_n 9.34899e-19 $X=2.555 $Y=2.405 $X2=3.25 $Y2=2.11
cc_398 N_A_c_336_n N_CI_c_825_n 0.00331391f $X=2.495 $Y=1.65 $X2=3.25 $Y2=2.11
cc_399 N_A_c_338_n N_CI_c_825_n 0.0704728f $X=2.35 $Y=1.74 $X2=3.25 $Y2=2.11
cc_400 N_A_c_340_n N_CI_c_825_n 0.0503961f $X=5.01 $Y=1.74 $X2=3.25 $Y2=2.11
cc_401 N_A_c_341_n N_CI_c_825_n 0.026793f $X=2.64 $Y=1.74 $X2=3.25 $Y2=2.11
cc_402 N_A_c_338_n N_CI_c_826_n 0.0262115f $X=2.35 $Y=1.74 $X2=1.48 $Y2=2.11
cc_403 N_A_c_340_n N_CI_c_827_n 0.0822815f $X=5.01 $Y=1.74 $X2=4.6 $Y2=2.11
cc_404 N_A_c_340_n N_CI_c_828_n 0.0308225f $X=5.01 $Y=1.74 $X2=3.585 $Y2=2.11
cc_405 N_A_c_330_n N_CI_c_829_n 0.00414468f $X=5.13 $Y=2.295 $X2=4.745 $Y2=2.11
cc_406 N_A_c_340_n N_CI_c_829_n 0.0251723f $X=5.01 $Y=1.74 $X2=4.745 $Y2=2.11
cc_407 N_A_c_340_n N_CON_M1005_g 0.0015506f $X=5.01 $Y=1.74 $X2=3.845 $Y2=3.235
cc_408 N_A_c_340_n N_CON_c_992_n 0.00199858f $X=5.01 $Y=1.74 $X2=3.845 $Y2=1.455
cc_409 N_A_c_311_n N_CON_c_997_n 6.2115e-19 $X=2.2 $Y=1.28 $X2=1.665 $Y2=1.37
cc_410 N_A_c_313_n N_CON_c_997_n 2.54894e-19 $X=2.2 $Y=2.405 $X2=1.665 $Y2=1.37
cc_411 N_A_c_314_n N_CON_c_997_n 8.87736e-19 $X=2.495 $Y=1.65 $X2=1.665 $Y2=1.37
cc_412 N_A_c_322_n N_CON_c_997_n 2.73498e-19 $X=2.495 $Y=1.815 $X2=1.665
+ $Y2=1.37
cc_413 N_A_c_336_n N_CON_c_997_n 0.00419634f $X=2.495 $Y=1.65 $X2=1.665 $Y2=1.37
cc_414 N_A_c_338_n N_CON_c_997_n 0.0131226f $X=2.35 $Y=1.74 $X2=1.665 $Y2=1.37
cc_415 N_A_c_305_n N_CON_c_999_n 0.00108488f $X=2.125 $Y=1.205 $X2=1.665 $Y2=1.2
cc_416 N_A_c_338_n N_CON_c_999_n 0.0024397f $X=2.35 $Y=1.74 $X2=1.665 $Y2=1.2
cc_417 N_A_c_347_n N_CON_c_1026_n 9.14995e-19 $X=2.125 $Y=2.48 $X2=1.665
+ $Y2=2.637
cc_418 N_A_c_340_n N_CON_c_1000_n 0.00387001f $X=5.01 $Y=1.74 $X2=3.845
+ $Y2=1.455
cc_419 N_A_c_309_n N_CON_c_1003_n 0.00539432f $X=2.36 $Y=1.28 $X2=3.855 $Y2=1.37
cc_420 N_A_c_311_n N_CON_c_1003_n 0.00787523f $X=2.2 $Y=1.28 $X2=3.855 $Y2=1.37
cc_421 N_A_c_314_n N_CON_c_1003_n 0.00341866f $X=2.495 $Y=1.65 $X2=3.855
+ $Y2=1.37
cc_422 N_A_c_321_n N_CON_c_1003_n 0.0105901f $X=2.495 $Y=1.28 $X2=3.855 $Y2=1.37
cc_423 N_A_c_336_n N_CON_c_1003_n 0.00717801f $X=2.495 $Y=1.65 $X2=3.855
+ $Y2=1.37
cc_424 N_A_c_338_n N_CON_c_1003_n 0.0459849f $X=2.35 $Y=1.74 $X2=3.855 $Y2=1.37
cc_425 N_A_c_340_n N_CON_c_1003_n 0.101275f $X=5.01 $Y=1.74 $X2=3.855 $Y2=1.37
cc_426 N_A_c_341_n N_CON_c_1003_n 0.0252711f $X=2.64 $Y=1.74 $X2=3.855 $Y2=1.37
cc_427 N_A_c_338_n N_CON_c_1005_n 0.0252795f $X=2.35 $Y=1.74 $X2=1.81 $Y2=1.37
cc_428 N_A_c_324_n N_CON_c_1006_n 0.009249f $X=5.155 $Y=1.4 $X2=5.995 $Y2=1.37
cc_429 N_A_c_333_n N_CON_c_1006_n 0.0198918f $X=5.155 $Y=1.485 $X2=5.995
+ $Y2=1.37
cc_430 N_A_c_340_n N_CON_c_1006_n 0.0756037f $X=5.01 $Y=1.74 $X2=5.995 $Y2=1.37
cc_431 N_A_c_342_n N_CON_c_1006_n 0.0247185f $X=5.155 $Y=1.74 $X2=5.995 $Y2=1.37
cc_432 N_A_c_340_n N_CON_c_1008_n 0.0217763f $X=5.01 $Y=1.74 $X2=4.1 $Y2=1.37
cc_433 N_A_c_324_n N_A_784_115#_M1018_g 0.0201282f $X=5.155 $Y=1.4 $X2=5.585
+ $Y2=0.85
cc_434 N_A_c_326_n N_A_784_115#_M1018_g 0.020327f $X=5.155 $Y=1.235 $X2=5.585
+ $Y2=0.85
cc_435 N_A_c_330_n N_A_784_115#_M1018_g 0.0249853f $X=5.13 $Y=2.295 $X2=5.585
+ $Y2=0.85
cc_436 N_A_c_333_n N_A_784_115#_M1018_g 0.00106683f $X=5.155 $Y=1.485 $X2=5.585
+ $Y2=0.85
cc_437 N_A_c_335_n N_A_784_115#_M1018_g 0.00146812f $X=5.155 $Y=1.74 $X2=5.585
+ $Y2=0.85
cc_438 N_A_c_342_n N_A_784_115#_M1018_g 0.00409904f $X=5.155 $Y=1.74 $X2=5.585
+ $Y2=0.85
cc_439 N_A_M1021_g N_A_784_115#_M1007_g 0.0423117f $X=5.095 $Y=3.235 $X2=5.585
+ $Y2=3.235
cc_440 N_A_c_330_n N_A_784_115#_c_1161_n 0.0197344f $X=5.13 $Y=2.295 $X2=5.585
+ $Y2=2.275
cc_441 N_A_c_335_n N_A_784_115#_c_1163_n 6.53915e-19 $X=5.155 $Y=1.74 $X2=4.225
+ $Y2=1.795
cc_442 N_A_c_340_n N_A_784_115#_c_1163_n 0.015473f $X=5.01 $Y=1.74 $X2=4.225
+ $Y2=1.795
cc_443 N_A_c_340_n N_A_784_115#_c_1164_n 0.00946022f $X=5.01 $Y=1.74 $X2=3.93
+ $Y2=1.795
cc_444 N_A_M1021_g N_A_784_115#_c_1181_n 0.0193311f $X=5.095 $Y=3.235 $X2=5.33
+ $Y2=2.855
cc_445 N_A_c_331_n N_A_784_115#_c_1181_n 0.0016251f $X=5.13 $Y=2.445 $X2=5.33
+ $Y2=2.855
cc_446 N_A_c_333_n N_A_784_115#_c_1165_n 0.00351293f $X=5.155 $Y=1.485 $X2=4.31
+ $Y2=1.71
cc_447 N_A_c_335_n N_A_784_115#_c_1165_n 0.00489504f $X=5.155 $Y=1.74 $X2=4.31
+ $Y2=1.71
cc_448 N_A_c_340_n N_A_784_115#_c_1165_n 0.00650611f $X=5.01 $Y=1.74 $X2=4.31
+ $Y2=1.71
cc_449 N_A_c_342_n N_A_784_115#_c_1165_n 6.49234e-19 $X=5.155 $Y=1.74 $X2=4.31
+ $Y2=1.71
cc_450 N_A_M1021_g N_A_784_115#_c_1183_n 0.00698879f $X=5.095 $Y=3.235 $X2=5.415
+ $Y2=2.77
cc_451 N_A_c_330_n N_A_784_115#_c_1169_n 0.00651436f $X=5.13 $Y=2.295 $X2=5.415
+ $Y2=2.275
cc_452 N_A_M1000_g N_A_27_521#_c_1288_n 0.0169496f $X=0.475 $Y=3.235 $X2=1.035
+ $Y2=2.98
cc_453 N_A_c_333_n N_S_c_1317_n 0.00568068f $X=5.155 $Y=1.485 $X2=5.8 $Y2=0.755
cc_454 N_A_c_335_n N_S_c_1317_n 0.00516363f $X=5.155 $Y=1.74 $X2=5.8 $Y2=0.755
cc_455 N_A_c_342_n N_S_c_1317_n 7.50607e-19 $X=5.155 $Y=1.74 $X2=5.8 $Y2=0.755
cc_456 N_A_c_342_n N_S_c_1321_n 0.00103006f $X=5.155 $Y=1.74 $X2=5.925 $Y2=2.685
cc_457 N_A_c_335_n N_S_c_1322_n 0.00335037f $X=5.155 $Y=1.74 $X2=5.925 $Y2=1.74
cc_458 N_A_c_342_n N_S_c_1322_n 0.00491314f $X=5.155 $Y=1.74 $X2=5.925 $Y2=1.74
cc_459 N_A_M1013_g N_A_27_115#_c_1387_n 0.0165142f $X=0.475 $Y=0.85 $X2=1.035
+ $Y2=1.16
cc_460 N_A_c_320_n N_A_27_115#_c_1387_n 0.00247554f $X=0.485 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_461 N_A_c_332_n N_A_27_115#_c_1387_n 0.00675159f $X=0.485 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_462 N_A_c_338_n N_A_27_115#_c_1387_n 0.0206117f $X=2.35 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_463 N_A_c_339_n N_A_27_115#_c_1387_n 0.00572534f $X=0.63 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_464 N_A_M1013_g N_A_27_115#_c_1394_n 0.00157308f $X=0.475 $Y=0.85 $X2=0.262
+ $Y2=1.16
cc_465 N_A_c_332_n N_A_27_115#_c_1394_n 0.00118386f $X=0.485 $Y=1.74 $X2=0.262
+ $Y2=1.16
cc_466 N_A_c_339_n N_A_27_115#_c_1394_n 2.32641e-19 $X=0.63 $Y=1.74 $X2=0.262
+ $Y2=1.16
cc_467 N_A_c_316_n N_A_526_115#_c_1410_n 3.74023e-19 $X=2.555 $Y=1.205 $X2=2.77
+ $Y2=0.755
cc_468 N_A_c_316_n N_A_526_115#_c_1418_n 0.00274649f $X=2.555 $Y=1.205 $X2=2.855
+ $Y2=1.115
cc_469 N_B_M1001_g N_CI_M1003_g 0.0343075f $X=0.905 $Y=0.85 $X2=1.335 $Y2=0.85
cc_470 N_B_M1025_g N_CI_M1003_g 0.0326327f $X=1.765 $Y=0.85 $X2=1.335 $Y2=0.85
cc_471 N_B_M1001_g N_CI_M1020_g 0.00863862f $X=0.905 $Y=0.85 $X2=1.335 $Y2=3.235
cc_472 N_B_M1019_g N_CI_M1020_g 0.0365393f $X=0.905 $Y=3.235 $X2=1.335 $Y2=3.235
cc_473 N_B_c_551_n N_CI_M1020_g 0.0185048f $X=0.895 $Y=2.28 $X2=1.335 $Y2=3.235
cc_474 N_B_c_552_n N_CI_M1020_g 0.0575121f $X=2.015 $Y=1.95 $X2=1.335 $Y2=3.235
cc_475 N_B_c_555_n N_CI_M1020_g 0.00161155f $X=0.895 $Y=2.28 $X2=1.335 $Y2=3.235
cc_476 N_B_c_561_n N_CI_M1020_g 0.0101401f $X=2.16 $Y=2.48 $X2=1.335 $Y2=3.235
cc_477 N_B_M1024_g N_CI_M1014_g 0.0336019f $X=2.985 $Y=0.85 $X2=3.415 $Y2=0.85
cc_478 N_B_M1011_g N_CI_M1014_g 0.00538306f $X=2.985 $Y=3.235 $X2=3.415 $Y2=0.85
cc_479 N_B_c_553_n N_CI_M1014_g 0.0197963f $X=2.975 $Y=1.655 $X2=3.415 $Y2=0.85
cc_480 N_B_c_557_n N_CI_M1014_g 0.00316322f $X=2.975 $Y=1.655 $X2=3.415 $Y2=0.85
cc_481 N_B_M1011_g N_CI_M1002_g 0.0624488f $X=2.985 $Y=3.235 $X2=3.415 $Y2=3.235
cc_482 N_B_c_557_n N_CI_M1002_g 0.00247376f $X=2.975 $Y=1.655 $X2=3.415
+ $Y2=3.235
cc_483 N_B_c_564_n N_CI_M1002_g 0.00637636f $X=4.12 $Y=2.48 $X2=3.415 $Y2=3.235
cc_484 N_B_c_565_n N_CI_M1002_g 8.82664e-19 $X=3.12 $Y=2.48 $X2=3.415 $Y2=3.235
cc_485 N_B_M1017_g N_CI_M1008_g 0.0755763f $X=4.275 $Y=0.85 $X2=4.685 $Y2=0.85
cc_486 N_B_M1006_g N_CI_M1026_g 0.0855548f $X=4.275 $Y=3.235 $X2=4.685 $Y2=3.235
cc_487 N_B_c_558_n N_CI_M1026_g 0.00297508f $X=4.265 $Y=2.48 $X2=4.685 $Y2=3.235
cc_488 N_B_c_566_n N_CI_M1026_g 0.0042599f $X=4.265 $Y=2.48 $X2=4.685 $Y2=3.235
cc_489 N_B_M1001_g N_CI_c_819_n 0.0219935f $X=0.905 $Y=0.85 $X2=1.325 $Y2=1.74
cc_490 N_B_M1025_g N_CI_c_819_n 0.0189858f $X=1.765 $Y=0.85 $X2=1.325 $Y2=1.74
cc_491 N_B_M1011_g N_CI_c_820_n 0.0205508f $X=2.985 $Y=3.235 $X2=3.415 $Y2=2.11
cc_492 N_B_c_557_n N_CI_c_820_n 0.00139232f $X=2.975 $Y=1.655 $X2=3.415 $Y2=2.11
cc_493 N_B_c_564_n N_CI_c_820_n 0.00186852f $X=4.12 $Y=2.48 $X2=3.415 $Y2=2.11
cc_494 N_B_c_554_n N_CI_c_821_n 0.0218143f $X=4.265 $Y=2.135 $X2=4.745 $Y2=1.92
cc_495 N_B_c_560_n N_CI_c_821_n 0.0011908f $X=4.265 $Y=2.135 $X2=4.745 $Y2=1.92
cc_496 N_B_M1001_g N_CI_c_822_n 0.00509772f $X=0.905 $Y=0.85 $X2=1.325 $Y2=1.74
cc_497 N_B_M1025_g N_CI_c_822_n 7.83117e-19 $X=1.765 $Y=0.85 $X2=1.325 $Y2=1.74
cc_498 N_B_c_551_n N_CI_c_822_n 0.00125384f $X=0.895 $Y=2.28 $X2=1.325 $Y2=1.74
cc_499 N_B_c_561_n N_CI_c_822_n 0.00261972f $X=2.16 $Y=2.48 $X2=1.325 $Y2=1.74
cc_500 N_B_M1011_g N_CI_c_823_n 6.71807e-19 $X=2.985 $Y=3.235 $X2=3.415 $Y2=2.11
cc_501 N_B_c_557_n N_CI_c_823_n 0.0102939f $X=2.975 $Y=1.655 $X2=3.415 $Y2=2.11
cc_502 N_B_c_564_n N_CI_c_823_n 0.00421142f $X=4.12 $Y=2.48 $X2=3.415 $Y2=2.11
cc_503 N_B_M1017_g N_CI_c_824_n 7.00026e-19 $X=4.275 $Y=0.85 $X2=4.745 $Y2=1.92
cc_504 N_B_c_554_n N_CI_c_824_n 9.49552e-19 $X=4.265 $Y=2.135 $X2=4.745 $Y2=1.92
cc_505 N_B_c_560_n N_CI_c_824_n 0.00724517f $X=4.265 $Y=2.135 $X2=4.745 $Y2=1.92
cc_506 N_B_M1012_g N_CI_c_825_n 0.00170136f $X=1.765 $Y=3.235 $X2=3.25 $Y2=2.11
cc_507 N_B_M1011_g N_CI_c_825_n 8.61868e-19 $X=2.985 $Y=3.235 $X2=3.25 $Y2=2.11
cc_508 N_B_c_552_n N_CI_c_825_n 0.00364968f $X=2.015 $Y=1.95 $X2=3.25 $Y2=2.11
cc_509 N_B_c_553_n N_CI_c_825_n 5.37679e-19 $X=2.975 $Y=1.655 $X2=3.25 $Y2=2.11
cc_510 N_B_c_556_n N_CI_c_825_n 0.0153524f $X=2.015 $Y=1.95 $X2=3.25 $Y2=2.11
cc_511 N_B_c_585_n N_CI_c_825_n 0.00372007f $X=2.305 $Y=2.48 $X2=3.25 $Y2=2.11
cc_512 N_B_c_557_n N_CI_c_825_n 0.0157783f $X=2.975 $Y=1.655 $X2=3.25 $Y2=2.11
cc_513 N_B_c_561_n N_CI_c_825_n 0.0544374f $X=2.16 $Y=2.48 $X2=3.25 $Y2=2.11
cc_514 N_B_c_563_n N_CI_c_825_n 0.0321777f $X=2.83 $Y=2.48 $X2=3.25 $Y2=2.11
cc_515 N_B_c_593_n N_CI_c_825_n 0.0265493f $X=2.45 $Y=2.48 $X2=3.25 $Y2=2.11
cc_516 N_B_c_564_n N_CI_c_825_n 0.0110545f $X=4.12 $Y=2.48 $X2=3.25 $Y2=2.11
cc_517 N_B_c_565_n N_CI_c_825_n 0.0253568f $X=3.12 $Y=2.48 $X2=3.25 $Y2=2.11
cc_518 N_B_M1001_g N_CI_c_826_n 0.0021686f $X=0.905 $Y=0.85 $X2=1.48 $Y2=2.11
cc_519 N_B_c_551_n N_CI_c_826_n 0.00159754f $X=0.895 $Y=2.28 $X2=1.48 $Y2=2.11
cc_520 N_B_c_555_n N_CI_c_826_n 0.00109446f $X=0.895 $Y=2.28 $X2=1.48 $Y2=2.11
cc_521 N_B_c_561_n N_CI_c_826_n 0.0277565f $X=2.16 $Y=2.48 $X2=1.48 $Y2=2.11
cc_522 N_B_c_554_n N_CI_c_827_n 0.00149553f $X=4.265 $Y=2.135 $X2=4.6 $Y2=2.11
cc_523 N_B_c_560_n N_CI_c_827_n 0.0133678f $X=4.265 $Y=2.135 $X2=4.6 $Y2=2.11
cc_524 N_B_c_564_n N_CI_c_827_n 0.0439483f $X=4.12 $Y=2.48 $X2=4.6 $Y2=2.11
cc_525 N_B_c_566_n N_CI_c_827_n 0.0251333f $X=4.265 $Y=2.48 $X2=4.6 $Y2=2.11
cc_526 N_B_M1011_g N_CI_c_828_n 9.12723e-19 $X=2.985 $Y=3.235 $X2=3.585 $Y2=2.11
cc_527 N_B_c_557_n N_CI_c_828_n 0.00268964f $X=2.975 $Y=1.655 $X2=3.585 $Y2=2.11
cc_528 N_B_c_564_n N_CI_c_828_n 0.0308225f $X=4.12 $Y=2.48 $X2=3.585 $Y2=2.11
cc_529 N_B_c_554_n N_CI_c_829_n 5.16714e-19 $X=4.265 $Y=2.135 $X2=4.745 $Y2=2.11
cc_530 N_B_c_560_n N_CI_c_829_n 0.00130045f $X=4.265 $Y=2.135 $X2=4.745 $Y2=2.11
cc_531 N_B_M1017_g N_CON_M1015_g 0.0230684f $X=4.275 $Y=0.85 $X2=3.845 $Y2=0.85
cc_532 N_B_M1017_g N_CON_M1005_g 0.0156819f $X=4.275 $Y=0.85 $X2=3.845 $Y2=3.235
cc_533 N_B_M1006_g N_CON_M1005_g 0.0421867f $X=4.275 $Y=3.235 $X2=3.845
+ $Y2=3.235
cc_534 N_B_c_554_n N_CON_M1005_g 0.0209816f $X=4.265 $Y=2.135 $X2=3.845
+ $Y2=3.235
cc_535 N_B_c_558_n N_CON_M1005_g 8.3458e-19 $X=4.265 $Y=2.48 $X2=3.845 $Y2=3.235
cc_536 N_B_c_560_n N_CON_M1005_g 4.50389e-19 $X=4.265 $Y=2.135 $X2=3.845
+ $Y2=3.235
cc_537 N_B_M1017_g N_CON_c_992_n 0.0199638f $X=4.275 $Y=0.85 $X2=3.845 $Y2=1.455
cc_538 N_B_M1025_g N_CON_c_994_n 7.48782e-19 $X=1.765 $Y=0.85 $X2=1.55 $Y2=0.755
cc_539 N_B_c_561_n N_CON_c_1020_n 8.38683e-19 $X=2.16 $Y=2.48 $X2=1.55 $Y2=3.295
cc_540 N_B_M1025_g N_CON_c_997_n 0.0137122f $X=1.765 $Y=0.85 $X2=1.665 $Y2=1.37
cc_541 N_B_M1012_g N_CON_c_997_n 0.00745479f $X=1.765 $Y=3.235 $X2=1.665
+ $Y2=1.37
cc_542 N_B_c_552_n N_CON_c_997_n 0.00755272f $X=2.015 $Y=1.95 $X2=1.665 $Y2=1.37
cc_543 N_B_c_555_n N_CON_c_997_n 0.00565241f $X=0.895 $Y=2.28 $X2=1.665 $Y2=1.37
cc_544 N_B_c_556_n N_CON_c_997_n 0.039273f $X=2.015 $Y=1.95 $X2=1.665 $Y2=1.37
cc_545 N_B_c_584_n N_CON_c_997_n 0.0097817f $X=2.1 $Y=2.48 $X2=1.665 $Y2=1.37
cc_546 N_B_c_561_n N_CON_c_997_n 0.0120419f $X=2.16 $Y=2.48 $X2=1.665 $Y2=1.37
cc_547 N_B_M1025_g N_CON_c_999_n 0.00764736f $X=1.765 $Y=0.85 $X2=1.665 $Y2=1.2
cc_548 N_B_M1012_g N_CON_c_1026_n 0.0075031f $X=1.765 $Y=3.235 $X2=1.665
+ $Y2=2.637
cc_549 N_B_c_584_n N_CON_c_1026_n 0.00124924f $X=2.1 $Y=2.48 $X2=1.665 $Y2=2.637
cc_550 N_B_c_561_n N_CON_c_1026_n 0.011664f $X=2.16 $Y=2.48 $X2=1.665 $Y2=2.637
cc_551 N_B_c_593_n N_CON_c_1026_n 9.96079e-19 $X=2.45 $Y=2.48 $X2=1.665
+ $Y2=2.637
cc_552 N_B_M1017_g N_CON_c_1000_n 0.00117535f $X=4.275 $Y=0.85 $X2=3.845
+ $Y2=1.455
cc_553 N_B_c_557_n N_CON_c_1000_n 0.00143014f $X=2.975 $Y=1.655 $X2=3.845
+ $Y2=1.455
cc_554 N_B_M1025_g N_CON_c_1003_n 0.00339936f $X=1.765 $Y=0.85 $X2=3.855
+ $Y2=1.37
cc_555 N_B_M1024_g N_CON_c_1003_n 0.00540482f $X=2.985 $Y=0.85 $X2=3.855
+ $Y2=1.37
cc_556 N_B_c_552_n N_CON_c_1003_n 5.24163e-19 $X=2.015 $Y=1.95 $X2=3.855
+ $Y2=1.37
cc_557 N_B_c_553_n N_CON_c_1003_n 0.00169614f $X=2.975 $Y=1.655 $X2=3.855
+ $Y2=1.37
cc_558 N_B_c_556_n N_CON_c_1003_n 0.00249638f $X=2.015 $Y=1.95 $X2=3.855
+ $Y2=1.37
cc_559 N_B_c_557_n N_CON_c_1003_n 0.00185056f $X=2.975 $Y=1.655 $X2=3.855
+ $Y2=1.37
cc_560 N_B_M1025_g N_CON_c_1005_n 0.00419948f $X=1.765 $Y=0.85 $X2=1.81 $Y2=1.37
cc_561 N_B_M1017_g N_CON_c_1006_n 0.00131714f $X=4.275 $Y=0.85 $X2=5.995
+ $Y2=1.37
cc_562 N_B_M1017_g N_CON_c_1008_n 9.0633e-19 $X=4.275 $Y=0.85 $X2=4.1 $Y2=1.37
cc_563 N_B_M1017_g N_A_784_115#_c_1162_n 0.00163203f $X=4.275 $Y=0.85 $X2=3.845
+ $Y2=2.55
cc_564 N_B_M1006_g N_A_784_115#_c_1162_n 7.03843e-19 $X=4.275 $Y=3.235 $X2=3.845
+ $Y2=2.55
cc_565 N_B_c_554_n N_A_784_115#_c_1162_n 0.00230204f $X=4.265 $Y=2.135 $X2=3.845
+ $Y2=2.55
cc_566 N_B_c_558_n N_A_784_115#_c_1162_n 0.016716f $X=4.265 $Y=2.48 $X2=3.845
+ $Y2=2.55
cc_567 N_B_c_560_n N_A_784_115#_c_1162_n 0.0122483f $X=4.265 $Y=2.135 $X2=3.845
+ $Y2=2.55
cc_568 N_B_c_564_n N_A_784_115#_c_1162_n 0.0129177f $X=4.12 $Y=2.48 $X2=3.845
+ $Y2=2.55
cc_569 N_B_c_566_n N_A_784_115#_c_1162_n 0.00102158f $X=4.265 $Y=2.48 $X2=3.845
+ $Y2=2.55
cc_570 N_B_M1017_g N_A_784_115#_c_1163_n 0.00761698f $X=4.275 $Y=0.85 $X2=4.225
+ $Y2=1.795
cc_571 N_B_c_554_n N_A_784_115#_c_1163_n 0.00287887f $X=4.265 $Y=2.135 $X2=4.225
+ $Y2=1.795
cc_572 N_B_c_560_n N_A_784_115#_c_1163_n 0.0193935f $X=4.265 $Y=2.135 $X2=4.225
+ $Y2=1.795
cc_573 N_B_M1006_g N_A_784_115#_c_1177_n 0.0013092f $X=4.275 $Y=3.235 $X2=4.06
+ $Y2=2.94
cc_574 N_B_c_554_n N_A_784_115#_c_1177_n 2.86796e-19 $X=4.265 $Y=2.135 $X2=4.06
+ $Y2=2.94
cc_575 N_B_c_558_n N_A_784_115#_c_1177_n 7.43237e-19 $X=4.265 $Y=2.48 $X2=4.06
+ $Y2=2.94
cc_576 N_B_c_560_n N_A_784_115#_c_1177_n 5.96301e-19 $X=4.265 $Y=2.135 $X2=4.06
+ $Y2=2.94
cc_577 N_B_c_564_n N_A_784_115#_c_1177_n 0.0184847f $X=4.12 $Y=2.48 $X2=4.06
+ $Y2=2.94
cc_578 N_B_c_566_n N_A_784_115#_c_1177_n 0.00255596f $X=4.265 $Y=2.48 $X2=4.06
+ $Y2=2.94
cc_579 N_B_M1006_g N_A_784_115#_c_1181_n 0.0149079f $X=4.275 $Y=3.235 $X2=5.33
+ $Y2=2.855
cc_580 N_B_c_558_n N_A_784_115#_c_1181_n 0.00784247f $X=4.265 $Y=2.48 $X2=5.33
+ $Y2=2.855
cc_581 N_B_c_560_n N_A_784_115#_c_1181_n 8.31144e-19 $X=4.265 $Y=2.135 $X2=5.33
+ $Y2=2.855
cc_582 N_B_c_566_n N_A_784_115#_c_1181_n 0.00727276f $X=4.265 $Y=2.48 $X2=5.33
+ $Y2=2.855
cc_583 N_B_M1017_g N_A_784_115#_c_1165_n 0.0187094f $X=4.275 $Y=0.85 $X2=4.31
+ $Y2=1.71
cc_584 N_B_M1017_g N_A_784_115#_c_1166_n 0.006753f $X=4.275 $Y=0.85 $X2=4.06
+ $Y2=0.74
cc_585 N_B_M1019_g N_A_27_521#_c_1288_n 0.0161147f $X=0.905 $Y=3.235 $X2=1.035
+ $Y2=2.98
cc_586 N_B_c_551_n N_A_27_521#_c_1288_n 6.80629e-19 $X=0.895 $Y=2.28 $X2=1.035
+ $Y2=2.98
cc_587 N_B_c_555_n N_A_27_521#_c_1288_n 0.00528048f $X=0.895 $Y=2.28 $X2=1.035
+ $Y2=2.98
cc_588 N_B_c_559_n N_A_27_521#_c_1288_n 0.00451483f $X=0.485 $Y=2.28 $X2=1.035
+ $Y2=2.98
cc_589 N_B_c_561_n N_A_27_521#_c_1288_n 0.0169669f $X=2.16 $Y=2.48 $X2=1.035
+ $Y2=2.98
cc_590 N_B_c_562_n N_A_27_521#_c_1288_n 0.00770039f $X=0.63 $Y=2.48 $X2=1.035
+ $Y2=2.98
cc_591 N_B_M1011_g N_A_526_521#_c_1300_n 0.01474f $X=2.985 $Y=3.235 $X2=3.545
+ $Y2=3.23
cc_592 N_B_c_557_n N_A_526_521#_c_1300_n 0.00208738f $X=2.975 $Y=1.655 $X2=3.545
+ $Y2=3.23
cc_593 N_B_c_564_n N_A_526_521#_c_1300_n 0.018439f $X=4.12 $Y=2.48 $X2=3.545
+ $Y2=3.23
cc_594 N_B_c_565_n N_A_526_521#_c_1300_n 0.00615328f $X=3.12 $Y=2.48 $X2=3.545
+ $Y2=3.23
cc_595 N_B_c_563_n N_A_526_521#_c_1305_n 0.00560026f $X=2.83 $Y=2.48 $X2=2.77
+ $Y2=3.295
cc_596 N_B_c_565_n N_A_526_521#_c_1305_n 9.8393e-19 $X=3.12 $Y=2.48 $X2=2.77
+ $Y2=3.295
cc_597 N_B_M1001_g N_A_27_115#_c_1387_n 0.0153084f $X=0.905 $Y=0.85 $X2=1.035
+ $Y2=1.16
cc_598 N_B_M1001_g N_A_27_115#_c_1390_n 5.63412e-19 $X=0.905 $Y=0.85 $X2=1.12
+ $Y2=0.755
cc_599 N_B_M1024_g N_A_526_115#_c_1410_n 3.74023e-19 $X=2.985 $Y=0.85 $X2=2.77
+ $Y2=0.755
cc_600 N_B_M1024_g N_A_526_115#_c_1415_n 0.0141303f $X=2.985 $Y=0.85 $X2=3.545
+ $Y2=1.115
cc_601 N_B_c_553_n N_A_526_115#_c_1415_n 0.00294604f $X=2.975 $Y=1.655 $X2=3.545
+ $Y2=1.115
cc_602 N_B_c_557_n N_A_526_115#_c_1415_n 0.00496839f $X=2.975 $Y=1.655 $X2=3.545
+ $Y2=1.115
cc_603 N_B_c_553_n N_A_526_115#_c_1418_n 5.77386e-19 $X=2.975 $Y=1.655 $X2=2.855
+ $Y2=1.115
cc_604 N_CI_M1014_g N_CON_M1015_g 0.0216753f $X=3.415 $Y=0.85 $X2=3.845 $Y2=0.85
cc_605 N_CI_M1014_g N_CON_M1005_g 0.0149568f $X=3.415 $Y=0.85 $X2=3.845
+ $Y2=3.235
cc_606 N_CI_M1002_g N_CON_M1005_g 0.0569699f $X=3.415 $Y=3.235 $X2=3.845
+ $Y2=3.235
cc_607 N_CI_c_820_n N_CON_M1005_g 0.0200144f $X=3.415 $Y=2.11 $X2=3.845
+ $Y2=3.235
cc_608 N_CI_c_823_n N_CON_M1005_g 4.36547e-19 $X=3.415 $Y=2.11 $X2=3.845
+ $Y2=3.235
cc_609 N_CI_M1014_g N_CON_c_992_n 0.0205382f $X=3.415 $Y=0.85 $X2=3.845
+ $Y2=1.455
cc_610 N_CI_M1003_g N_CON_c_994_n 7.31757e-19 $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=0.755
cc_611 N_CI_M1003_g N_CON_c_997_n 0.00525468f $X=1.335 $Y=0.85 $X2=1.665
+ $Y2=1.37
cc_612 N_CI_M1020_g N_CON_c_997_n 0.00601328f $X=1.335 $Y=3.235 $X2=1.665
+ $Y2=1.37
cc_613 N_CI_c_819_n N_CON_c_997_n 0.00175448f $X=1.325 $Y=1.74 $X2=1.665
+ $Y2=1.37
cc_614 N_CI_c_822_n N_CON_c_997_n 0.0427337f $X=1.325 $Y=1.74 $X2=1.665 $Y2=1.37
cc_615 N_CI_c_825_n N_CON_c_997_n 0.011693f $X=3.25 $Y=2.11 $X2=1.665 $Y2=1.37
cc_616 N_CI_c_826_n N_CON_c_997_n 0.00204819f $X=1.48 $Y=2.11 $X2=1.665 $Y2=1.37
cc_617 N_CI_M1003_g N_CON_c_999_n 0.00211843f $X=1.335 $Y=0.85 $X2=1.665 $Y2=1.2
cc_618 N_CI_M1020_g N_CON_c_1026_n 0.0019658f $X=1.335 $Y=3.235 $X2=1.665
+ $Y2=2.637
cc_619 N_CI_c_825_n N_CON_c_1026_n 6.01856e-19 $X=3.25 $Y=2.11 $X2=1.665
+ $Y2=2.637
cc_620 N_CI_M1014_g N_CON_c_1000_n 0.00334783f $X=3.415 $Y=0.85 $X2=3.845
+ $Y2=1.455
cc_621 N_CI_M1014_g N_CON_c_1003_n 0.0055726f $X=3.415 $Y=0.85 $X2=3.855
+ $Y2=1.37
cc_622 N_CI_M1003_g N_CON_c_1005_n 0.00394781f $X=1.335 $Y=0.85 $X2=1.81
+ $Y2=1.37
cc_623 N_CI_M1008_g N_CON_c_1006_n 0.010613f $X=4.685 $Y=0.85 $X2=5.995 $Y2=1.37
cc_624 N_CI_c_821_n N_CON_c_1006_n 2.41418e-19 $X=4.745 $Y=1.92 $X2=5.995
+ $Y2=1.37
cc_625 N_CI_c_824_n N_CON_c_1006_n 0.0023884f $X=4.745 $Y=1.92 $X2=5.995
+ $Y2=1.37
cc_626 N_CI_M1014_g N_A_784_115#_c_1162_n 0.0011736f $X=3.415 $Y=0.85 $X2=3.845
+ $Y2=2.55
cc_627 N_CI_M1002_g N_A_784_115#_c_1162_n 0.00427742f $X=3.415 $Y=3.235
+ $X2=3.845 $Y2=2.55
cc_628 N_CI_c_820_n N_A_784_115#_c_1162_n 0.00347943f $X=3.415 $Y=2.11 $X2=3.845
+ $Y2=2.55
cc_629 N_CI_c_823_n N_A_784_115#_c_1162_n 0.0113765f $X=3.415 $Y=2.11 $X2=3.845
+ $Y2=2.55
cc_630 N_CI_c_827_n N_A_784_115#_c_1162_n 0.0124958f $X=4.6 $Y=2.11 $X2=3.845
+ $Y2=2.55
cc_631 N_CI_c_828_n N_A_784_115#_c_1162_n 0.00295734f $X=3.585 $Y=2.11 $X2=3.845
+ $Y2=2.55
cc_632 N_CI_M1008_g N_A_784_115#_c_1163_n 0.00112503f $X=4.685 $Y=0.85 $X2=4.225
+ $Y2=1.795
cc_633 N_CI_c_824_n N_A_784_115#_c_1163_n 0.00608653f $X=4.745 $Y=1.92 $X2=4.225
+ $Y2=1.795
cc_634 N_CI_c_827_n N_A_784_115#_c_1163_n 0.0064487f $X=4.6 $Y=2.11 $X2=4.225
+ $Y2=1.795
cc_635 N_CI_M1014_g N_A_784_115#_c_1164_n 0.00310209f $X=3.415 $Y=0.85 $X2=3.93
+ $Y2=1.795
cc_636 N_CI_M1002_g N_A_784_115#_c_1177_n 0.00185418f $X=3.415 $Y=3.235 $X2=4.06
+ $Y2=2.94
cc_637 N_CI_M1026_g N_A_784_115#_c_1181_n 0.0164402f $X=4.685 $Y=3.235 $X2=5.33
+ $Y2=2.855
cc_638 N_CI_c_821_n N_A_784_115#_c_1181_n 9.74133e-19 $X=4.745 $Y=1.92 $X2=5.33
+ $Y2=2.855
cc_639 N_CI_c_824_n N_A_784_115#_c_1181_n 0.00204032f $X=4.745 $Y=1.92 $X2=5.33
+ $Y2=2.855
cc_640 N_CI_c_827_n N_A_784_115#_c_1181_n 0.00554537f $X=4.6 $Y=2.11 $X2=5.33
+ $Y2=2.855
cc_641 N_CI_c_829_n N_A_784_115#_c_1181_n 0.00692907f $X=4.745 $Y=2.11 $X2=5.33
+ $Y2=2.855
cc_642 N_CI_M1008_g N_A_784_115#_c_1165_n 0.0072079f $X=4.685 $Y=0.85 $X2=4.31
+ $Y2=1.71
cc_643 N_CI_c_824_n N_A_784_115#_c_1169_n 0.00112894f $X=4.745 $Y=1.92 $X2=5.415
+ $Y2=2.275
cc_644 N_CI_c_829_n N_A_784_115#_c_1169_n 0.00318599f $X=4.745 $Y=2.11 $X2=5.415
+ $Y2=2.275
cc_645 N_CI_M1002_g N_A_526_521#_c_1300_n 0.0160555f $X=3.415 $Y=3.235 $X2=3.545
+ $Y2=3.23
cc_646 N_CI_M1003_g N_A_27_115#_c_1387_n 0.00138916f $X=1.335 $Y=0.85 $X2=1.035
+ $Y2=1.16
cc_647 N_CI_c_819_n N_A_27_115#_c_1387_n 5.57939e-19 $X=1.325 $Y=1.74 $X2=1.035
+ $Y2=1.16
cc_648 N_CI_M1003_g N_A_27_115#_c_1390_n 5.63412e-19 $X=1.335 $Y=0.85 $X2=1.12
+ $Y2=0.755
cc_649 N_CI_M1014_g N_A_526_115#_c_1415_n 0.0138152f $X=3.415 $Y=0.85 $X2=3.545
+ $Y2=1.115
cc_650 N_CI_M1014_g N_A_526_115#_c_1419_n 3.74023e-19 $X=3.415 $Y=0.85 $X2=3.63
+ $Y2=0.755
cc_651 N_CON_c_998_n N_A_784_115#_M1018_g 0.00118029f $X=6.41 $Y=2.26 $X2=5.585
+ $Y2=0.85
cc_652 N_CON_c_1006_n N_A_784_115#_M1018_g 0.0166629f $X=5.995 $Y=1.37 $X2=5.585
+ $Y2=0.85
cc_653 N_CON_c_993_n N_A_784_115#_c_1161_n 0.00451843f $X=6.41 $Y=2.26 $X2=5.585
+ $Y2=2.275
cc_654 N_CON_M1005_g N_A_784_115#_c_1162_n 0.0125625f $X=3.845 $Y=3.235
+ $X2=3.845 $Y2=2.55
cc_655 N_CON_c_992_n N_A_784_115#_c_1163_n 0.00120777f $X=3.845 $Y=1.455
+ $X2=4.225 $Y2=1.795
cc_656 N_CON_c_1000_n N_A_784_115#_c_1163_n 0.0081374f $X=3.845 $Y=1.455
+ $X2=4.225 $Y2=1.795
cc_657 N_CON_c_1006_n N_A_784_115#_c_1163_n 9.69195e-19 $X=5.995 $Y=1.37
+ $X2=4.225 $Y2=1.795
cc_658 N_CON_c_1008_n N_A_784_115#_c_1163_n 4.37195e-19 $X=4.1 $Y=1.37 $X2=4.225
+ $Y2=1.795
cc_659 N_CON_M1005_g N_A_784_115#_c_1164_n 0.00603753f $X=3.845 $Y=3.235
+ $X2=3.93 $Y2=1.795
cc_660 N_CON_c_992_n N_A_784_115#_c_1164_n 4.92662e-19 $X=3.845 $Y=1.455
+ $X2=3.93 $Y2=1.795
cc_661 N_CON_c_1000_n N_A_784_115#_c_1164_n 0.0104493f $X=3.845 $Y=1.455
+ $X2=3.93 $Y2=1.795
cc_662 N_CON_M1005_g N_A_784_115#_c_1177_n 0.0172636f $X=3.845 $Y=3.235 $X2=4.06
+ $Y2=2.94
cc_663 N_CON_M1015_g N_A_784_115#_c_1165_n 0.00139535f $X=3.845 $Y=0.85 $X2=4.31
+ $Y2=1.71
cc_664 N_CON_M1005_g N_A_784_115#_c_1165_n 6.92976e-19 $X=3.845 $Y=3.235
+ $X2=4.31 $Y2=1.71
cc_665 N_CON_c_992_n N_A_784_115#_c_1165_n 8.69455e-19 $X=3.845 $Y=1.455
+ $X2=4.31 $Y2=1.71
cc_666 N_CON_c_1000_n N_A_784_115#_c_1165_n 0.0176297f $X=3.845 $Y=1.455
+ $X2=4.31 $Y2=1.71
cc_667 N_CON_c_1006_n N_A_784_115#_c_1165_n 0.0201151f $X=5.995 $Y=1.37 $X2=4.31
+ $Y2=1.71
cc_668 N_CON_c_1008_n N_A_784_115#_c_1165_n 0.00225703f $X=4.1 $Y=1.37 $X2=4.31
+ $Y2=1.71
cc_669 N_CON_c_1000_n N_A_784_115#_c_1166_n 0.0027165f $X=3.845 $Y=1.455
+ $X2=4.06 $Y2=0.74
cc_670 N_CON_c_1006_n N_A_784_115#_c_1166_n 0.00481242f $X=5.995 $Y=1.37
+ $X2=4.06 $Y2=0.74
cc_671 N_CON_c_1008_n N_A_784_115#_c_1166_n 0.00414256f $X=4.1 $Y=1.37 $X2=4.06
+ $Y2=0.74
cc_672 N_CON_M1023_g N_S_c_1317_n 0.0102543f $X=6.535 $Y=0.85 $X2=5.8 $Y2=0.755
cc_673 N_CON_c_998_n N_S_c_1317_n 0.00716033f $X=6.41 $Y=2.26 $X2=5.8 $Y2=0.755
cc_674 N_CON_c_1001_n N_S_c_1317_n 0.0121035f $X=6.41 $Y=1.37 $X2=5.8 $Y2=0.755
cc_675 N_CON_c_1006_n N_S_c_1317_n 0.0196259f $X=5.995 $Y=1.37 $X2=5.8 $Y2=0.755
cc_676 CON N_S_c_1317_n 0.00260317f $X=6.14 $Y=1.37 $X2=5.8 $Y2=0.755
cc_677 N_CON_M1023_g N_S_c_1321_n 0.00130367f $X=6.535 $Y=0.85 $X2=5.925
+ $Y2=2.685
cc_678 N_CON_M1010_g N_S_c_1321_n 0.00437761f $X=6.535 $Y=3.235 $X2=5.925
+ $Y2=2.685
cc_679 N_CON_c_993_n N_S_c_1321_n 0.00305399f $X=6.41 $Y=2.26 $X2=5.925
+ $Y2=2.685
cc_680 N_CON_c_998_n N_S_c_1321_n 0.0278588f $X=6.41 $Y=2.26 $X2=5.925 $Y2=2.685
cc_681 N_CON_M1023_g N_S_c_1322_n 8.65886e-19 $X=6.535 $Y=0.85 $X2=5.925
+ $Y2=1.74
cc_682 N_CON_c_998_n N_S_c_1322_n 0.00863446f $X=6.41 $Y=2.26 $X2=5.925 $Y2=1.74
cc_683 N_CON_c_1006_n N_S_c_1322_n 0.00569656f $X=5.995 $Y=1.37 $X2=5.925
+ $Y2=1.74
cc_684 CON N_S_c_1322_n 7.15106e-19 $X=6.14 $Y=1.37 $X2=5.925 $Y2=1.74
cc_685 N_CON_M1010_g N_S_c_1328_n 9.292e-19 $X=6.535 $Y=3.235 $X2=5.925 $Y2=2.77
cc_686 N_CON_M1023_g N_CO_c_1368_n 0.0434637f $X=6.535 $Y=0.85 $X2=6.75
+ $Y2=0.755
cc_687 N_CON_c_998_n N_CO_c_1368_n 0.0686303f $X=6.41 $Y=2.26 $X2=6.75 $Y2=0.755
cc_688 N_CON_c_1001_n N_CO_c_1368_n 0.0122992f $X=6.41 $Y=1.37 $X2=6.75
+ $Y2=0.755
cc_689 CON N_CO_c_1368_n 0.00209642f $X=6.14 $Y=1.37 $X2=6.75 $Y2=0.755
cc_690 N_CON_M1010_g CO 0.00944261f $X=6.535 $Y=3.235 $X2=6.75 $Y2=2.48
cc_691 N_CON_c_993_n CO 0.00612215f $X=6.41 $Y=2.26 $X2=6.75 $Y2=2.48
cc_692 N_CON_c_998_n CO 0.0017516f $X=6.41 $Y=2.26 $X2=6.75 $Y2=2.48
cc_693 N_CON_c_999_n N_A_27_115#_c_1387_n 0.00774941f $X=1.665 $Y=1.2 $X2=1.035
+ $Y2=1.16
cc_694 N_CON_c_994_n N_A_27_115#_c_1390_n 2.23682e-19 $X=1.55 $Y=0.755 $X2=1.12
+ $Y2=0.755
cc_695 N_CON_M1015_g N_A_526_115#_c_1415_n 0.00145663f $X=3.845 $Y=0.85
+ $X2=3.545 $Y2=1.115
cc_696 N_CON_c_1000_n N_A_526_115#_c_1415_n 0.00251315f $X=3.845 $Y=1.455
+ $X2=3.545 $Y2=1.115
cc_697 N_CON_c_1003_n N_A_526_115#_c_1415_n 0.038473f $X=3.855 $Y=1.37 $X2=3.545
+ $Y2=1.115
cc_698 N_CON_c_1003_n N_A_526_115#_c_1418_n 0.00984552f $X=3.855 $Y=1.37
+ $X2=2.855 $Y2=1.115
cc_699 N_CON_M1015_g N_A_526_115#_c_1419_n 3.73968e-19 $X=3.845 $Y=0.85 $X2=3.63
+ $Y2=0.755
cc_700 N_A_784_115#_c_1181_n A_870_521# 0.00836716f $X=5.33 $Y=2.855 $X2=4.35
+ $Y2=2.605
cc_701 N_A_784_115#_c_1181_n A_952_521# 0.00920662f $X=5.33 $Y=2.855 $X2=4.76
+ $Y2=2.605
cc_702 N_A_784_115#_M1018_g N_S_c_1317_n 0.0186398f $X=5.585 $Y=0.85 $X2=5.8
+ $Y2=0.755
cc_703 N_A_784_115#_M1007_g N_S_c_1323_n 0.00542992f $X=5.585 $Y=3.235 $X2=5.8
+ $Y2=3.295
cc_704 N_A_784_115#_M1018_g N_S_c_1321_n 0.00949101f $X=5.585 $Y=0.85 $X2=5.925
+ $Y2=2.685
cc_705 N_A_784_115#_M1007_g N_S_c_1321_n 0.00506137f $X=5.585 $Y=3.235 $X2=5.925
+ $Y2=2.685
cc_706 N_A_784_115#_c_1161_n N_S_c_1321_n 0.00346737f $X=5.585 $Y=2.275
+ $X2=5.925 $Y2=2.685
cc_707 N_A_784_115#_c_1183_n N_S_c_1321_n 0.0093653f $X=5.415 $Y=2.77 $X2=5.925
+ $Y2=2.685
cc_708 N_A_784_115#_c_1169_n N_S_c_1321_n 0.0246408f $X=5.415 $Y=2.275 $X2=5.925
+ $Y2=2.685
cc_709 N_A_784_115#_M1018_g N_S_c_1322_n 0.00451626f $X=5.585 $Y=0.85 $X2=5.925
+ $Y2=1.74
cc_710 N_A_784_115#_M1007_g N_S_c_1328_n 0.00309508f $X=5.585 $Y=3.235 $X2=5.925
+ $Y2=2.77
cc_711 N_A_784_115#_M1007_g S 0.0115125f $X=5.585 $Y=3.235 $X2=5.8 $Y2=2.855
cc_712 N_A_784_115#_c_1161_n S 0.00106713f $X=5.585 $Y=2.275 $X2=5.8 $Y2=2.855
cc_713 N_A_784_115#_c_1181_n S 0.00567717f $X=5.33 $Y=2.855 $X2=5.8 $Y2=2.855
cc_714 N_A_784_115#_c_1183_n S 7.73713e-19 $X=5.415 $Y=2.77 $X2=5.8 $Y2=2.855
cc_715 N_A_784_115#_c_1169_n S 0.00443271f $X=5.415 $Y=2.275 $X2=5.8 $Y2=2.855
cc_716 N_A_784_115#_c_1165_n N_A_526_115#_c_1415_n 0.00394379f $X=4.31 $Y=1.71
+ $X2=3.545 $Y2=1.115
cc_717 N_A_784_115#_c_1166_n N_A_526_115#_c_1419_n 2.24479e-19 $X=4.06 $Y=0.74
+ $X2=3.63 $Y2=0.755
cc_718 N_S_c_1321_n N_CO_c_1368_n 0.00396474f $X=5.925 $Y=2.685 $X2=6.75
+ $Y2=0.755
cc_719 N_S_c_1321_n CO 0.00370359f $X=5.925 $Y=2.685 $X2=6.75 $Y2=2.48
