* File: sky130_osu_sc_12T_ls__buf_4.pex.spice
* Created: Fri Nov 12 15:35:14 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__BUF_4%GND 1 2 3 31 35 39 41 42 49 63 65
r61 63 65 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r62 47 49 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.755
r63 41 47 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.325 $Y=0.152
+ $X2=2.41 $Y2=0.305
r64 37 42 3.38889 $w=3.06e-07 $l=8.6487e-08 $layer=LI1_cond $X=1.55 $Y=0.155
+ $X2=1.635 $Y2=0.152
r65 37 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.755
r66 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r67 31 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r68 31 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r69 31 37 21.1307 $w=3.06e-07 $l=5.3e-07 $layer=LI1_cond $X=1.02 $Y=0.155
+ $X2=1.55 $Y2=0.155
r70 31 33 13.1569 $w=3.06e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=0.155
+ $X2=0.69 $Y2=0.155
r71 31 33 13.9542 $w=3.06e-07 $l=3.5e-07 $layer=LI1_cond $X=0.34 $Y=0.155
+ $X2=0.69 $Y2=0.155
r72 31 41 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r73 31 42 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r74 3 49 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.27 $Y=0.575
+ $X2=2.41 $Y2=0.755
r75 2 39 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41 $Y=0.575
+ $X2=1.55 $Y2=0.755
r76 1 35 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__BUF_4%VDD 1 2 3 25 27 34 36 42 46 53 60 64
r44 60 64 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.7 $Y2=4.287
r45 53 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=2.955
+ $X2=2.41 $Y2=3.635
r46 51 56 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.41 $Y=4.135 $X2=2.41
+ $Y2=3.635
r47 49 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=4.25 $X2=1.7
+ $Y2=4.25
r48 47 58 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=4.287
+ $X2=1.55 $Y2=4.287
r49 47 49 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=4.287
+ $X2=1.7 $Y2=4.287
r50 46 51 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.325 $Y=4.287
+ $X2=2.41 $Y2=4.135
r51 46 49 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=4.287
+ $X2=1.7 $Y2=4.287
r52 42 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r53 40 58 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=4.287
r54 40 45 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.55 $Y=4.135 $X2=1.55
+ $Y2=3.635
r55 37 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r56 37 39 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r57 36 58 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=4.287
+ $X2=1.55 $Y2=4.287
r58 36 39 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=4.287
+ $X2=1.02 $Y2=4.287
r59 32 57 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r60 32 34 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135 $X2=0.69
+ $Y2=3.635
r61 29 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r62 27 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r63 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r64 25 49 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r65 25 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r66 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r67 3 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=3.635
r68 3 53 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=2.955
r69 2 45 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r70 2 42 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r71 1 34 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__BUF_4%A 3 7 10 14 20
r39 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=2.85
+ $X2=0.635 $Y2=2.85
r40 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2 $X2=0.635
+ $Y2=2.85
r41 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635 $Y=2
+ $X2=0.635 $Y2=2
r42 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=2.165
r43 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2
+ $X2=0.585 $Y2=1.835
r44 7 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.475 $Y=3.235
+ $X2=0.475 $Y2=2.165
r45 3 11 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=0.475 $Y=0.835
+ $X2=0.475 $Y2=1.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__BUF_4%A_27_115# 1 3 11 13 15 17 20 22 24 25 26
+ 27 28 31 33 35 36 38 42 44 46 56 57 60 64 68 70 73
c118 33 0 1.33323e-19 $X=1.765 $Y=2.53
c119 31 0 1.33323e-19 $X=1.765 $Y=0.835
c120 22 0 1.33323e-19 $X=1.335 $Y=2.53
c121 20 0 1.33323e-19 $X=1.335 $Y=0.835
r122 69 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.455
+ $X2=0.26 $Y2=1.455
r123 68 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.965 $Y2=1.455
r124 68 69 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.455
+ $X2=0.345 $Y2=1.455
r125 64 66 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r126 62 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.54
+ $X2=0.26 $Y2=1.455
r127 62 64 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=0.26 $Y=1.54
+ $X2=0.26 $Y2=2.955
r128 58 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=1.455
r129 58 60 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.26 $Y=1.37
+ $X2=0.26 $Y2=0.755
r130 53 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.455 $X2=0.965 $Y2=1.455
r131 53 54 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.455
+ $X2=1.18 $Y2=1.455
r132 51 53 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.455
+ $X2=0.965 $Y2=1.455
r133 49 50 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.455
+ $X2=1.335 $Y2=2.455
r134 47 49 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.455
+ $X2=1.18 $Y2=2.455
r135 44 46 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.195 $Y=2.53
+ $X2=2.195 $Y2=3.235
r136 40 42 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.195 $Y=1.29
+ $X2=2.195 $Y2=0.835
r137 39 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.455
+ $X2=1.765 $Y2=2.455
r138 38 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=2.455
+ $X2=2.195 $Y2=2.53
r139 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.455
+ $X2=1.84 $Y2=2.455
r140 37 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.365
+ $X2=1.765 $Y2=1.365
r141 36 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=2.195 $Y2=1.29
r142 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.365
+ $X2=1.84 $Y2=1.365
r143 33 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.53
+ $X2=1.765 $Y2=2.455
r144 33 35 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.765 $Y=2.53
+ $X2=1.765 $Y2=3.235
r145 29 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=1.365
r146 29 31 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.765 $Y=1.29
+ $X2=1.765 $Y2=0.835
r147 28 50 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.455
+ $X2=1.335 $Y2=2.455
r148 27 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.455
+ $X2=1.765 $Y2=2.455
r149 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.455
+ $X2=1.41 $Y2=2.455
r150 25 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.365
+ $X2=1.765 $Y2=1.365
r151 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.365
+ $X2=1.41 $Y2=1.365
r152 22 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.53
+ $X2=1.335 $Y2=2.455
r153 22 24 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.335 $Y=2.53
+ $X2=1.335 $Y2=3.235
r154 18 26 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.41 $Y2=1.365
r155 18 54 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.18 $Y2=1.455
r156 18 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=1.29
+ $X2=1.335 $Y2=0.835
r157 17 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.38
+ $X2=1.18 $Y2=2.455
r158 16 54 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=1.455
r159 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=2.38
r160 13 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=2.455
r161 13 15 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=2.53
+ $X2=0.905 $Y2=3.235
r162 9 51 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=1.455
r163 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=1.29
+ $X2=0.905 $Y2=0.835
r164 3 66 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r165 3 64 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r166 1 60 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__BUF_4%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c84 55 0 1.33323e-19 $X=1.98 $Y=2.365
c85 54 0 1.33323e-19 $X=1.98 $Y=1.115
c86 46 0 1.33323e-19 $X=1.12 $Y=2.365
c87 45 0 1.33323e-19 $X=1.12 $Y=1.115
r88 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.365
+ $X2=1.98 $Y2=2.48
r89 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.115
+ $X2=1.98 $Y2=1
r90 54 55 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.115
+ $X2=1.98 $Y2=2.365
r91 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.48
+ $X2=1.12 $Y2=2.48
r92 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.48
+ $X2=1.98 $Y2=2.48
r93 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.48
+ $X2=1.265 $Y2=2.48
r94 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1
+ $X2=1.12 $Y2=1
r95 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1
+ $X2=1.98 $Y2=1
r96 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1
+ $X2=1.265 $Y2=1
r97 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=2.48
r98 46 48 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.365
+ $X2=1.12 $Y2=1.79
r99 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1
r100 45 48 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.115
+ $X2=1.12 $Y2=1.79
r101 41 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r102 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.48
+ $X2=1.98 $Y2=2.48
r103 38 41 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.98 $Y=2.48
+ $X2=1.98 $Y2=2.955
r104 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1 $X2=1.98
+ $Y2=1
r105 32 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.98 $Y=0.755
+ $X2=1.98 $Y2=1
r106 27 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r107 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.48
r108 24 27 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.12 $Y=2.48
+ $X2=1.12 $Y2=2.955
r109 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1 $X2=1.12
+ $Y2=1
r110 18 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.12 $Y=0.755
+ $X2=1.12 $Y2=1
r111 6 43 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r112 6 41 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r113 5 29 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r114 5 27 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r115 2 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.755
r116 1 18 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.755
.ends

