* File: sky130_osu_sc_18T_hs__dff_1.pex.spice
* Created: Fri Nov 12 13:48:41 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%GND 1 2 3 4 5 81 83 91 93 103 105 115 117
+ 124 126 133 152 154
c171 81 0 1.27355e-19 $X=-0.045 $Y=0
r172 152 154 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r173 131 133 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.545 $Y=0.305
+ $X2=6.545 $Y2=0.825
r174 122 124 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.165 $Y=0.305
+ $X2=5.165 $Y2=0.825
r175 118 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.152
+ $X2=4.215 $Y2=0.152
r176 113 141 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.152
r177 113 115 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.825
r178 105 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.152
+ $X2=4.215 $Y2=0.152
r179 101 103 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.465 $Y=0.305
+ $X2=2.465 $Y2=0.825
r180 94 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.152
+ $X2=0.715 $Y2=0.152
r181 89 137 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.152
r182 89 91 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.825
r183 83 137 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.152
+ $X2=0.715 $Y2=0.152
r184 81 154 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r185 81 152 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r186 81 131 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.545 $Y2=0.305
r187 81 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.46 $Y2=0.152
r188 81 122 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.165 $Y2=0.305
r189 81 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.08 $Y2=0.152
r190 81 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.25 $Y2=0.152
r191 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.465 $Y2=0.305
r192 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.38 $Y2=0.152
r193 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.55 $Y2=0.152
r194 81 126 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.46 $Y2=0.152
r195 81 127 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.25 $Y2=0.152
r196 81 117 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=5.08 $Y2=0.152
r197 81 118 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.3 $Y2=0.152
r198 81 105 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.13 $Y2=0.152
r199 81 106 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.55 $Y2=0.152
r200 81 93 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.38 $Y2=0.152
r201 81 94 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.8 $Y2=0.152
r202 81 83 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.63 $Y2=0.152
r203 5 133 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.405
+ $Y=0.575 $X2=6.545 $Y2=0.825
r204 4 124 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=5.04
+ $Y=0.575 $X2=5.165 $Y2=0.825
r205 3 115 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.075
+ $Y=0.575 $X2=4.215 $Y2=0.825
r206 2 103 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.825
r207 1 91 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.575 $X2=0.715 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%VDD 1 2 3 4 5 61 63 70 74 82 86 94 98 104
+ 108 114 127 130 134
c99 114 0 1.98165e-19 $X=6.545 $Y=3.455
c100 70 0 5.41559e-20 $X=0.715 $Y=3.795
c101 1 0 1.59851e-19 $X=0.575 $Y=3.085
r102 130 134 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=6.46 $Y2=6.507
r103 127 134 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=6.47
+ $X2=6.46 $Y2=6.47
r104 114 117 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.545 $Y=3.455
+ $X2=6.545 $Y2=5.835
r105 112 127 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=6.355
+ $X2=6.545 $Y2=6.507
r106 112 117 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.545 $Y=6.355
+ $X2=6.545 $Y2=5.835
r107 109 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.25 $Y=6.507
+ $X2=5.165 $Y2=6.507
r108 109 111 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.25 $Y=6.507
+ $X2=5.78 $Y2=6.507
r109 108 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=6.507
+ $X2=6.545 $Y2=6.507
r110 108 111 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.46 $Y=6.507
+ $X2=5.78 $Y2=6.507
r111 104 107 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=5.165 $Y=3.795
+ $X2=5.165 $Y2=5.835
r112 102 125 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.165 $Y=6.355
+ $X2=5.165 $Y2=6.507
r113 102 107 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.165 $Y=6.355
+ $X2=5.165 $Y2=5.835
r114 99 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=6.507
+ $X2=4.215 $Y2=6.507
r115 99 101 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.3 $Y=6.507
+ $X2=4.42 $Y2=6.507
r116 98 125 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=6.507
+ $X2=5.165 $Y2=6.507
r117 98 101 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.08 $Y=6.507
+ $X2=4.42 $Y2=6.507
r118 94 97 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.215 $Y=3.455
+ $X2=4.215 $Y2=5.835
r119 92 123 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.215 $Y=6.355
+ $X2=4.215 $Y2=6.507
r120 92 97 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.215 $Y=6.355
+ $X2=4.215 $Y2=5.835
r121 89 91 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=6.507
+ $X2=3.74 $Y2=6.507
r122 87 122 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=6.507
+ $X2=2.465 $Y2=6.507
r123 87 89 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=2.55 $Y=6.507
+ $X2=3.06 $Y2=6.507
r124 86 123 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=6.507
+ $X2=4.215 $Y2=6.507
r125 86 91 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=4.13 $Y=6.507
+ $X2=3.74 $Y2=6.507
r126 82 85 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.465 $Y=3.795
+ $X2=2.465 $Y2=5.835
r127 80 122 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.465 $Y=6.355
+ $X2=2.465 $Y2=6.507
r128 80 85 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.465 $Y=6.355
+ $X2=2.465 $Y2=5.835
r129 77 79 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r130 75 120 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=6.507
+ $X2=0.715 $Y2=6.507
r131 75 77 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=0.8 $Y=6.507
+ $X2=1.02 $Y2=6.507
r132 74 122 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=6.507
+ $X2=2.465 $Y2=6.507
r133 74 79 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=6.507
+ $X2=1.7 $Y2=6.507
r134 70 73 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.715 $Y=3.795
+ $X2=0.715 $Y2=5.835
r135 68 120 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.715 $Y=6.355
+ $X2=0.715 $Y2=6.507
r136 68 73 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.715 $Y=6.355
+ $X2=0.715 $Y2=5.835
r137 65 130 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r138 63 120 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=6.507
+ $X2=0.715 $Y2=6.507
r139 63 65 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.63 $Y=6.507
+ $X2=0.34 $Y2=6.507
r140 61 127 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=6.355 $X2=6.46 $Y2=6.44
r141 61 111 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=6.355 $X2=5.78 $Y2=6.44
r142 61 125 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=6.355 $X2=5.1 $Y2=6.44
r143 61 101 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r144 61 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r145 61 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r146 61 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r147 61 79 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r148 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r149 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r150 5 117 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.405
+ $Y=3.085 $X2=6.545 $Y2=5.835
r151 5 114 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.405
+ $Y=3.085 $X2=6.545 $Y2=3.455
r152 4 107 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=5.04 $Y=3.085 $X2=5.165 $Y2=5.835
r153 4 104 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=5.04 $Y=3.085 $X2=5.165 $Y2=3.795
r154 3 97 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.075
+ $Y=3.085 $X2=4.215 $Y2=5.835
r155 3 94 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.075
+ $Y=3.085 $X2=4.215 $Y2=3.455
r156 2 85 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=2.325 $Y=3.085 $X2=2.465 $Y2=5.835
r157 2 82 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=2.325 $Y=3.085 $X2=2.465 $Y2=3.795
r158 1 73 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=0.575 $Y=3.085 $X2=0.715 $Y2=5.835
r159 1 70 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=0.575 $Y=3.085 $X2=0.715 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%A_75_344# 1 3 13 17 20 22 23 28 29 30 31
+ 32 34 37 41 46 47 50
c86 29 0 1.29912e-19 $X=1.405 $Y=1.765
c87 28 0 1.59851e-19 $X=0.625 $Y=3.1
c88 22 0 5.41559e-20 $X=0.51 $Y=2.765
r89 49 50 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.582 $Y=1.245
+ $X2=1.582 $Y2=1.415
r90 46 48 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.765
+ $X2=0.567 $Y2=2.93
r91 46 47 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.765
+ $X2=0.567 $Y2=2.6
r92 41 43 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.59 $Y=3.455
+ $X2=1.59 $Y2=5.835
r93 39 41 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=1.59 $Y=3.375 $X2=1.59
+ $Y2=3.455
r94 37 49 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.59 $Y=0.825
+ $X2=1.59 $Y2=1.245
r95 34 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.49 $Y=1.68
+ $X2=1.49 $Y2=1.415
r96 31 39 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=1.42 $Y=3.185
+ $X2=1.59 $Y2=3.375
r97 31 32 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.42 $Y=3.185
+ $X2=0.71 $Y2=3.185
r98 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.765
+ $X2=1.49 $Y2=1.68
r99 29 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.405 $Y=1.765
+ $X2=0.71 $Y2=1.765
r100 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=3.1
+ $X2=0.71 $Y2=3.185
r101 28 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.625 $Y=3.1
+ $X2=0.625 $Y2=2.93
r102 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.85
+ $X2=0.71 $Y2=1.765
r103 25 47 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.625 $Y=1.85
+ $X2=0.625 $Y2=2.6
r104 22 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=2.765 $X2=0.51 $Y2=2.765
r105 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.765
+ $X2=0.51 $Y2=2.93
r106 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.765
+ $X2=0.51 $Y2=2.6
r107 20 23 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.45 $Y=1.87
+ $X2=0.45 $Y2=2.6
r108 19 20 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.475 $Y=1.72
+ $X2=0.475 $Y2=1.87
r109 17 24 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.5 $Y=4.585
+ $X2=0.5 $Y2=2.93
r110 13 19 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.5 $Y=1.075
+ $X2=0.5 $Y2=1.72
r111 3 43 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.365
+ $Y=3.085 $X2=1.59 $Y2=5.835
r112 3 41 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.365
+ $Y=3.085 $X2=1.59 $Y2=3.455
r113 1 37 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.365
+ $Y=0.575 $X2=1.59 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%D 3 7 10 14 19
c43 19 0 1.41836e-19 $X=0.99 $Y=2.22
c44 10 0 1.12321e-19 $X=0.99 $Y=2.22
r45 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=2.22
+ $X2=0.99 $Y2=2.22
r46 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.22 $X2=0.99 $Y2=2.22
r47 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=2.22
+ $X2=0.99 $Y2=2.385
r48 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=2.22
+ $X2=0.99 $Y2=2.055
r49 7 12 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.93 $Y=4.585
+ $X2=0.93 $Y2=2.385
r50 3 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.93 $Y=1.075
+ $X2=0.93 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c213 55 0 6.79641e-20 $X=3.185 $Y=2.59
c214 48 0 1.98654e-19 $X=1.83 $Y=1.85
c215 44 0 1.86602e-19 $X=1.745 $Y=2.59
c216 30 0 1.29912e-19 $X=1.83 $Y=1.685
c217 25 0 1.41836e-19 $X=1.35 $Y=2.765
r218 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.725 $Y=2.59
+ $X2=3.58 $Y2=2.59
r219 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.43 $Y=2.59
+ $X2=4.575 $Y2=2.59
r220 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=4.43 $Y=2.59
+ $X2=3.725 $Y2=2.59
r221 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.495 $Y=2.59
+ $X2=1.35 $Y2=2.59
r222 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.435 $Y=2.59
+ $X2=3.58 $Y2=2.59
r223 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=3.435 $Y=2.59
+ $X2=1.495 $Y2=2.59
r224 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.59
+ $X2=3.58 $Y2=2.59
r225 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.58 $Y=2.59
+ $X2=3.58 $Y2=2.765
r226 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.35 $Y=2.59
+ $X2=1.35 $Y2=2.59
r227 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.35 $Y=2.59
+ $X2=1.35 $Y2=2.765
r228 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.575 $Y=2.59
+ $X2=4.575 $Y2=2.59
r229 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.59
+ $X2=4.575 $Y2=2.765
r230 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.59
+ $X2=3.58 $Y2=2.59
r231 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.495 $Y=2.59
+ $X2=3.185 $Y2=2.59
r232 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.505
+ $X2=3.185 $Y2=2.59
r233 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.1 $Y=2.505
+ $X2=3.1 $Y2=1.85
r234 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.83 $Y=2.505
+ $X2=1.83 $Y2=1.85
r235 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.59
+ $X2=1.35 $Y2=2.59
r236 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=2.59
+ $X2=1.83 $Y2=2.505
r237 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.745 $Y=2.59
+ $X2=1.435 $Y2=2.59
r238 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=2.765 $X2=4.575 $Y2=2.765
r239 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=4.457 $Y=1.685
+ $X2=4.457 $Y2=1.835
r240 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=2.765 $X2=3.58 $Y2=2.765
r241 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=2.765
+ $X2=3.58 $Y2=2.93
r242 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.85 $X2=3.1 $Y2=1.85
r243 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.85
+ $X2=3.1 $Y2=1.685
r244 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.85 $X2=1.83 $Y2=1.85
r245 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.85
+ $X2=1.83 $Y2=1.685
r246 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=2.765 $X2=1.35 $Y2=2.765
r247 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=2.765
+ $X2=1.35 $Y2=2.93
r248 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=4.485 $Y=2.6
+ $X2=4.532 $Y2=2.765
r249 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.485 $Y=2.6
+ $X2=4.485 $Y2=1.835
r250 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=4.43 $Y=2.93
+ $X2=4.532 $Y2=2.765
r251 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=4.43 $Y=2.93
+ $X2=4.43 $Y2=4.585
r252 17 40 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.43 $Y=1.075
+ $X2=4.43 $Y2=1.685
r253 13 39 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.64 $Y=4.585
+ $X2=3.64 $Y2=2.93
r254 10 34 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.04 $Y=1.075
+ $X2=3.04 $Y2=1.685
r255 7 30 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.89 $Y=1.075
+ $X2=1.89 $Y2=1.685
r256 3 27 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.29 $Y=4.585
+ $X2=1.29 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%A_32_115# 1 3 11 15 17 18 21 22 27 31 34
+ 37 41 47 52 56 61 62 63 68
c115 47 0 1.5821e-19 $X=2.42 $Y=2.765
c116 31 0 6.36774e-20 $X=2.68 $Y=4.585
c117 22 0 1.86602e-19 $X=2.325 $Y=2.765
c118 21 0 6.79641e-20 $X=2.605 $Y=2.765
c119 15 0 6.36774e-20 $X=2.25 $Y=4.585
r120 63 65 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.43 $Y=1.85
+ $X2=0.285 $Y2=1.85
r121 62 68 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.185 $Y=1.85
+ $X2=2.33 $Y2=1.85
r122 62 63 1.68986 $w=1.7e-07 $l=1.755e-06 $layer=MET1_cond $X=2.185 $Y=1.85
+ $X2=0.43 $Y2=1.85
r123 59 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.33 $Y=1.85
+ $X2=2.33 $Y2=1.85
r124 59 61 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=2.33 $Y=1.81 $X2=2.42
+ $Y2=1.81
r125 54 56 6.22173 $w=2.03e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=3.242
+ $X2=0.285 $Y2=3.242
r126 52 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.285 $Y=1.85
+ $X2=0.285 $Y2=1.85
r127 49 52 4.81931 $w=2.73e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=1.797
+ $X2=0.285 $Y2=1.797
r128 45 61 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.42 $Y=1.935
+ $X2=2.42 $Y2=1.81
r129 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.42 $Y=1.935
+ $X2=2.42 $Y2=2.765
r130 41 43 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.285 $Y=3.455
+ $X2=0.285 $Y2=5.835
r131 39 56 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.285 $Y=3.345
+ $X2=0.285 $Y2=3.242
r132 39 41 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.285 $Y=3.345
+ $X2=0.285 $Y2=3.455
r133 35 52 3.55113 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.285 $Y=1.66
+ $X2=0.285 $Y2=1.797
r134 35 37 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.285 $Y=1.66
+ $X2=0.285 $Y2=0.825
r135 34 54 1.83547 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=0.17 $Y=3.14
+ $X2=0.17 $Y2=3.242
r136 33 49 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.17 $Y=1.935
+ $X2=0.17 $Y2=1.797
r137 33 34 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=0.17 $Y=1.935
+ $X2=0.17 $Y2=3.14
r138 29 31 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=2.68 $Y=2.9
+ $X2=2.68 $Y2=4.585
r139 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.68 $Y=1.715
+ $X2=2.68 $Y2=1.075
r140 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=2.765 $X2=2.42 $Y2=2.765
r141 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=2.765
+ $X2=2.42 $Y2=2.765
r142 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=2.765
+ $X2=2.68 $Y2=2.9
r143 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=2.765
+ $X2=2.42 $Y2=2.765
r144 20 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.85 $X2=2.42 $Y2=1.85
r145 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=1.85
+ $X2=2.42 $Y2=1.85
r146 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.605 $Y=1.85
+ $X2=2.68 $Y2=1.715
r147 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=1.85
+ $X2=2.42 $Y2=1.85
r148 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=2.9
+ $X2=2.325 $Y2=2.765
r149 13 15 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=2.25 $Y=2.9
+ $X2=2.25 $Y2=4.585
r150 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=1.715
+ $X2=2.325 $Y2=1.85
r151 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.25 $Y=1.715
+ $X2=2.25 $Y2=1.075
r152 3 43 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.16
+ $Y=3.085 $X2=0.285 $Y2=5.835
r153 3 41 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.16
+ $Y=3.085 $X2=0.285 $Y2=3.455
r154 1 37 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%A_243_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c174 35 0 1.98654e-19 $X=1.41 $Y=1.76
c175 18 0 1.12321e-19 $X=1.89 $Y=4.585
r176 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=3.185
+ $X2=4.915 $Y2=3.185
r177 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=2.19
+ $X2=4.915 $Y2=2.19
r178 60 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=3.1
+ $X2=4.915 $Y2=3.185
r179 59 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.275
+ $X2=4.915 $Y2=2.19
r180 59 60 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.915 $Y=2.275
+ $X2=4.915 $Y2=3.1
r181 55 57 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.645 $Y=3.455
+ $X2=4.645 $Y2=5.835
r182 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=3.27
+ $X2=4.645 $Y2=3.185
r183 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.645 $Y=3.27
+ $X2=4.645 $Y2=3.455
r184 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=2.105
+ $X2=4.645 $Y2=2.19
r185 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.935
+ $X2=4.645 $Y2=1.85
r186 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.645 $Y=1.935
+ $X2=4.645 $Y2=2.105
r187 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=1.85
r188 47 49 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=0.825
r189 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=1.85
+ $X2=4.645 $Y2=1.85
r190 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.56 $Y=1.85
+ $X2=3.58 $Y2=1.85
r191 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.85 $X2=3.58 $Y2=1.85
r192 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.85
+ $X2=3.58 $Y2=2.015
r193 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.85
+ $X2=3.58 $Y2=1.685
r194 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.29 $Y=1.76
+ $X2=1.41 $Y2=1.76
r195 32 41 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.64 $Y=1.075
+ $X2=3.64 $Y2=1.685
r196 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.52 $Y=2.225
+ $X2=3.52 $Y2=2.015
r197 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.115 $Y=2.3
+ $X2=3.04 $Y2=2.3
r198 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.445 $Y=2.3
+ $X2=3.52 $Y2=2.225
r199 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.445 $Y=2.3
+ $X2=3.115 $Y2=2.3
r200 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.04 $Y=2.375
+ $X2=3.04 $Y2=2.3
r201 22 24 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=3.04 $Y=2.375
+ $X2=3.04 $Y2=4.585
r202 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=2.3
+ $X2=1.89 $Y2=2.3
r203 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.965 $Y=2.3
+ $X2=3.04 $Y2=2.3
r204 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.965 $Y=2.3
+ $X2=1.965 $Y2=2.3
r205 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=2.375
+ $X2=1.89 $Y2=2.3
r206 16 18 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=1.89 $Y=2.375
+ $X2=1.89 $Y2=4.585
r207 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=2.3
+ $X2=1.89 $Y2=2.3
r208 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.815 $Y=2.3
+ $X2=1.485 $Y2=2.3
r209 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=2.225
+ $X2=1.485 $Y2=2.3
r210 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.835
+ $X2=1.41 $Y2=1.76
r211 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.41 $Y=1.835
+ $X2=1.41 $Y2=2.225
r212 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.685
+ $X2=1.29 $Y2=1.76
r213 9 11 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.29 $Y=1.685
+ $X2=1.29 $Y2=1.075
r214 3 57 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.505
+ $Y=3.085 $X2=4.645 $Y2=5.835
r215 3 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.505
+ $Y=3.085 $X2=4.645 $Y2=3.455
r216 1 49 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.505
+ $Y=0.575 $X2=4.645 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%A_785_89# 1 3 11 15 23 26 28 32 33 35 36
+ 37 38 40 46 50 56 59 60 61 66
c131 37 0 8.77106e-20 $X=6.305 $Y=2.855
c132 32 0 2.20654e-19 $X=6.215 $Y=2.19
r133 61 63 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.205 $Y=2.19
+ $X2=4.06 $Y2=2.19
r134 60 66 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.07 $Y=2.19
+ $X2=6.215 $Y2=2.19
r135 60 61 1.79578 $w=1.7e-07 $l=1.865e-06 $layer=MET1_cond $X=6.07 $Y=2.19
+ $X2=4.205 $Y2=2.19
r136 56 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=2.19
+ $X2=6.215 $Y2=2.19
r137 54 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=2.19
+ $X2=5.595 $Y2=2.19
r138 54 56 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.68 $Y=2.19
+ $X2=6.215 $Y2=2.19
r139 50 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.595 $Y=3.455
+ $X2=5.595 $Y2=5.835
r140 48 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=2.275
+ $X2=5.595 $Y2=2.19
r141 48 50 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=5.595 $Y=2.275
+ $X2=5.595 $Y2=3.455
r142 44 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=2.105
+ $X2=5.595 $Y2=2.19
r143 44 46 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=5.595 $Y=2.105
+ $X2=5.595 $Y2=0.825
r144 40 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.06 $Y=2.19
+ $X2=4.06 $Y2=2.19
r145 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=2.855
+ $X2=6.305 $Y2=3.005
r146 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=1.65
+ $X2=6.305 $Y2=1.8
r147 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.28 $Y=2.355
+ $X2=6.28 $Y2=2.855
r148 33 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.28 $Y=2.025
+ $X2=6.28 $Y2=1.8
r149 32 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=2.19 $X2=6.215 $Y2=2.19
r150 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.217 $Y=2.19
+ $X2=6.217 $Y2=2.355
r151 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.217 $Y=2.19
+ $X2=6.217 $Y2=2.025
r152 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=2.19 $X2=4.06 $Y2=2.19
r153 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=2.19
+ $X2=4.06 $Y2=2.355
r154 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=2.19
+ $X2=4.06 $Y2=2.025
r155 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=6.33 $Y=4.585
+ $X2=6.33 $Y2=3.005
r156 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.33 $Y=1.075
+ $X2=6.33 $Y2=1.65
r157 15 30 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=4 $Y=4.585 $X2=4
+ $Y2=2.355
r158 11 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4 $Y=1.075 $X2=4
+ $Y2=2.025
r159 3 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5.455
+ $Y=3.085 $X2=5.595 $Y2=5.835
r160 3 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5.455
+ $Y=3.085 $X2=5.595 $Y2=3.455
r161 1 46 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.455
+ $Y=0.575 $X2=5.595 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%A_623_115# 1 3 9 11 14 19 24 25 26 27 28
+ 31 35 40 44 45 50
c115 45 0 1.5821e-19 $X=2.905 $Y=1.85
c116 24 0 1.57671e-19 $X=2.76 $Y=1.85
r117 45 47 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.905 $Y=1.85
+ $X2=2.76 $Y2=1.85
r118 44 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.85
+ $X2=5.175 $Y2=1.85
r119 44 45 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=5.03 $Y=1.85
+ $X2=2.905 $Y2=1.85
r120 40 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.85
+ $X2=5.175 $Y2=1.85
r121 35 37 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=3.34 $Y=3.455
+ $X2=3.34 $Y2=5.835
r122 33 35 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=3.34 $Y=3.27
+ $X2=3.34 $Y2=3.455
r123 29 31 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=3.34 $Y=1.345
+ $X2=3.34 $Y2=0.825
r124 27 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=3.185
+ $X2=3.34 $Y2=3.27
r125 27 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=3.185
+ $X2=2.845 $Y2=3.185
r126 25 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=1.43
+ $X2=3.34 $Y2=1.345
r127 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=1.43
+ $X2=2.845 $Y2=1.43
r128 24 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.76 $Y=1.85
+ $X2=2.76 $Y2=1.85
r129 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=3.1
+ $X2=2.845 $Y2=3.185
r130 22 24 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.76 $Y=3.1
+ $X2=2.76 $Y2=1.85
r131 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.76 $Y=1.515
+ $X2=2.845 $Y2=1.43
r132 21 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.76 $Y=1.515
+ $X2=2.76 $Y2=1.85
r133 17 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.85 $X2=5.175 $Y2=1.85
r134 17 19 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.175 $Y=1.85
+ $X2=5.38 $Y2=1.85
r135 12 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=2.015
+ $X2=5.38 $Y2=1.85
r136 12 14 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=5.38 $Y=2.015
+ $X2=5.38 $Y2=4.585
r137 9 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.685
+ $X2=5.38 $Y2=1.85
r138 9 11 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.38 $Y=1.685
+ $X2=5.38 $Y2=1.075
r139 3 37 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=3.115
+ $Y=3.085 $X2=3.34 $Y2=5.835
r140 3 35 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=3.115
+ $Y=3.085 $X2=3.34 $Y2=3.455
r141 1 31 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=3.115
+ $Y=0.575 $X2=3.34 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c75 44 0 8.77106e-20 $X=6.12 $Y=2.96
c76 35 0 9.99996e-20 $X=6.615 $Y=2.765
c77 33 0 1.20654e-19 $X=6.615 $Y=1.85
c78 18 0 1.98165e-19 $X=6.7 $Y=2.395
r79 42 44 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=6.115 $Y=2.96
+ $X2=6.12 $Y2=2.96
r80 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.7 $Y=2.68 $X2=6.7
+ $Y2=2.395
r81 37 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.7 $Y=1.935 $X2=6.7
+ $Y2=2.395
r82 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=2.765
+ $X2=6.7 $Y2=2.68
r83 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=2.765
+ $X2=6.2 $Y2=2.765
r84 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=1.85
+ $X2=6.7 $Y2=1.935
r85 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=1.85
+ $X2=6.2 $Y2=1.85
r86 29 31 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.115 $Y=3.455
+ $X2=6.115 $Y2=5.835
r87 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.115 $Y=2.96
+ $X2=6.115 $Y2=2.96
r88 27 29 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.115 $Y=2.96
+ $X2=6.115 $Y2=3.455
r89 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=2.85
+ $X2=6.2 $Y2=2.765
r90 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.115 $Y=2.85
+ $X2=6.115 $Y2=2.96
r91 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=1.765
+ $X2=6.2 $Y2=1.85
r92 21 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.115 $Y=1.765
+ $X2=6.115 $Y2=0.825
r93 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=2.395 $X2=6.7 $Y2=2.395
r94 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.395
+ $X2=6.7 $Y2=2.56
r95 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.395
+ $X2=6.7 $Y2=2.23
r96 15 20 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=6.76 $Y=4.585
+ $X2=6.76 $Y2=2.56
r97 11 19 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=6.76 $Y=1.075
+ $X2=6.76 $Y2=2.23
r98 3 31 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=5.99
+ $Y=3.085 $X2=6.115 $Y2=5.835
r99 3 29 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=5.99
+ $Y=3.085 $X2=6.115 $Y2=3.455
r100 1 23 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=5.99
+ $Y=0.575 $X2=6.115 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFF_1%Q 1 3 11 17 22 25 29 32
r20 27 29 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=3.245
+ $X2=7.09 $Y2=3.245
r21 23 25 7.08586 $w=1.78e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=1.52
+ $X2=7.09 $Y2=1.52
r22 22 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=3.16
+ $X2=7.09 $Y2=3.245
r23 21 25 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.09 $Y=1.61 $X2=7.09
+ $Y2=1.52
r24 21 22 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=7.09 $Y=1.61
+ $X2=7.09 $Y2=3.16
r25 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.975 $Y=3.455
+ $X2=6.975 $Y2=5.835
r26 15 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.975 $Y=3.33
+ $X2=6.975 $Y2=3.33
r27 15 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=6.975 $Y2=3.245
r28 15 17 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=6.975 $Y2=3.455
r29 9 23 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.975 $Y=1.43 $X2=6.975
+ $Y2=1.52
r30 9 11 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.975 $Y=1.43
+ $X2=6.975 $Y2=0.825
r31 3 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.835
+ $Y=3.085 $X2=6.975 $Y2=5.835
r32 3 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.835
+ $Y=3.085 $X2=6.975 $Y2=3.455
r33 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.835
+ $Y=0.575 $X2=6.975 $Y2=0.825
.ends

