magic
tech sky130A
magscale 1 2
timestamp 1606864622
<< checkpaint >>
rect -1209 -1243 1753 2575
<< nwell >>
rect -9 581 638 1341
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 238 617 268 1217
rect 358 617 388 1217
rect 430 617 460 1217
rect 516 617 546 1217
<< nmoslvt >>
rect 80 115 110 315
rect 166 115 196 315
rect 238 115 268 315
rect 358 115 388 315
rect 430 115 460 315
rect 516 115 546 315
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 199 166 315
rect 110 131 121 199
rect 155 131 166 199
rect 110 115 166 131
rect 196 115 238 315
rect 268 267 358 315
rect 268 131 279 267
rect 347 131 358 267
rect 268 115 358 131
rect 388 115 430 315
rect 460 199 516 315
rect 460 131 471 199
rect 505 131 516 199
rect 460 115 516 131
rect 546 267 599 315
rect 546 131 557 267
rect 591 131 599 267
rect 546 115 599 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 657 35 1201
rect 69 657 80 1201
rect 27 617 80 657
rect 110 1201 166 1217
rect 110 657 121 1201
rect 155 657 166 1201
rect 110 617 166 657
rect 196 617 238 1217
rect 268 1201 358 1217
rect 268 657 279 1201
rect 347 657 358 1201
rect 268 617 358 657
rect 388 617 430 1217
rect 460 1201 516 1217
rect 460 657 471 1201
rect 505 657 516 1201
rect 460 617 516 657
rect 546 1201 599 1217
rect 546 658 557 1201
rect 591 658 599 1201
rect 546 617 599 658
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 199
rect 279 131 347 267
rect 471 131 505 199
rect 557 131 591 267
<< pdiffc >>
rect 35 657 69 1201
rect 121 657 155 1201
rect 279 657 347 1201
rect 471 657 505 1201
rect 557 658 591 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 238 1217 268 1243
rect 358 1217 388 1243
rect 430 1217 460 1243
rect 516 1217 546 1243
rect 80 602 110 617
rect 70 572 110 602
rect 70 360 100 572
rect 166 511 196 617
rect 142 495 196 511
rect 142 461 152 495
rect 186 461 196 495
rect 142 445 196 461
rect 238 586 268 617
rect 238 570 292 586
rect 238 536 248 570
rect 282 536 292 570
rect 238 520 292 536
rect 142 387 196 403
rect 142 360 152 387
rect 70 353 152 360
rect 186 353 196 387
rect 70 330 196 353
rect 80 315 110 330
rect 166 315 196 330
rect 238 315 268 520
rect 358 511 388 617
rect 430 602 460 617
rect 516 602 546 617
rect 430 572 546 602
rect 358 495 472 511
rect 358 481 428 495
rect 418 461 428 481
rect 462 461 472 495
rect 418 445 472 461
rect 516 403 546 572
rect 326 387 380 403
rect 326 353 336 387
rect 370 360 380 387
rect 479 387 546 403
rect 479 360 489 387
rect 370 353 388 360
rect 326 337 388 353
rect 358 315 388 337
rect 430 353 489 360
rect 523 353 546 387
rect 430 330 546 353
rect 430 315 460 330
rect 516 315 546 330
rect 80 89 110 115
rect 166 89 196 115
rect 238 89 268 115
rect 358 89 388 115
rect 430 89 460 115
rect 516 89 546 115
<< polycont >>
rect 152 461 186 495
rect 248 536 282 570
rect 152 353 186 387
rect 428 461 462 495
rect 336 353 370 387
rect 489 353 523 387
<< locali >>
rect 0 1311 638 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 638 1311
rect 35 1201 69 1217
rect 35 495 69 657
rect 121 1201 155 1271
rect 279 1201 347 1217
rect 121 641 155 657
rect 268 683 279 689
rect 302 649 347 657
rect 279 641 347 649
rect 471 1201 505 1271
rect 471 641 505 657
rect 557 1201 591 1217
rect 557 570 591 658
rect 232 536 248 570
rect 282 536 591 570
rect 35 461 152 495
rect 186 461 370 495
rect 35 267 69 461
rect 152 387 186 403
rect 336 387 370 461
rect 152 313 186 353
rect 268 283 302 353
rect 336 337 370 353
rect 412 461 428 495
rect 462 461 478 495
rect 412 313 446 461
rect 489 387 523 403
rect 489 337 523 353
rect 268 267 347 283
rect 268 249 279 267
rect 35 115 69 131
rect 121 199 155 215
rect 121 61 155 131
rect 557 267 591 536
rect 279 115 347 131
rect 471 199 505 215
rect 471 61 505 131
rect 557 115 591 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 638 61
rect 0 0 638 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 268 657 279 683
rect 279 657 302 683
rect 268 649 302 657
rect 152 279 186 313
rect 268 353 302 387
rect 489 353 523 387
rect 412 279 446 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1311 638 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 638 1311
rect 0 1271 638 1277
rect 256 683 314 689
rect 256 649 268 683
rect 302 649 314 683
rect 256 643 314 649
rect 268 393 302 643
rect 256 387 314 393
rect 477 387 535 393
rect 256 353 268 387
rect 302 353 314 387
rect 455 353 489 387
rect 523 353 535 387
rect 256 347 314 353
rect 477 347 535 353
rect 140 313 198 319
rect 400 313 458 319
rect 140 279 152 313
rect 186 279 412 313
rect 446 279 458 313
rect 140 273 198 279
rect 400 273 458 279
rect 0 55 638 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 638 55
rect 0 0 638 21
<< labels >>
rlabel metal1 170 296 170 296 1 A
port 1 n
rlabel metal1 506 370 506 370 1 B
port 2 n
rlabel metal1 284 427 284 427 1 Y
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
