magic
tech sky130A
magscale 1 2
timestamp 1606864590
<< checkpaint >>
rect -1209 -1243 1753 2575
<< nwell >>
rect -9 581 638 1341
<< nmos >>
rect 80 115 110 315
rect 152 115 182 315
rect 252 115 282 315
rect 338 115 368 315
rect 424 115 454 315
rect 510 115 540 315
<< pmoshvt >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
rect 338 617 368 1217
rect 424 617 454 1217
rect 510 617 540 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 115 152 315
rect 182 267 252 315
rect 182 131 193 267
rect 227 131 252 267
rect 182 115 252 131
rect 282 267 338 315
rect 282 131 293 267
rect 327 131 338 267
rect 282 115 338 131
rect 368 267 424 315
rect 368 131 379 267
rect 413 131 424 267
rect 368 115 424 131
rect 454 267 510 315
rect 454 131 465 267
rect 499 131 510 267
rect 454 115 510 131
rect 540 267 593 315
rect 540 131 551 267
rect 585 131 593 267
rect 540 115 593 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 166 1217
rect 110 725 121 1201
rect 155 725 166 1201
rect 110 617 166 725
rect 196 1201 252 1217
rect 196 725 207 1201
rect 241 725 252 1201
rect 196 617 252 725
rect 282 1201 338 1217
rect 282 657 293 1201
rect 327 657 338 1201
rect 282 617 338 657
rect 368 1201 424 1217
rect 368 657 379 1201
rect 413 657 424 1201
rect 368 617 424 657
rect 454 1201 510 1217
rect 454 657 465 1201
rect 499 657 510 1201
rect 454 617 510 657
rect 540 1201 593 1217
rect 540 657 551 1201
rect 585 657 593 1201
rect 540 617 593 657
<< ndiffc >>
rect 35 131 69 267
rect 193 131 227 267
rect 293 131 327 267
rect 379 131 413 267
rect 465 131 499 267
rect 551 131 585 267
<< pdiffc >>
rect 35 793 69 1201
rect 121 725 155 1201
rect 207 725 241 1201
rect 293 657 327 1201
rect 379 657 413 1201
rect 465 657 499 1201
rect 551 657 585 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 338 1217 368 1244
rect 424 1217 454 1243
rect 510 1217 540 1243
rect 80 586 110 617
rect 27 570 110 586
rect 27 536 37 570
rect 71 536 110 570
rect 27 520 110 536
rect 80 315 110 520
rect 166 518 196 617
rect 252 592 282 617
rect 338 592 368 617
rect 424 592 454 617
rect 510 592 540 617
rect 252 562 540 592
rect 152 502 217 518
rect 152 468 173 502
rect 207 468 217 502
rect 152 452 217 468
rect 152 315 182 452
rect 259 420 289 562
rect 259 404 313 420
rect 259 384 269 404
rect 252 370 269 384
rect 303 384 313 404
rect 303 370 540 384
rect 252 354 540 370
rect 252 315 282 354
rect 338 315 368 354
rect 424 315 454 354
rect 510 315 540 354
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
rect 338 89 368 115
rect 424 89 454 115
rect 510 89 540 115
<< polycont >>
rect 37 536 71 570
rect 173 468 207 502
rect 269 370 303 404
<< locali >>
rect 0 1311 638 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 638 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 105 725 121 743
rect 105 709 155 725
rect 207 1201 241 1271
rect 207 709 241 725
rect 293 1201 327 1217
rect 37 570 71 649
rect 37 520 71 536
rect 105 404 139 709
rect 173 502 207 575
rect 293 535 327 657
rect 379 1201 413 1271
rect 379 641 413 657
rect 465 1201 499 1217
rect 465 535 499 657
rect 551 1201 585 1271
rect 551 641 585 657
rect 173 452 207 468
rect 35 370 269 404
rect 303 370 319 404
rect 35 267 69 370
rect 35 115 69 131
rect 193 267 227 283
rect 193 61 227 131
rect 293 267 327 279
rect 293 115 327 131
rect 379 267 413 283
rect 379 61 413 131
rect 465 267 499 279
rect 465 115 499 131
rect 551 267 585 283
rect 551 61 585 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 638 61
rect 0 0 638 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 37 649 71 683
rect 173 575 207 609
rect 293 501 327 535
rect 465 501 499 535
rect 293 279 327 313
rect 465 279 499 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1311 638 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 638 1311
rect 0 1271 638 1277
rect 25 683 83 689
rect 25 649 37 683
rect 71 649 105 683
rect 25 643 83 649
rect 161 609 219 615
rect 140 575 173 609
rect 207 575 219 609
rect 161 569 219 575
rect 281 535 339 541
rect 453 535 511 541
rect 281 501 293 535
rect 327 501 465 535
rect 499 501 511 535
rect 281 495 339 501
rect 453 495 511 501
rect 293 319 327 495
rect 465 319 499 495
rect 281 313 339 319
rect 453 313 511 319
rect 281 279 293 313
rect 327 279 465 313
rect 499 279 511 313
rect 281 273 339 279
rect 453 273 511 279
rect 0 55 638 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 638 55
rect 0 0 638 21
<< labels >>
rlabel metal1 311 444 311 444 1 Y
port 1 n
rlabel metal1 55 666 55 666 1 A
port 2 n
rlabel metal1 191 592 191 592 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
