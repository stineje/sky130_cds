* File: sky130_osu_sc_12T_ls__ant.pxi.spice
* Created: Fri Nov 12 15:34:32 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__ANT%GND N_GND_M1001_b N_GND_c_2_p N_GND_c_7_p GND
+ PM_SKY130_OSU_SC_12T_LS__ANT%GND
x_PM_SKY130_OSU_SC_12T_LS__ANT%VDD N_VDD_M1000_d N_VDD_M1000_b N_VDD_c_18_p
+ N_VDD_c_19_p VDD PM_SKY130_OSU_SC_12T_LS__ANT%VDD
x_PM_SKY130_OSU_SC_12T_LS__ANT%A N_A_M1001_s N_A_M1000_s N_A_M1001_g N_A_M1000_g
+ N_A_c_27_n N_A_c_28_n N_A_c_31_n N_A_c_32_n N_A_c_33_n N_A_c_34_n N_A_c_37_n
+ N_A_c_38_n A PM_SKY130_OSU_SC_12T_LS__ANT%A
cc_1 N_GND_M1001_b N_A_M1001_g 0.0789999f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1001_g 0.00607478f $X=0.34 $Y=0.19 $X2=0.475 $Y2=0.835
cc_3 N_GND_M1001_b N_A_M1000_g 0.0125577f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_4 N_GND_M1001_b N_A_c_27_n 0.0562319f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.11
cc_5 N_GND_M1001_b N_A_c_28_n 0.0162383f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.755
cc_6 N_GND_c_2_p N_A_c_28_n 0.00739457f $X=0.34 $Y=0.19 $X2=0.26 $Y2=0.755
cc_7 N_GND_c_7_p N_A_c_28_n 0.00138205f $X=0.34 $Y=0.19 $X2=0.26 $Y2=0.755
cc_8 N_GND_M1001_b N_A_c_31_n 0.0149833f $X=-0.045 $Y=0 $X2=0.26 $Y2=2.025
cc_9 N_GND_M1001_b N_A_c_32_n 0.00651531f $X=-0.045 $Y=0 $X2=0.26 $Y2=2.955
cc_10 N_GND_M1001_b N_A_c_33_n 0.0199494f $X=-0.045 $Y=0 $X2=0.605 $Y2=1.52
cc_11 N_GND_M1001_b N_A_c_34_n 0.0162383f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.755
cc_12 N_GND_c_2_p N_A_c_34_n 0.00761023f $X=0.34 $Y=0.19 $X2=0.69 $Y2=0.755
cc_13 N_GND_c_7_p N_A_c_34_n 0.00138205f $X=0.34 $Y=0.19 $X2=0.69 $Y2=0.755
cc_14 N_GND_M1001_b N_A_c_37_n 0.0076399f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.11
cc_15 N_GND_M1001_b N_A_c_38_n 0.00710193f $X=-0.045 $Y=0 $X2=0.26 $Y2=1.52
cc_16 N_GND_M1001_b A 0.00241298f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.11
cc_17 N_VDD_M1000_b N_A_M1000_g 0.0299903f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_18 N_VDD_c_18_p N_A_M1000_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=3.235
cc_19 N_VDD_c_19_p N_A_M1000_g 0.00636672f $X=0.69 $Y=2.955 $X2=0.475 $Y2=3.235
cc_20 VDD N_A_M1000_g 0.00468827f $X=0.34 $Y=4.2 $X2=0.475 $Y2=3.235
cc_21 N_VDD_M1000_b N_A_c_32_n 0.0103018f $X=-0.045 $Y=2.425 $X2=0.26 $Y2=2.955
cc_22 N_VDD_c_18_p N_A_c_32_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26 $Y2=2.955
cc_23 VDD N_A_c_32_n 0.00476261f $X=0.34 $Y=4.2 $X2=0.26 $Y2=2.955
