* File: sky130_osu_sc_18T_hs__inv_6.pex.spice
* Created: Thu Oct 29 17:08:37 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__INV_6%GND 1 2 3 4 29 33 35 42 44 51 55 60 65 67
r82 65 67 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r83 58 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r84 53 60 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.755 $Y2=0.152
r85 53 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.825
r86 49 59 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r87 49 51 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r88 45 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r89 44 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r90 40 57 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r91 40 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r92 35 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r93 31 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r94 29 31 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r95 29 36 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r96 29 60 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r97 29 58 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r98 29 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.17
+ $X2=2.38 $Y2=0.17
r99 29 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r100 29 44 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r101 29 45 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r102 29 35 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r103 29 36 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r104 4 55 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r105 3 51 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r106 2 42 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r107 1 33 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__INV_6%VDD 1 2 3 4 25 29 33 39 43 49 55 62 64 69
r58 69 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=6.49
+ $X2=2.38 $Y2=6.49
r59 64 69 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=2.38 $Y2=6.507
r60 64 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r61 62 73 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=6.507
+ $X2=2.38 $Y2=6.507
r62 60 73 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=2.38 $Y2=6.507
r63 60 61 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=6.507
+ $X2=1.98 $Y2=6.507
r64 55 58 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r65 53 62 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.755 $Y2=6.507
r66 53 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.84 $Y=6.355
+ $X2=2.84 $Y2=5.835
r67 49 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r68 47 61 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=6.507
r69 47 52 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r70 44 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r71 44 46 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r72 43 61 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.98 $Y2=6.507
r73 43 46 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r74 39 42 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r75 37 59 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r76 37 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r77 34 67 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r78 34 36 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r79 33 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r80 33 36 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r81 29 32 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r82 27 67 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r83 27 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r84 25 67 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r85 25 73 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r86 25 46 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r87 25 36 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r88 4 58 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r89 4 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r90 3 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r91 3 49 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r92 2 42 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r93 2 39 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r94 1 32 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r95 1 29 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__INV_6%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 45 47 49 50 52 53 55 57 59 60 62 63 64 65 66
+ 67 68 69 70 71 72 73 75 76 80 83 85
c179 50 0 1.33323e-19 $X=2.195 $Y=2.96
c180 45 0 1.33323e-19 $X=2.195 $Y=1.7
c181 38 0 1.33323e-19 $X=1.765 $Y=2.96
c182 35 0 1.33323e-19 $X=1.765 $Y=1.7
c183 28 0 1.33323e-19 $X=1.335 $Y=2.96
c184 25 0 1.33323e-19 $X=1.335 $Y=1.7
c185 18 0 1.33323e-19 $X=0.905 $Y=2.96
c186 15 0 1.33323e-19 $X=0.905 $Y=1.7
r187 80 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r188 78 83 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.39
+ $X2=0.32 $Y2=3.33
r189 76 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.47
r190 76 85 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.14
r191 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.305 $X2=0.535 $Y2=2.305
r192 73 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.405 $Y=2.305
+ $X2=0.32 $Y2=2.39
r193 73 75 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.305
+ $X2=0.535 $Y2=2.305
r194 60 62 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.625 $Y=2.96
+ $X2=2.625 $Y2=4.585
r195 57 59 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.625 $Y=1.7
+ $X2=2.625 $Y2=1.075
r196 56 72 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.885
+ $X2=2.195 $Y2=2.885
r197 55 60 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.625 $Y2=2.96
r198 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.885
+ $X2=2.27 $Y2=2.885
r199 54 71 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.775
+ $X2=2.195 $Y2=1.775
r200 53 57 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=1.775
+ $X2=2.625 $Y2=1.7
r201 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.775
+ $X2=2.27 $Y2=1.775
r202 50 72 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=2.885
r203 50 52 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.195 $Y=2.96
+ $X2=2.195 $Y2=4.585
r204 49 72 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.81
+ $X2=2.195 $Y2=2.885
r205 48 71 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.85
+ $X2=2.195 $Y2=1.775
r206 48 49 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.85
+ $X2=2.195 $Y2=2.81
r207 45 71 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.7 $X2=2.195
+ $Y2=1.775
r208 45 47 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.195 $Y=1.7
+ $X2=2.195 $Y2=1.075
r209 44 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.885
+ $X2=1.765 $Y2=2.885
r210 43 72 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=2.195 $Y2=2.885
r211 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.885
+ $X2=1.84 $Y2=2.885
r212 42 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.775
+ $X2=1.765 $Y2=1.775
r213 41 71 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.775
+ $X2=2.195 $Y2=1.775
r214 41 42 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.775
+ $X2=1.84 $Y2=1.775
r215 38 70 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=2.885
r216 38 40 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r217 35 69 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.7
+ $X2=1.765 $Y2=1.775
r218 35 37 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.765 $Y=1.7
+ $X2=1.765 $Y2=1.075
r219 34 68 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.885
+ $X2=1.335 $Y2=2.885
r220 33 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.885
r221 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.41 $Y2=2.885
r222 32 67 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.775
+ $X2=1.335 $Y2=1.775
r223 31 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.775
+ $X2=1.765 $Y2=1.775
r224 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.775
+ $X2=1.41 $Y2=1.775
r225 28 68 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=2.885
r226 28 30 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r227 25 67 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.7
+ $X2=1.335 $Y2=1.775
r228 25 27 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.335 $Y=1.7
+ $X2=1.335 $Y2=1.075
r229 24 66 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.885
+ $X2=0.905 $Y2=2.885
r230 23 68 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=1.335 $Y2=2.885
r231 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=0.98 $Y2=2.885
r232 22 65 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.775
+ $X2=0.905 $Y2=1.775
r233 21 67 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=1.335 $Y2=1.775
r234 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=0.98 $Y2=1.775
r235 18 66 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=2.885
r236 18 20 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=4.585
r237 15 65 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.775
r238 15 17 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.075
r239 14 64 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.885
+ $X2=0.475 $Y2=2.885
r240 13 66 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.905 $Y2=2.885
r241 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.55 $Y2=2.885
r242 12 63 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.775
+ $X2=0.475 $Y2=1.775
r243 11 65 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.905 $Y2=1.775
r244 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.55 $Y2=1.775
r245 8 64 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=2.885
r246 8 10 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=4.585
r247 7 64 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.885
r248 7 86 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.47
r249 4 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=1.775
r250 4 85 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=2.14
r251 1 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.775
r252 1 3 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__INV_6%Y 1 2 3 4 5 6 19 20 22 24 26 29 30 31 32
+ 33 34 35 41 47 53 55 67 79
c129 35 0 1.33323e-19 $X=2.41 $Y=2.845
c130 34 0 1.33323e-19 $X=2.41 $Y=1.595
c131 33 0 2.66647e-19 $X=1.695 $Y=2.96
c132 31 0 2.66647e-19 $X=1.695 $Y=1.48
c133 20 0 1.33323e-19 $X=0.69 $Y=2.845
c134 19 0 1.33323e-19 $X=0.69 $Y=1.595
r135 86 88 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r136 74 76 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r137 62 64 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r138 53 86 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.41 $Y=2.96
+ $X2=2.41 $Y2=3.455
r139 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.96
+ $X2=2.41 $Y2=2.96
r140 50 79 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.41 $Y=1.48
+ $X2=2.41 $Y2=0.825
r141 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.48
+ $X2=2.41 $Y2=1.48
r142 47 74 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=3.455
r143 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=2.96
r144 44 67 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r145 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r146 41 62 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=3.455
r147 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=2.96
r148 38 55 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=0.825
r149 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.48
r150 35 52 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.845
+ $X2=2.41 $Y2=2.96
r151 34 49 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=1.48
r152 34 35 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.595
+ $X2=2.41 $Y2=2.845
r153 33 46 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.96
+ $X2=1.55 $Y2=2.96
r154 32 52 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.96
+ $X2=2.41 $Y2=2.96
r155 32 33 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.96
+ $X2=1.695 $Y2=2.96
r156 31 43 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.48
+ $X2=1.55 $Y2=1.48
r157 30 49 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=2.41 $Y2=1.48
r158 30 31 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.48
+ $X2=1.695 $Y2=1.48
r159 29 46 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.845
+ $X2=1.55 $Y2=2.96
r160 28 43 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r161 28 29 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.845
r162 27 40 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.96
+ $X2=0.69 $Y2=2.96
r163 26 46 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=1.55 $Y2=2.96
r164 26 27 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=0.835 $Y2=2.96
r165 25 37 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.48
+ $X2=0.69 $Y2=1.48
r166 24 43 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=1.55 $Y2=1.48
r167 24 25 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=0.835 $Y2=1.48
r168 20 40 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.96
r169 20 22 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.2
r170 19 37 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.48
r171 19 22 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=2.2
r172 6 88 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r173 6 86 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r174 5 76 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r175 5 74 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r176 4 64 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r177 4 62 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r178 3 79 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r179 2 67 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r180 1 55 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

