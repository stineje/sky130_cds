magic
tech sky130A
magscale 1 2
timestamp 1638810222
<< nwell >>
rect 75 1340 1020 1341
rect 71 581 1020 1340
<< nmos >>
rect 171 115 201 315
rect 257 115 287 315
rect 329 115 359 315
rect 449 115 479 315
rect 521 115 551 315
rect 607 115 637 315
rect 815 115 845 315
rect 901 115 931 315
<< pmos >>
rect 171 617 201 1217
rect 257 617 287 1217
rect 329 617 359 1217
rect 449 617 479 1217
rect 521 617 551 1217
rect 607 617 637 1217
rect 815 617 845 1217
rect 901 617 931 1217
<< ndiff >>
rect 118 267 171 315
rect 118 131 126 267
rect 160 131 171 267
rect 118 115 171 131
rect 201 267 257 315
rect 201 131 212 267
rect 246 131 257 267
rect 201 115 257 131
rect 287 115 329 315
rect 359 267 449 315
rect 359 131 370 267
rect 438 131 449 267
rect 359 115 449 131
rect 479 115 521 315
rect 551 267 607 315
rect 551 131 562 267
rect 596 131 607 267
rect 551 115 607 131
rect 637 267 690 315
rect 637 131 648 267
rect 682 131 690 267
rect 637 115 690 131
rect 762 267 815 315
rect 762 131 770 267
rect 804 131 815 267
rect 762 115 815 131
rect 845 267 901 315
rect 845 131 856 267
rect 890 131 901 267
rect 845 115 901 131
rect 931 267 984 315
rect 931 131 942 267
rect 976 131 984 267
rect 931 115 984 131
<< pdiff >>
rect 118 1201 171 1217
rect 118 725 126 1201
rect 160 725 171 1201
rect 118 617 171 725
rect 201 1201 257 1217
rect 201 725 212 1201
rect 246 725 257 1201
rect 201 617 257 725
rect 287 617 329 1217
rect 359 1201 449 1217
rect 359 657 370 1201
rect 438 657 449 1201
rect 359 617 449 657
rect 479 617 521 1217
rect 551 1201 607 1217
rect 551 657 562 1201
rect 596 657 607 1201
rect 551 617 607 657
rect 637 1201 690 1217
rect 637 657 648 1201
rect 682 657 690 1201
rect 637 617 690 657
rect 762 1201 815 1217
rect 762 657 770 1201
rect 804 657 815 1201
rect 762 617 815 657
rect 845 1201 901 1217
rect 845 657 856 1201
rect 890 657 901 1201
rect 845 617 901 657
rect 931 1201 984 1217
rect 931 657 942 1201
rect 976 657 984 1201
rect 931 617 984 657
<< ndiffc >>
rect 126 131 160 267
rect 212 131 246 267
rect 370 131 438 267
rect 562 131 596 267
rect 648 131 682 267
rect 770 131 804 267
rect 856 131 890 267
rect 942 131 976 267
<< pdiffc >>
rect 126 725 160 1201
rect 212 725 246 1201
rect 370 657 438 1201
rect 562 657 596 1201
rect 648 657 682 1201
rect 770 657 804 1201
rect 856 657 890 1201
rect 942 657 976 1201
<< psubdiff >>
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
<< nsubdiff >>
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
rect 707 1271 731 1305
rect 765 1271 789 1305
rect 843 1271 867 1305
rect 901 1271 925 1305
<< psubdiffcont >>
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
<< nsubdiffcont >>
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
rect 731 1271 765 1305
rect 867 1271 901 1305
<< poly >>
rect 171 1217 201 1243
rect 257 1217 287 1243
rect 329 1217 359 1243
rect 449 1217 479 1243
rect 521 1217 551 1243
rect 607 1217 637 1243
rect 815 1217 845 1243
rect 901 1217 931 1243
rect 171 595 201 617
rect 161 561 201 595
rect 161 403 191 561
rect 257 518 287 617
rect 329 586 359 617
rect 449 586 479 617
rect 329 570 383 586
rect 329 536 339 570
rect 373 536 383 570
rect 329 520 383 536
rect 425 570 479 586
rect 425 536 435 570
rect 469 536 479 570
rect 425 520 479 536
rect 233 502 287 518
rect 233 468 243 502
rect 277 468 287 502
rect 425 475 455 520
rect 233 452 287 468
rect 161 387 215 403
rect 161 353 171 387
rect 205 353 215 387
rect 161 337 215 353
rect 171 315 201 337
rect 257 315 287 452
rect 329 445 455 475
rect 521 477 551 617
rect 607 586 637 617
rect 815 601 845 617
rect 607 570 678 586
rect 607 556 634 570
rect 618 536 634 556
rect 668 536 678 570
rect 618 520 678 536
rect 805 571 845 601
rect 521 461 575 477
rect 329 315 359 445
rect 521 427 531 461
rect 565 427 575 461
rect 521 411 575 427
rect 425 387 479 403
rect 425 353 435 387
rect 469 353 479 387
rect 425 337 479 353
rect 449 315 479 337
rect 521 315 551 411
rect 618 363 648 520
rect 805 477 835 571
rect 901 477 931 617
rect 780 461 835 477
rect 780 427 790 461
rect 824 427 835 461
rect 780 411 835 427
rect 877 461 931 477
rect 877 427 887 461
rect 921 427 931 461
rect 877 411 931 427
rect 607 333 648 363
rect 805 360 835 411
rect 607 315 637 333
rect 805 330 845 360
rect 815 315 845 330
rect 901 315 931 411
rect 171 89 201 115
rect 257 89 287 115
rect 329 89 359 115
rect 449 89 479 115
rect 521 89 551 115
rect 607 89 637 115
rect 815 89 845 115
rect 901 89 931 115
<< polycont >>
rect 339 536 373 570
rect 435 536 469 570
rect 243 468 277 502
rect 171 353 205 387
rect 634 536 668 570
rect 531 427 565 461
rect 435 353 469 387
rect 790 427 824 461
rect 887 427 921 461
<< locali >>
rect 71 1311 1017 1332
rect 71 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 595 1311
rect 629 1271 731 1311
rect 765 1271 867 1311
rect 901 1271 1017 1311
rect 126 1201 160 1217
rect 103 725 126 791
rect 103 708 160 725
rect 212 1201 246 1271
rect 212 709 246 725
rect 370 1201 438 1217
rect 103 461 137 708
rect 370 654 438 657
rect 103 296 137 427
rect 171 620 438 654
rect 562 1201 596 1271
rect 562 641 596 657
rect 648 1201 682 1217
rect 648 654 682 657
rect 770 1201 804 1217
rect 648 620 736 654
rect 171 387 205 620
rect 435 570 469 586
rect 323 536 339 570
rect 373 536 389 570
rect 243 452 277 468
rect 355 387 389 536
rect 435 535 469 536
rect 634 570 668 586
rect 634 535 668 536
rect 702 461 736 620
rect 770 609 804 657
rect 856 1201 890 1271
rect 856 641 890 657
rect 942 1201 976 1217
rect 976 649 989 666
rect 942 632 989 649
rect 770 570 804 575
rect 770 536 921 570
rect 887 461 921 536
rect 515 427 531 461
rect 565 427 581 461
rect 648 427 736 461
rect 774 427 790 461
rect 824 427 840 461
rect 648 387 682 427
rect 887 387 921 427
rect 205 353 314 387
rect 355 353 435 387
rect 469 353 682 387
rect 171 337 205 353
rect 280 303 314 353
rect 103 267 160 296
rect 103 262 126 267
rect 126 115 160 131
rect 212 267 246 283
rect 280 269 438 303
rect 212 61 246 131
rect 370 267 438 269
rect 370 115 438 131
rect 562 267 596 283
rect 562 61 596 131
rect 648 267 682 353
rect 648 115 682 131
rect 770 353 921 387
rect 770 267 804 353
rect 955 319 989 632
rect 942 285 989 319
rect 770 115 804 131
rect 856 267 890 283
rect 856 61 890 131
rect 942 267 976 285
rect 942 115 976 131
rect 71 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1016 61
rect 71 0 1016 21
<< viali >>
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 595 1305 629 1311
rect 595 1277 629 1305
rect 731 1305 765 1311
rect 731 1277 765 1305
rect 867 1305 901 1311
rect 867 1277 901 1305
rect 103 427 137 461
rect 243 502 277 536
rect 435 501 469 535
rect 634 501 668 535
rect 942 657 976 683
rect 942 649 976 657
rect 770 575 804 609
rect 531 427 565 461
rect 790 427 824 461
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
<< metal1 >>
rect 71 1311 1017 1332
rect 71 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 595 1311
rect 629 1277 731 1311
rect 765 1277 867 1311
rect 901 1277 1017 1311
rect 71 1271 1017 1277
rect 930 683 988 689
rect 907 649 942 683
rect 976 649 988 683
rect 930 643 988 649
rect 758 609 816 615
rect 751 608 770 609
rect 736 576 770 608
rect 751 575 770 576
rect 804 575 816 609
rect 758 569 816 575
rect 231 536 290 542
rect 231 502 243 536
rect 277 502 310 536
rect 423 535 481 541
rect 622 535 680 541
rect 231 496 290 502
rect 423 501 435 535
rect 469 501 634 535
rect 668 501 680 535
rect 423 495 481 501
rect 622 495 680 501
rect 90 461 149 467
rect 90 427 103 461
rect 137 454 149 461
rect 519 461 578 467
rect 519 454 531 461
rect 137 427 531 454
rect 565 458 578 461
rect 778 461 836 467
rect 778 458 790 461
rect 565 430 790 458
rect 565 427 578 430
rect 90 426 578 427
rect 90 421 149 426
rect 519 421 578 426
rect 778 427 790 430
rect 824 427 836 461
rect 778 421 836 427
rect 71 55 1016 61
rect 71 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1016 55
rect 71 0 1016 21
<< labels >>
rlabel metal1 651 518 651 518 1 CK
port 1 n
rlabel metal1 260 518 260 518 1 D
port 2 n
rlabel metal1 959 666 959 666 1 Q
port 3 n
rlabel metal1 788 592 788 592 1 QN
port 4 n
<< end >>
