* File: sky130_osu_sc_18T_ls__inv_2.pxi.spice
* Created: Thu Oct 29 17:36:25 2020
* 
x_PM_SKY130_OSU_SC_18T_LS__INV_2%GND N_GND_M1000_d N_GND_M1002_d N_GND_M1000_b
+ N_GND_c_2_p N_GND_c_9_p N_GND_c_3_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_LS__INV_2%GND
x_PM_SKY130_OSU_SC_18T_LS__INV_2%VDD N_VDD_M1001_s N_VDD_M1003_s N_VDD_M1001_b
+ N_VDD_c_27_p N_VDD_c_33_p N_VDD_c_28_p VDD N_VDD_c_29_p
+ PM_SKY130_OSU_SC_18T_LS__INV_2%VDD
x_PM_SKY130_OSU_SC_18T_LS__INV_2%A N_A_c_47_n N_A_M1000_g N_A_c_51_n N_A_c_65_n
+ N_A_M1001_g N_A_c_52_n N_A_c_53_n N_A_c_54_n N_A_M1002_g N_A_c_70_n
+ N_A_M1003_g N_A_c_58_n N_A_c_59_n N_A_c_60_n N_A_c_61_n N_A_c_62_n A
+ N_A_c_63_n N_A_c_64_n PM_SKY130_OSU_SC_18T_LS__INV_2%A
x_PM_SKY130_OSU_SC_18T_LS__INV_2%Y N_Y_M1000_s N_Y_M1001_d Y N_Y_c_115_n
+ N_Y_c_121_n N_Y_c_122_n N_Y_c_118_n PM_SKY130_OSU_SC_18T_LS__INV_2%Y
cc_1 N_GND_M1000_b N_A_c_47_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.7
cc_2 N_GND_c_2_p N_A_c_47_n 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.7
cc_3 N_GND_c_3_p N_A_c_47_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.7
cc_4 N_GND_c_4_p N_A_c_47_n 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=1.7
cc_5 N_GND_M1000_b N_A_c_51_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.81
cc_6 N_GND_M1000_b N_A_c_52_n 0.0349926f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.775
cc_7 N_GND_M1000_b N_A_c_53_n 0.0263741f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.885
cc_8 N_GND_M1000_b N_A_c_54_n 0.0208613f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.7
cc_9 N_GND_c_9_p N_A_c_54_n 0.00713292f $X=1.12 $Y=0.825 $X2=0.905 $Y2=1.7
cc_10 N_GND_c_3_p N_A_c_54_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.7
cc_11 N_GND_c_4_p N_A_c_54_n 0.00468827f $X=1.02 $Y=0.17 $X2=0.905 $Y2=1.7
cc_12 N_GND_M1000_b N_A_c_58_n 0.0104975f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.775
cc_13 N_GND_M1000_b N_A_c_59_n 0.00422485f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.885
cc_14 N_GND_M1000_b N_A_c_60_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.305
cc_15 N_GND_M1000_b N_A_c_61_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_16 N_GND_M1000_b N_A_c_62_n 0.0348407f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_17 N_GND_M1000_b N_A_c_63_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.33
cc_18 N_GND_M1000_b N_A_c_64_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.14
cc_19 N_GND_M1000_b Y 0.0458015f $X=-0.045 $Y=0 $X2=0.76 $Y2=2.2
cc_20 N_GND_M1000_b N_Y_c_115_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.48
cc_21 N_GND_c_2_p N_Y_c_115_n 0.00125659f $X=0.26 $Y=0.825 $X2=0.69 $Y2=1.48
cc_22 N_GND_c_9_p N_Y_c_115_n 0.00125659f $X=1.12 $Y=0.825 $X2=0.69 $Y2=1.48
cc_23 N_GND_M1000_b N_Y_c_118_n 0.00155118f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_24 N_GND_c_3_p N_Y_c_118_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.825
cc_25 N_GND_c_4_p N_Y_c_118_n 0.00475776f $X=1.02 $Y=0.17 $X2=0.69 $Y2=0.825
cc_26 N_VDD_M1001_b N_A_c_65_n 0.0181616f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=2.96
cc_27 N_VDD_c_27_p N_A_c_65_n 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=2.96
cc_28 N_VDD_c_28_p N_A_c_65_n 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=2.96
cc_29 N_VDD_c_29_p N_A_c_65_n 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=2.96
cc_30 N_VDD_M1001_b N_A_c_53_n 0.00833572f $X=-0.045 $Y=2.905 $X2=0.83 $Y2=2.885
cc_31 N_VDD_M1001_b N_A_c_70_n 0.0207946f $X=-0.045 $Y=2.905 $X2=0.905 $Y2=2.96
cc_32 N_VDD_c_27_p N_A_c_70_n 3.67508e-19 $X=0.26 $Y=4.135 $X2=0.905 $Y2=2.96
cc_33 N_VDD_c_33_p N_A_c_70_n 0.00732698f $X=1.12 $Y=3.455 $X2=0.905 $Y2=2.96
cc_34 N_VDD_c_28_p N_A_c_70_n 0.00610567f $X=1.035 $Y=6.507 $X2=0.905 $Y2=2.96
cc_35 N_VDD_c_29_p N_A_c_70_n 0.00470215f $X=1.02 $Y=6.49 $X2=0.905 $Y2=2.96
cc_36 N_VDD_M1001_b N_A_c_59_n 0.00244597f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.885
cc_37 N_VDD_M1001_s A 0.0162774f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.325
cc_38 N_VDD_c_27_p A 0.00522047f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.325
cc_39 N_VDD_c_33_p A 9.09141e-19 $X=1.12 $Y=3.455 $X2=0.32 $Y2=3.325
cc_40 N_VDD_M1001_s N_A_c_63_n 0.00953431f $X=0.135 $Y=3.085 $X2=0.32 $Y2=3.33
cc_41 N_VDD_M1001_b N_A_c_63_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=3.33
cc_42 N_VDD_c_27_p N_A_c_63_n 0.00252874f $X=0.26 $Y=4.135 $X2=0.32 $Y2=3.33
cc_43 N_VDD_M1001_b N_Y_c_121_n 0.00248543f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_44 N_VDD_M1001_b N_Y_c_122_n 0.00361433f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_45 N_VDD_c_28_p N_Y_c_122_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69 $Y2=2.96
cc_46 N_VDD_c_29_p N_Y_c_122_n 0.00475776f $X=1.02 $Y=6.49 $X2=0.69 $Y2=2.96
cc_47 A N_Y_M1001_d 0.00251573f $X=0.32 $Y=3.325 $X2=0.55 $Y2=3.085
cc_48 N_A_c_47_n Y 0.00150089f $X=0.475 $Y=1.7 $X2=0.76 $Y2=2.2
cc_49 N_A_c_51_n Y 0.00792324f $X=0.475 $Y=2.81 $X2=0.76 $Y2=2.2
cc_50 N_A_c_52_n Y 0.0155521f $X=0.83 $Y=1.775 $X2=0.76 $Y2=2.2
cc_51 N_A_c_53_n Y 0.00371247f $X=0.83 $Y=2.885 $X2=0.76 $Y2=2.2
cc_52 N_A_c_54_n Y 0.00150089f $X=0.905 $Y=1.7 $X2=0.76 $Y2=2.2
cc_53 N_A_c_61_n Y 0.0178517f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_54 N_A_c_62_n Y 0.00610708f $X=0.535 $Y=2.305 $X2=0.76 $Y2=2.2
cc_55 N_A_c_63_n Y 0.0182346f $X=0.32 $Y=3.33 $X2=0.76 $Y2=2.2
cc_56 N_A_c_64_n Y 0.00675469f $X=0.535 $Y=2.14 $X2=0.76 $Y2=2.2
cc_57 N_A_c_47_n N_Y_c_115_n 0.00910659f $X=0.475 $Y=1.7 $X2=0.69 $Y2=1.48
cc_58 N_A_c_54_n N_Y_c_115_n 0.00908049f $X=0.905 $Y=1.7 $X2=0.69 $Y2=1.48
cc_59 N_A_c_62_n N_Y_c_115_n 6.32153e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=1.48
cc_60 N_A_c_65_n N_Y_c_121_n 0.00166042f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.96
cc_61 N_A_c_53_n N_Y_c_121_n 0.00715376f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.96
cc_62 N_A_c_70_n N_Y_c_121_n 0.00524573f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.96
cc_63 N_A_c_59_n N_Y_c_121_n 9.8958e-19 $X=0.475 $Y=2.885 $X2=0.69 $Y2=2.96
cc_64 N_A_c_61_n N_Y_c_121_n 0.00173027f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_65 N_A_c_62_n N_Y_c_121_n 2.98633e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_66 A N_Y_c_121_n 0.00815006f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.96
cc_67 N_A_c_63_n N_Y_c_121_n 0.00637867f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_68 N_A_c_65_n N_Y_c_122_n 0.00199065f $X=0.475 $Y=2.96 $X2=0.69 $Y2=2.96
cc_69 N_A_c_53_n N_Y_c_122_n 0.00839237f $X=0.83 $Y=2.885 $X2=0.69 $Y2=2.96
cc_70 N_A_c_70_n N_Y_c_122_n 0.0035213f $X=0.905 $Y=2.96 $X2=0.69 $Y2=2.96
cc_71 N_A_c_61_n N_Y_c_122_n 0.00165526f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_72 N_A_c_62_n N_Y_c_122_n 2.38128e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_73 A N_Y_c_122_n 0.00938699f $X=0.32 $Y=3.325 $X2=0.69 $Y2=2.96
cc_74 N_A_c_63_n N_Y_c_122_n 0.0226156f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_75 N_A_c_47_n N_Y_c_118_n 0.00231637f $X=0.475 $Y=1.7 $X2=0.69 $Y2=0.825
cc_76 N_A_c_52_n N_Y_c_118_n 0.00256118f $X=0.83 $Y=1.775 $X2=0.69 $Y2=0.825
cc_77 N_A_c_54_n N_Y_c_118_n 0.00231637f $X=0.905 $Y=1.7 $X2=0.69 $Y2=0.825
cc_78 N_A_c_61_n N_Y_c_118_n 0.00110256f $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
