magic
tech sky130A
magscale 1 2
timestamp 1606864602
<< checkpaint >>
rect -1209 -1243 1345 2575
<< nwell >>
rect -9 581 199 1341
<< nmos >>
rect 80 115 110 315
<< pmos >>
rect 80 1017 110 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 163 315
rect 110 131 121 267
rect 155 131 163 267
rect 110 115 163 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 1065 35 1201
rect 69 1065 80 1201
rect 27 1017 80 1065
rect 110 1201 163 1217
rect 110 1065 121 1201
rect 155 1065 163 1201
rect 110 1017 163 1065
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
<< pdiffc >>
rect 35 1065 69 1201
rect 121 1065 155 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1271 85 1305
<< poly >>
rect 80 1217 110 1243
rect 80 315 110 1017
rect 80 80 110 115
<< locali >>
rect 0 1311 198 1332
rect 0 1271 51 1311
rect 85 1271 198 1311
rect 35 1201 69 1271
rect 35 1049 69 1065
rect 121 1201 155 1271
rect 121 1049 155 1065
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 283
rect 121 61 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1311 198 1332
rect 0 1277 51 1311
rect 85 1277 198 1311
rect 0 1271 198 1277
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
