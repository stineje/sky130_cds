* File: sky130_osu_sc_15T_ms__dffsr_l.pex.spice
* Created: Fri Nov 12 14:43:13 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%GND 1 2 3 4 5 6 7 8 9 127 131 133 140
+ 142 152 158 160 170 172 182 184 191 193 203 205 212 238 240
c249 191 0 1.63226e-19 $X=7.47 $Y=0.865
c250 182 0 1.67294e-19 $X=6.52 $Y=0.865
c251 158 0 3.07193e-19 $X=3.02 $Y=0.865
c252 152 0 2.98797e-19 $X=2.5 $Y=0.865
c253 127 0 1.91032e-19 $X=-0.05 $Y=0
r254 238 240 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.855 $Y2=0.152
r255 214 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=0.152
+ $X2=9.71 $Y2=0.152
r256 210 234 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.152
r257 210 212 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.74
r258 206 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.152
+ $X2=8.75 $Y2=0.152
r259 205 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=0.152
+ $X2=9.71 $Y2=0.152
r260 201 233 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.152
r261 201 203 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.74
r262 194 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.152
+ $X2=7.47 $Y2=0.152
r263 193 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.152
+ $X2=8.75 $Y2=0.152
r264 189 232 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.152
r265 189 191 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.865
r266 184 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=0.152
+ $X2=7.47 $Y2=0.152
r267 180 182 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.52 $Y=0.305
+ $X2=6.52 $Y2=0.865
r268 173 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.152
+ $X2=4.77 $Y2=0.152
r269 168 228 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.152
r270 168 170 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.74
r271 160 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.152
+ $X2=4.77 $Y2=0.152
r272 156 158 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.02 $Y=0.305
+ $X2=3.02 $Y2=0.865
r273 155 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.152
+ $X2=2.5 $Y2=0.152
r274 154 155 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=2.935 $Y=0.152
+ $X2=2.585 $Y2=0.152
r275 150 224 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.152
r276 150 152 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.865
r277 143 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0.152
+ $X2=1.22 $Y2=0.152
r278 142 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.152
+ $X2=2.5 $Y2=0.152
r279 138 223 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.152
r280 138 140 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.74
r281 133 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.152
+ $X2=1.22 $Y2=0.152
r282 129 131 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r283 127 240 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=0.19
+ $X2=9.855 $Y2=0.19
r284 127 238 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r285 127 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.52 $Y2=0.305
r286 127 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.435 $Y2=0.152
r287 127 185 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.605 $Y2=0.152
r288 127 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.02 $Y2=0.305
r289 127 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=2.935 $Y2=0.152
r290 127 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.105 $Y2=0.152
r291 127 129 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r292 127 134 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r293 127 214 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.855 $Y=0.152
+ $X2=9.795 $Y2=0.152
r294 127 205 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=9.625 $Y2=0.152
r295 127 206 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.835 $Y2=0.152
r296 127 193 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.665 $Y2=0.152
r297 127 194 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=7.815 $Y=0.152
+ $X2=7.555 $Y2=0.152
r298 127 184 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.385 $Y2=0.152
r299 127 185 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.605 $Y2=0.152
r300 127 172 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.435 $Y2=0.152
r301 127 173 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.855 $Y2=0.152
r302 127 160 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=4.685 $Y2=0.152
r303 127 161 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.105 $Y2=0.152
r304 127 142 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.415 $Y2=0.152
r305 127 143 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.305 $Y2=0.152
r306 127 133 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.135 $Y2=0.152
r307 127 134 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r308 9 212 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.57
+ $Y=0.575 $X2=9.71 $Y2=0.74
r309 8 203 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.61
+ $Y=0.575 $X2=8.75 $Y2=0.74
r310 7 191 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.865
r311 6 182 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.865
r312 5 170 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.575 $X2=4.77 $Y2=0.74
r313 4 158 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.575 $X2=3.02 $Y2=0.865
r314 3 152 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.575 $X2=2.5 $Y2=0.865
r315 2 140 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.575 $X2=1.22 $Y2=0.74
r316 1 131 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%VDD 1 2 3 4 5 6 7 89 93 97 105 109 115
+ 119 127 131 139 143 149 153 161 165 180 184
r144 180 184 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=5.397
+ $X2=9.855 $Y2=5.397
r145 168 180 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=5.36
+ $X2=0.335 $Y2=5.36
r146 165 184 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=5.36
+ $X2=9.855 $Y2=5.36
r147 163 178 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=5.397
+ $X2=9.71 $Y2=5.397
r148 163 165 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.795 $Y=5.397
+ $X2=9.855 $Y2=5.397
r149 159 178 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.71 $Y=5.245
+ $X2=9.71 $Y2=5.397
r150 159 161 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=9.71 $Y=5.245
+ $X2=9.71 $Y2=4.225
r151 156 158 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=8.495 $Y=5.397
+ $X2=9.175 $Y2=5.397
r152 154 177 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=5.397
+ $X2=7.9 $Y2=5.397
r153 154 156 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=7.985 $Y=5.397
+ $X2=8.495 $Y2=5.397
r154 153 178 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=5.397
+ $X2=9.71 $Y2=5.397
r155 153 158 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.625 $Y=5.397
+ $X2=9.175 $Y2=5.397
r156 149 152 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.9 $Y=3.885
+ $X2=7.9 $Y2=4.565
r157 147 177 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=5.245
+ $X2=7.9 $Y2=5.397
r158 147 152 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.9 $Y=5.245
+ $X2=7.9 $Y2=4.565
r159 144 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=5.397
+ $X2=6.52 $Y2=5.397
r160 144 146 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=6.605 $Y=5.397
+ $X2=7.135 $Y2=5.397
r161 143 177 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=5.397
+ $X2=7.9 $Y2=5.397
r162 143 146 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=5.397
+ $X2=7.135 $Y2=5.397
r163 139 142 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.52 $Y=3.205
+ $X2=6.52 $Y2=4.565
r164 137 175 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.52 $Y=5.245
+ $X2=6.52 $Y2=5.397
r165 137 142 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.52 $Y=5.245
+ $X2=6.52 $Y2=4.565
r166 134 136 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=5.397
+ $X2=5.775 $Y2=5.397
r167 132 173 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=5.397
+ $X2=4.77 $Y2=5.397
r168 132 134 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=4.855 $Y=5.397
+ $X2=5.095 $Y2=5.397
r169 131 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=5.397
+ $X2=6.52 $Y2=5.397
r170 131 136 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=6.435 $Y=5.397
+ $X2=5.775 $Y2=5.397
r171 127 130 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.77 $Y=3.545
+ $X2=4.77 $Y2=4.565
r172 125 173 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.77 $Y=5.245
+ $X2=4.77 $Y2=5.397
r173 125 130 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.77 $Y=5.245
+ $X2=4.77 $Y2=4.565
r174 122 124 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=5.397
+ $X2=4.415 $Y2=5.397
r175 120 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=5.397
+ $X2=3.02 $Y2=5.397
r176 120 122 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.105 $Y=5.397
+ $X2=3.735 $Y2=5.397
r177 119 173 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=5.397
+ $X2=4.77 $Y2=5.397
r178 119 124 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.685 $Y=5.397
+ $X2=4.415 $Y2=5.397
r179 115 118 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.02 $Y=3.545
+ $X2=3.02 $Y2=4.565
r180 113 172 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.02 $Y=5.245
+ $X2=3.02 $Y2=5.397
r181 113 118 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.02 $Y=5.245
+ $X2=3.02 $Y2=4.565
r182 110 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=5.397
+ $X2=2.07 $Y2=5.397
r183 110 112 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.155 $Y=5.397
+ $X2=2.375 $Y2=5.397
r184 109 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=5.397
+ $X2=3.02 $Y2=5.397
r185 109 112 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=2.935 $Y=5.397
+ $X2=2.375 $Y2=5.397
r186 105 108 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.07 $Y=3.885
+ $X2=2.07 $Y2=4.565
r187 103 170 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.07 $Y=5.245
+ $X2=2.07 $Y2=5.397
r188 103 108 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.07 $Y=5.245
+ $X2=2.07 $Y2=4.565
r189 100 102 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=5.397
+ $X2=1.695 $Y2=5.397
r190 98 168 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r191 98 100 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.015 $Y2=5.397
r192 97 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=5.397
+ $X2=2.07 $Y2=5.397
r193 97 102 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.985 $Y=5.397
+ $X2=1.695 $Y2=5.397
r194 93 96 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.885
+ $X2=0.26 $Y2=4.565
r195 91 168 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r196 91 96 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.565
r197 89 165 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=9.65 $Y=5.245 $X2=9.855 $Y2=5.33
r198 89 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=5.245 $X2=9.175 $Y2=5.33
r199 89 156 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=5.245 $X2=8.495 $Y2=5.33
r200 89 177 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=5.245 $X2=7.815 $Y2=5.33
r201 89 146 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=5.245 $X2=7.135 $Y2=5.33
r202 89 175 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=5.245 $X2=6.455 $Y2=5.33
r203 89 136 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=5.245 $X2=5.775 $Y2=5.33
r204 89 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=5.245 $X2=5.095 $Y2=5.33
r205 89 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=5.245 $X2=4.415 $Y2=5.33
r206 89 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=5.245 $X2=3.735 $Y2=5.33
r207 89 172 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=5.245 $X2=3.055 $Y2=5.33
r208 89 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=5.245 $X2=2.375 $Y2=5.33
r209 89 102 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=5.245 $X2=1.695 $Y2=5.33
r210 89 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=5.245 $X2=1.015 $Y2=5.33
r211 89 168 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=5.245 $X2=0.335 $Y2=5.33
r212 7 161 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=9.57
+ $Y=3.565 $X2=9.71 $Y2=4.225
r213 6 152 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.825 $X2=7.9 $Y2=4.565
r214 6 149 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.825 $X2=7.9 $Y2=3.885
r215 5 142 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=2.825 $X2=6.52 $Y2=4.565
r216 5 139 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=2.825 $X2=6.52 $Y2=3.205
r217 4 130 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.63
+ $Y=2.825 $X2=4.77 $Y2=4.565
r218 4 127 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=4.63
+ $Y=2.825 $X2=4.77 $Y2=3.545
r219 3 118 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.825 $X2=3.02 $Y2=4.565
r220 3 115 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.825 $X2=3.02 $Y2=3.545
r221 2 108 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.825 $X2=2.07 $Y2=4.565
r222 2 105 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.825 $X2=2.07 $Y2=3.885
r223 1 96 400 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r224 1 93 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%RN 3 5 7 13 15 21
c40 21 0 7.48684e-20 $X=0.325 $Y=3.07
c41 3 0 1.63751e-20 $X=0.475 $Y=0.945
r42 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=3.07
+ $X2=0.325 $Y2=3.07
r43 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=2.045
+ $X2=0.53 $Y2=2.045
r44 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.07
+ $X2=0.32 $Y2=3.07
r45 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.21
+ $X2=0.32 $Y2=2.045
r46 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=2.21 $X2=0.32
+ $Y2=3.07
r47 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=2.045 $X2=0.53 $Y2=2.045
r48 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=2.21
+ $X2=0.53 $Y2=2.045
r49 5 7 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=0.475 $Y=2.21
+ $X2=0.475 $Y2=3.825
r50 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.875
+ $X2=0.53 $Y2=2.045
r51 1 3 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.475 $Y=1.875
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_110_115# 1 3 10 13 15 17 18 20 23 26
+ 29 33 37 40 45 49 54 55 56 62 67 69 72 73 78
c211 78 0 1.95146e-19 $X=8.86 $Y=1.22
c212 73 0 1.63751e-20 $X=1.375 $Y=1.22
c213 62 0 7.48684e-20 $X=0.87 $Y=2.48
r214 73 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.375 $Y=1.22
+ $X2=1.23 $Y2=1.22
r215 72 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.715 $Y=1.22
+ $X2=8.86 $Y2=1.22
r216 72 73 7.06756 $w=1.7e-07 $l=7.34e-06 $layer=MET1_cond $X=8.715 $Y=1.22
+ $X2=1.375 $Y2=1.22
r217 69 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.86 $Y=1.22
+ $X2=8.86 $Y2=1.22
r218 69 71 7.17647 $w=2.55e-07 $l=1.5e-07 $layer=LI1_cond $X=8.86 $Y=1.22
+ $X2=8.86 $Y2=1.37
r219 65 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.22
+ $X2=1.23 $Y2=1.22
r220 65 67 8.63208 $w=2.12e-07 $l=1.5e-07 $layer=LI1_cond $X=1.27 $Y=1.22
+ $X2=1.27 $Y2=1.37
r221 60 62 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.87 $Y2=2.48
r222 57 59 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.87 $Y2=1.37
r223 56 59 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.37
+ $X2=0.87 $Y2=1.37
r224 55 67 2.03271 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.145 $Y=1.37
+ $X2=1.27 $Y2=1.37
r225 55 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.145 $Y=1.37
+ $X2=0.955 $Y2=1.37
r226 54 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.395
+ $X2=0.87 $Y2=2.48
r227 53 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.455
+ $X2=0.87 $Y2=1.37
r228 53 54 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.87 $Y=1.455
+ $X2=0.87 $Y2=2.395
r229 49 51 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=3.205
+ $X2=0.69 $Y2=4.565
r230 47 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.565
+ $X2=0.69 $Y2=2.48
r231 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.69 $Y=2.565
+ $X2=0.69 $Y2=3.205
r232 43 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.285
+ $X2=0.69 $Y2=1.37
r233 43 45 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.69 $Y=1.285
+ $X2=0.69 $Y2=0.865
r234 42 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.86
+ $Y=1.37 $X2=8.86 $Y2=1.37
r235 40 42 12.05 $w=2.4e-07 $l=6e-08 $layer=POLY_cond $X=8.8 $Y=1.37 $X2=8.86
+ $Y2=1.37
r236 35 37 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.545 $Y=2.56
+ $X2=8.8 $Y2=2.56
r237 32 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.37 $X2=1.23 $Y2=1.37
r238 32 33 10.8315 $w=2.67e-07 $l=6e-08 $layer=POLY_cond $X=1.23 $Y=1.37
+ $X2=1.29 $Y2=1.37
r239 27 29 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.29 $Y=2.56
+ $X2=1.425 $Y2=2.56
r240 26 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.8 $Y=2.485
+ $X2=8.8 $Y2=2.56
r241 25 40 13.7767 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=1.535
+ $X2=8.8 $Y2=1.37
r242 25 26 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.8 $Y=1.535
+ $X2=8.8 $Y2=2.485
r243 21 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.545 $Y=2.635
+ $X2=8.545 $Y2=2.56
r244 21 23 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=8.545 $Y=2.635
+ $X2=8.545 $Y2=3.825
r245 18 40 53.2208 $w=2.4e-07 $l=3.37565e-07 $layer=POLY_cond $X=8.535 $Y=1.205
+ $X2=8.8 $Y2=1.37
r246 18 20 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.535 $Y=1.205
+ $X2=8.535 $Y2=0.835
r247 15 33 26.176 $w=2.67e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.435 $Y=1.205
+ $X2=1.29 $Y2=1.37
r248 15 17 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.435 $Y=1.205
+ $X2=1.435 $Y2=0.835
r249 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=2.635
+ $X2=1.425 $Y2=2.56
r250 11 13 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=1.425 $Y=2.635
+ $X2=1.425 $Y2=3.825
r251 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=2.485
+ $X2=1.29 $Y2=2.56
r252 9 33 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.535
+ $X2=1.29 $Y2=1.37
r253 9 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.29 $Y=1.535
+ $X2=1.29 $Y2=2.485
r254 3 51 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.565
r255 3 49 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.205
r256 1 45 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%SN 5 9 13 17 20 21 24 26 31 35 38 43 45
+ 46 51
c172 46 0 2.97185e-19 $X=1.855 $Y=2.7
c173 21 0 1.55885e-19 $X=1.752 $Y=1.945
r174 46 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=2.7
+ $X2=1.71 $Y2=2.7
r175 45 51 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.79 $Y=2.7
+ $X2=7.935 $Y2=2.7
r176 45 46 5.71471 $w=1.7e-07 $l=5.935e-06 $layer=MET1_cond $X=7.79 $Y=2.7
+ $X2=1.855 $Y2=2.7
r177 40 43 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.935 $Y=2.035
+ $X2=8.025 $Y2=2.035
r178 35 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.935 $Y=2.7
+ $X2=7.935 $Y2=2.7
r179 33 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=2.16
+ $X2=7.935 $Y2=2.035
r180 33 35 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.935 $Y=2.16
+ $X2=7.935 $Y2=2.7
r181 31 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=2.7
+ $X2=1.71 $Y2=2.7
r182 29 38 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.195
+ $X2=1.71 $Y2=2.11
r183 29 31 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.71 $Y=2.195
+ $X2=1.71 $Y2=2.7
r184 26 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.025
+ $Y=1.995 $X2=8.025 $Y2=1.995
r185 26 28 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=1.995
+ $X2=8.035 $Y2=2.16
r186 26 27 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=8.035 $Y=1.995
+ $X2=8.035 $Y2=1.83
r187 23 24 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.89 $Y=1.515
+ $X2=1.89 $Y2=1.665
r188 21 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.855 $Y=1.945
+ $X2=1.855 $Y2=1.665
r189 20 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=2.11 $X2=1.71 $Y2=2.11
r190 20 22 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.752 $Y=2.11
+ $X2=1.752 $Y2=2.275
r191 20 21 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.752 $Y=2.11
+ $X2=1.752 $Y2=1.945
r192 17 28 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=8.115 $Y=3.825
+ $X2=8.115 $Y2=2.16
r193 13 27 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=8.045 $Y=0.945
+ $X2=8.045 $Y2=1.83
r194 9 23 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.925 $Y=0.945
+ $X2=1.925 $Y2=1.515
r195 5 22 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=1.855 $Y=3.825
+ $X2=1.855 $Y2=2.275
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_432_468# 1 3 11 15 18 24 25 26 27 28
+ 30 33 37 42
c90 42 0 1.71621e-19 $X=3.887 $Y=1.155
c91 25 0 1.29912e-19 $X=3.71 $Y=1.505
c92 18 0 1.52962e-19 $X=2.295 $Y=2.505
c93 15 0 1.44224e-19 $X=2.285 $Y=3.825
c94 11 0 1.44224e-19 $X=2.285 $Y=0.945
r95 41 42 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.887 $Y=0.985
+ $X2=3.887 $Y2=1.155
r96 37 39 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=3.895 $Y=3.205
+ $X2=3.895 $Y2=4.565
r97 35 37 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=3.895 $Y=3.115
+ $X2=3.895 $Y2=3.205
r98 33 41 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.895 $Y=0.865
+ $X2=3.895 $Y2=0.985
r99 30 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.795 $Y=1.42
+ $X2=3.795 $Y2=1.155
r100 27 35 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=3.725 $Y=2.925
+ $X2=3.895 $Y2=3.115
r101 27 28 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=3.725 $Y=2.925
+ $X2=2.38 $Y2=2.925
r102 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=1.505
+ $X2=3.795 $Y2=1.42
r103 25 26 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.71 $Y=1.505
+ $X2=2.38 $Y2=1.505
r104 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=2.84
+ $X2=2.38 $Y2=2.925
r105 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.295 $Y=2.84
+ $X2=2.295 $Y2=2.505
r106 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=1.59
+ $X2=2.38 $Y2=1.505
r107 21 24 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.295 $Y=1.59
+ $X2=2.295 $Y2=2.505
r108 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=2.505 $X2=2.295 $Y2=2.505
r109 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.505
+ $X2=2.295 $Y2=2.67
r110 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.505
+ $X2=2.295 $Y2=2.34
r111 15 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=2.285 $Y=3.825
+ $X2=2.285 $Y2=2.67
r112 11 19 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=2.285 $Y=0.945
+ $X2=2.285 $Y2=2.34
r113 3 39 240 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=3.67
+ $Y=2.825 $X2=3.895 $Y2=4.565
r114 3 37 240 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=2 $X=3.67
+ $Y=2.825 $X2=3.895 $Y2=3.205
r115 1 33 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.575 $X2=3.895 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%D 3 7 10 14 19
c39 19 0 1.41836e-19 $X=3.295 $Y=1.96
c40 10 0 1.12321e-19 $X=3.295 $Y=1.96
r41 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.295 $Y=1.96
+ $X2=3.295 $Y2=1.96
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.96 $X2=3.295 $Y2=1.96
r43 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.96
+ $X2=3.295 $Y2=2.125
r44 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.96
+ $X2=3.295 $Y2=1.795
r45 7 12 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=3.235 $Y=3.825
+ $X2=3.235 $Y2=2.125
r46 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.235 $Y=0.945
+ $X2=3.235 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c233 55 0 6.79641e-20 $X=5.49 $Y=2.33
c234 48 0 1.98654e-19 $X=4.135 $Y=1.59
c235 44 0 1.86602e-19 $X=4.05 $Y=2.33
c236 30 0 1.29912e-19 $X=4.135 $Y=1.425
c237 25 0 1.41836e-19 $X=3.655 $Y=2.505
r238 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.03 $Y=2.33
+ $X2=5.885 $Y2=2.33
r239 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.735 $Y=2.33
+ $X2=6.88 $Y2=2.33
r240 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.735 $Y=2.33
+ $X2=6.03 $Y2=2.33
r241 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.8 $Y=2.33
+ $X2=3.655 $Y2=2.33
r242 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.74 $Y=2.33
+ $X2=5.885 $Y2=2.33
r243 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.74 $Y=2.33
+ $X2=3.8 $Y2=2.33
r244 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=2.33
+ $X2=5.885 $Y2=2.33
r245 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.885 $Y=2.33
+ $X2=5.885 $Y2=2.505
r246 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.655 $Y=2.33
+ $X2=3.655 $Y2=2.33
r247 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.655 $Y=2.33
+ $X2=3.655 $Y2=2.505
r248 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.88 $Y=2.33
+ $X2=6.88 $Y2=2.33
r249 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.88 $Y=2.33
+ $X2=6.88 $Y2=2.505
r250 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.33
+ $X2=5.885 $Y2=2.33
r251 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.8 $Y=2.33
+ $X2=5.49 $Y2=2.33
r252 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.405 $Y=2.245
+ $X2=5.49 $Y2=2.33
r253 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.405 $Y=2.245
+ $X2=5.405 $Y2=1.59
r254 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.135 $Y=2.245
+ $X2=4.135 $Y2=1.59
r255 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=2.33
+ $X2=3.655 $Y2=2.33
r256 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.05 $Y=2.33
+ $X2=4.135 $Y2=2.245
r257 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.05 $Y=2.33
+ $X2=3.74 $Y2=2.33
r258 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=2.505 $X2=6.88 $Y2=2.505
r259 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.762 $Y=1.425
+ $X2=6.762 $Y2=1.575
r260 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=2.505 $X2=5.885 $Y2=2.505
r261 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=2.505
+ $X2=5.885 $Y2=2.67
r262 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.59 $X2=5.405 $Y2=1.59
r263 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.59
+ $X2=5.405 $Y2=1.425
r264 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.59 $X2=4.135 $Y2=1.59
r265 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.59
+ $X2=4.135 $Y2=1.425
r266 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=2.505 $X2=3.655 $Y2=2.505
r267 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=2.505
+ $X2=3.655 $Y2=2.67
r268 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.79 $Y=2.34
+ $X2=6.837 $Y2=2.505
r269 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.79 $Y=2.34
+ $X2=6.79 $Y2=1.575
r270 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.735 $Y=2.67
+ $X2=6.837 $Y2=2.505
r271 18 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=6.735 $Y=2.67
+ $X2=6.735 $Y2=3.825
r272 17 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.735 $Y=0.945
+ $X2=6.735 $Y2=1.425
r273 13 39 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=5.945 $Y=3.825
+ $X2=5.945 $Y2=2.67
r274 10 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.345 $Y=0.945
+ $X2=5.345 $Y2=1.425
r275 7 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.195 $Y=0.945
+ $X2=4.195 $Y2=1.425
r276 3 27 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=3.595 $Y=3.825
+ $X2=3.595 $Y2=2.67
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_217_565# 1 3 11 15 17 18 21 22 27 31
+ 35 39 40 43 49 54 55 56 61
c164 56 0 1.44224e-19 $X=1.855 $Y=1.59
c165 55 0 2.71143e-19 $X=4.49 $Y=1.59
c166 49 0 1.5821e-19 $X=4.725 $Y=2.505
c167 43 0 3.19111e-19 $X=1.71 $Y=0.865
c168 31 0 6.36774e-20 $X=4.985 $Y=3.825
c169 22 0 1.86602e-19 $X=4.63 $Y=2.505
c170 21 0 6.79641e-20 $X=4.91 $Y=2.505
c171 15 0 6.36774e-20 $X=4.555 $Y=3.825
r172 56 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.59
+ $X2=1.71 $Y2=1.59
r173 55 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.49 $Y=1.59
+ $X2=4.635 $Y2=1.59
r174 55 56 2.53719 $w=1.7e-07 $l=2.635e-06 $layer=MET1_cond $X=4.49 $Y=1.59
+ $X2=1.855 $Y2=1.59
r175 52 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.59
+ $X2=4.635 $Y2=1.59
r176 52 54 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=4.635 $Y=1.55
+ $X2=4.725 $Y2=1.55
r177 47 54 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.725 $Y=1.675
+ $X2=4.725 $Y2=1.55
r178 47 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.725 $Y=1.675
+ $X2=4.725 $Y2=2.505
r179 46 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.59
+ $X2=1.71 $Y2=1.59
r180 43 46 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.71 $Y=0.865
+ $X2=1.71 $Y2=1.59
r181 41 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.675
+ $X2=1.71 $Y2=1.59
r182 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=1.76
+ $X2=1.71 $Y2=1.675
r183 39 40 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.625 $Y=1.76
+ $X2=1.295 $Y2=1.76
r184 35 37 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.21 $Y=3.545
+ $X2=1.21 $Y2=4.565
r185 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.845
+ $X2=1.295 $Y2=1.76
r186 33 35 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.21 $Y=1.845
+ $X2=1.21 $Y2=3.545
r187 29 31 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=4.985 $Y=2.64
+ $X2=4.985 $Y2=3.825
r188 25 27 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.985 $Y=1.455
+ $X2=4.985 $Y2=0.945
r189 24 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=2.505 $X2=4.725 $Y2=2.505
r190 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=2.505
+ $X2=4.725 $Y2=2.505
r191 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=2.505
+ $X2=4.985 $Y2=2.64
r192 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=2.505
+ $X2=4.725 $Y2=2.505
r193 20 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=1.59 $X2=4.725 $Y2=1.59
r194 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=1.59
+ $X2=4.725 $Y2=1.59
r195 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=1.59
+ $X2=4.985 $Y2=1.455
r196 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=1.59
+ $X2=4.725 $Y2=1.59
r197 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.64
+ $X2=4.63 $Y2=2.505
r198 13 15 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=4.555 $Y=2.64
+ $X2=4.555 $Y2=3.825
r199 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.455
+ $X2=4.63 $Y2=1.59
r200 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.555 $Y=1.455
+ $X2=4.555 $Y2=0.945
r201 3 37 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.825 $X2=1.21 $Y2=4.565
r202 3 35 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.825 $X2=1.21 $Y2=3.545
r203 1 43 182 $w=1.7e-07 $l=3.76962e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.575 $X2=1.71 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_704_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c191 35 0 1.98654e-19 $X=3.715 $Y=1.5
c192 18 0 1.12321e-19 $X=4.195 $Y=3.825
r193 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=2.925
+ $X2=7.22 $Y2=2.925
r194 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=1.93
+ $X2=7.22 $Y2=1.93
r195 60 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.84
+ $X2=7.22 $Y2=2.925
r196 59 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.015
+ $X2=7.22 $Y2=1.93
r197 59 60 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=7.22 $Y=2.015
+ $X2=7.22 $Y2=2.84
r198 55 57 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.95 $Y=3.205
+ $X2=6.95 $Y2=4.565
r199 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=3.01
+ $X2=6.95 $Y2=2.925
r200 53 55 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.95 $Y=3.01
+ $X2=6.95 $Y2=3.205
r201 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.845
+ $X2=6.95 $Y2=1.93
r202 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.675
+ $X2=6.95 $Y2=1.59
r203 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.95 $Y=1.675
+ $X2=6.95 $Y2=1.845
r204 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.505
+ $X2=6.95 $Y2=1.59
r205 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.95 $Y=1.505
+ $X2=6.95 $Y2=0.865
r206 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=1.59
+ $X2=6.95 $Y2=1.59
r207 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.865 $Y=1.59
+ $X2=5.885 $Y2=1.59
r208 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=1.59 $X2=5.885 $Y2=1.59
r209 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.59
+ $X2=5.885 $Y2=1.755
r210 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.59
+ $X2=5.885 $Y2=1.425
r211 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.595 $Y=1.5
+ $X2=3.715 $Y2=1.5
r212 32 41 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.945 $Y=0.945
+ $X2=5.945 $Y2=1.425
r213 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.825 $Y=1.965
+ $X2=5.825 $Y2=1.755
r214 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=2.04
+ $X2=5.345 $Y2=2.04
r215 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.75 $Y=2.04
+ $X2=5.825 $Y2=1.965
r216 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.75 $Y=2.04
+ $X2=5.42 $Y2=2.04
r217 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.345 $Y=2.115
+ $X2=5.345 $Y2=2.04
r218 22 24 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=5.345 $Y=2.115
+ $X2=5.345 $Y2=3.825
r219 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=2.04
+ $X2=4.195 $Y2=2.04
r220 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=2.04
+ $X2=5.345 $Y2=2.04
r221 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.27 $Y=2.04 $X2=4.27
+ $Y2=2.04
r222 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=2.115
+ $X2=4.195 $Y2=2.04
r223 16 18 876.83 $w=1.5e-07 $l=1.71e-06 $layer=POLY_cond $X=4.195 $Y=2.115
+ $X2=4.195 $Y2=3.825
r224 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=2.04
+ $X2=4.195 $Y2=2.04
r225 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.12 $Y=2.04
+ $X2=3.79 $Y2=2.04
r226 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=1.965
+ $X2=3.79 $Y2=2.04
r227 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.715 $Y=1.575
+ $X2=3.715 $Y2=1.5
r228 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.715 $Y=1.575
+ $X2=3.715 $Y2=1.965
r229 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.425
+ $X2=3.595 $Y2=1.5
r230 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.595 $Y=1.425
+ $X2=3.595 $Y2=0.945
r231 3 57 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=2.825 $X2=6.95 $Y2=4.565
r232 3 55 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=2.825 $X2=6.95 $Y2=3.205
r233 1 49 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.575 $X2=6.95 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_1246_89# 1 3 11 15 23 27 30 34 35 38
+ 39 40 42 48 52 56 58 63 64 69
c175 58 0 1.95146e-19 $X=9.38 $Y=1.93
c176 48 0 1.63226e-19 $X=8.26 $Y=0.865
c177 39 0 8.77106e-20 $X=9.47 $Y=2.595
c178 34 0 2.20654e-19 $X=9.38 $Y=1.93
r179 64 66 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.51 $Y=1.93
+ $X2=6.365 $Y2=1.93
r180 63 69 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.235 $Y=1.93
+ $X2=9.38 $Y2=1.93
r181 63 64 2.62385 $w=1.7e-07 $l=2.725e-06 $layer=MET1_cond $X=9.235 $Y=1.93
+ $X2=6.51 $Y2=1.93
r182 58 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.38 $Y=1.93
+ $X2=9.38 $Y2=1.93
r183 56 58 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.845 $Y=1.93
+ $X2=9.38 $Y2=1.93
r184 52 54 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.76 $Y=3.545
+ $X2=8.76 $Y2=4.565
r185 50 56 5.37722 $w=2.41e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=2.015
+ $X2=8.845 $Y2=1.93
r186 50 52 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=8.76 $Y=2.015
+ $X2=8.76 $Y2=3.545
r187 46 50 25.3112 $w=2.41e-07 $l=6.89202e-07 $layer=LI1_cond $X=8.26 $Y=1.565
+ $X2=8.76 $Y2=2.015
r188 46 48 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.26 $Y=1.565
+ $X2=8.26 $Y2=0.865
r189 42 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.365 $Y=1.93
+ $X2=6.365 $Y2=1.93
r190 39 40 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=2.595
+ $X2=9.47 $Y2=2.745
r191 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=1.39 $X2=9.47
+ $Y2=1.54
r192 36 39 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.445 $Y=2.095
+ $X2=9.445 $Y2=2.595
r193 35 38 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.445 $Y=1.765
+ $X2=9.445 $Y2=1.54
r194 34 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.38
+ $Y=1.93 $X2=9.38 $Y2=1.93
r195 34 36 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=1.93
+ $X2=9.382 $Y2=2.095
r196 34 35 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=1.93
+ $X2=9.382 $Y2=1.765
r197 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=1.93 $X2=6.365 $Y2=1.93
r198 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.93
+ $X2=6.365 $Y2=2.095
r199 30 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.93
+ $X2=6.365 $Y2=1.765
r200 27 40 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=9.495 $Y=4.195
+ $X2=9.495 $Y2=2.745
r201 23 37 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=9.495 $Y=0.835
+ $X2=9.495 $Y2=1.39
r202 15 32 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=6.305 $Y=3.825
+ $X2=6.305 $Y2=2.095
r203 11 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.305 $Y=0.945
+ $X2=6.305 $Y2=1.765
r204 3 54 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=8.62
+ $Y=2.825 $X2=8.76 $Y2=4.565
r205 3 52 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=8.62
+ $Y=2.825 $X2=8.76 $Y2=3.545
r206 1 48 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=8.12
+ $Y=0.575 $X2=8.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_1084_115# 1 3 10 11 13 16 20 26 31 32
+ 33 34 35 38 42 47 52 53 58
c157 53 0 1.5821e-19 $X=5.21 $Y=1.59
c158 32 0 1.67294e-19 $X=5.475 $Y=1.17
c159 31 0 1.57671e-19 $X=5.065 $Y=1.59
c160 16 0 6.36774e-20 $X=7.685 $Y=3.825
r161 53 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.21 $Y=1.59
+ $X2=5.065 $Y2=1.59
r162 52 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=1.59
+ $X2=7.595 $Y2=1.59
r163 52 53 2.15686 $w=1.7e-07 $l=2.24e-06 $layer=MET1_cond $X=7.45 $Y=1.59
+ $X2=5.21 $Y2=1.59
r164 47 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=1.59
+ $X2=7.595 $Y2=1.59
r165 47 50 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.595 $Y=1.59
+ $X2=7.595 $Y2=2.505
r166 42 44 34.5733 $w=3.38e-07 $l=1.02e-06 $layer=LI1_cond $X=5.645 $Y=3.545
+ $X2=5.645 $Y2=4.565
r167 40 42 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=5.645 $Y=3.01
+ $X2=5.645 $Y2=3.545
r168 36 38 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=5.645 $Y=1.085
+ $X2=5.645 $Y2=0.865
r169 34 40 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=2.925
+ $X2=5.645 $Y2=3.01
r170 34 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=2.925
+ $X2=5.15 $Y2=2.925
r171 32 36 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=1.17
+ $X2=5.645 $Y2=1.085
r172 32 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=1.17
+ $X2=5.15 $Y2=1.17
r173 31 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.065 $Y=1.59
+ $X2=5.065 $Y2=1.59
r174 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=2.84
+ $X2=5.15 $Y2=2.925
r175 29 31 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.065 $Y=2.84
+ $X2=5.065 $Y2=1.59
r176 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=1.255
+ $X2=5.15 $Y2=1.17
r177 28 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.065 $Y=1.255
+ $X2=5.065 $Y2=1.59
r178 25 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=2.505 $X2=7.595 $Y2=2.505
r179 25 26 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=2.505
+ $X2=7.685 $Y2=2.505
r180 22 25 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=2.505
+ $X2=7.595 $Y2=2.505
r181 18 20 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=7.505 $Y=1.51
+ $X2=7.685 $Y2=1.51
r182 14 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.685 $Y=2.64
+ $X2=7.685 $Y2=2.505
r183 14 16 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=7.685 $Y=2.64
+ $X2=7.685 $Y2=3.825
r184 11 20 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.685 $Y=1.43
+ $X2=7.685 $Y2=1.51
r185 11 13 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.685 $Y=1.43
+ $X2=7.685 $Y2=0.945
r186 10 22 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.505 $Y=2.37
+ $X2=7.505 $Y2=2.505
r187 9 18 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.505 $Y=1.59
+ $X2=7.505 $Y2=1.51
r188 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.505 $Y=1.59
+ $X2=7.505 $Y2=2.37
r189 3 44 300 $w=1.7e-07 $l=1.84908e-06 $layer=licon1_PDIFF $count=2 $X=5.42
+ $Y=2.825 $X2=5.645 $Y2=4.565
r190 3 42 300 $w=1.7e-07 $l=8.24864e-07 $layer=licon1_PDIFF $count=2 $X=5.42
+ $Y=2.825 $X2=5.645 $Y2=3.545
r191 1 38 182 $w=1.7e-07 $l=3.86458e-07 $layer=licon1_NDIFF $count=1 $X=5.42
+ $Y=0.575 $X2=5.645 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c86 42 0 8.77106e-20 $X=9.285 $Y=2.7
c87 33 0 9.99996e-20 $X=9.78 $Y=2.505
c88 31 0 1.20654e-19 $X=9.78 $Y=1.59
r89 40 42 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=9.28 $Y=2.7
+ $X2=9.285 $Y2=2.7
r90 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.865 $Y=2.42
+ $X2=9.865 $Y2=2.135
r91 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.865 $Y=1.675
+ $X2=9.865 $Y2=2.135
r92 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=2.505
+ $X2=9.865 $Y2=2.42
r93 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=2.505
+ $X2=9.365 $Y2=2.505
r94 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.59
+ $X2=9.865 $Y2=1.675
r95 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=1.59
+ $X2=9.365 $Y2=1.59
r96 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=2.7 $X2=9.28
+ $Y2=2.7
r97 27 29 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=9.28 $Y=2.7
+ $X2=9.28 $Y2=4.225
r98 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=2.59
+ $X2=9.365 $Y2=2.505
r99 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.28 $Y=2.59
+ $X2=9.28 $Y2=2.7
r100 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=1.505
+ $X2=9.365 $Y2=1.59
r101 21 23 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=9.28 $Y=1.505
+ $X2=9.28 $Y2=0.74
r102 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.865
+ $Y=2.135 $X2=9.865 $Y2=2.135
r103 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=2.135
+ $X2=9.865 $Y2=2.3
r104 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=2.135
+ $X2=9.865 $Y2=1.97
r105 15 20 971.691 $w=1.5e-07 $l=1.895e-06 $layer=POLY_cond $X=9.925 $Y=4.195
+ $X2=9.925 $Y2=2.3
r106 11 19 581.989 $w=1.5e-07 $l=1.135e-06 $layer=POLY_cond $X=9.925 $Y=0.835
+ $X2=9.925 $Y2=1.97
r107 3 29 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=9.155
+ $Y=3.565 $X2=9.28 $Y2=4.225
r108 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.575 $X2=9.28 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_300_565# 1 2 11 15 16 19
r20 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.5 $Y=3.545
+ $X2=2.5 $Y2=4.565
r21 17 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.5 $Y=3.455 $X2=2.5
+ $Y2=3.545
r22 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=3.37
+ $X2=2.5 $Y2=3.455
r23 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.415 $Y=3.37
+ $X2=1.725 $Y2=3.37
r24 11 13 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.64 $Y=3.545
+ $X2=1.64 $Y2=4.565
r25 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.455
+ $X2=1.725 $Y2=3.37
r26 9 11 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.64 $Y=3.455 $X2=1.64
+ $Y2=3.545
r27 2 21 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=2.825 $X2=2.5 $Y2=4.565
r28 2 19 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=2.825 $X2=2.5 $Y2=3.545
r29 1 13 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.825 $X2=1.64 $Y2=4.565
r30 1 11 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.825 $X2=1.64 $Y2=3.545
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%A_1469_565# 1 2 11 15 16 19
r19 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.33 $Y=3.545
+ $X2=8.33 $Y2=4.565
r20 17 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.33 $Y=3.455 $X2=8.33
+ $Y2=3.545
r21 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.245 $Y=3.37
+ $X2=8.33 $Y2=3.455
r22 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.245 $Y=3.37
+ $X2=7.555 $Y2=3.37
r23 11 13 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.47 $Y=3.545
+ $X2=7.47 $Y2=4.565
r24 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=3.455
+ $X2=7.555 $Y2=3.37
r25 9 11 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.47 $Y=3.455 $X2=7.47
+ $Y2=3.545
r26 2 21 300 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=2.825 $X2=8.33 $Y2=4.565
r27 2 19 300 $w=1.7e-07 $l=7.86893e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=2.825 $X2=8.33 $Y2=3.545
r28 1 13 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=2.825 $X2=7.47 $Y2=4.565
r29 1 11 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=2.825 $X2=7.47 $Y2=3.545
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__DFFSR_L%Q 1 3 11 15 18 21 25 28
r22 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=3.027
+ $X2=10.255 $Y2=3.027
r23 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.135 $Y=3.07
+ $X2=10.135 $Y2=3.07
r24 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=10.135 $Y=3.027
+ $X2=10.14 $Y2=3.027
r25 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=1.255
+ $X2=10.255 $Y2=1.255
r26 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=10.255 $Y=2.9
+ $X2=10.255 $Y2=3.027
r27 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=1.34
+ $X2=10.255 $Y2=1.255
r28 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=10.255 $Y=1.34
+ $X2=10.255 $Y2=2.9
r29 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.14 $Y=3.155
+ $X2=10.14 $Y2=3.027
r30 13 15 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=10.14 $Y=3.155
+ $X2=10.14 $Y2=4.225
r31 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=1.17
+ $X2=10.14 $Y2=1.255
r32 9 11 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.14 $Y=1.17
+ $X2=10.14 $Y2=0.74
r33 3 15 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=10
+ $Y=3.565 $X2=10.14 $Y2=4.225
r34 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=10
+ $Y=0.575 $X2=10.14 $Y2=0.74
.ends

