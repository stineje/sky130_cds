* File: sky130_osu_sc_12T_ls__mux2_1.pex.spice
* Created: Fri Nov 12 15:38:30 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%GND 1 29 33 54 56
r36 54 56 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r37 31 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r38 29 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r39 29 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r40 29 31 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r41 29 35 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r42 29 35 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r43 1 33 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%VDD 1 9 13 17 21
r30 21 24 0.00227273 $w=2.75e-06 $l=5e-08 $layer=MET1_cond $X=1.375 $Y=4.2
+ $X2=1.375 $Y2=4.25
r31 17 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.38 $Y=4.25
+ $X2=2.38 $Y2=4.25
r32 15 17 76.8925 $w=3.03e-07 $l=2.035e-06 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=2.38 $Y2=4.287
r33 11 15 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.345 $Y2=4.287
r34 11 13 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135 $X2=0.26
+ $Y2=3.635
r35 9 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r36 1 13 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%A_110_115# 1 3 9 11 15 19 24 28 31 34 37
+ 44 49
c69 9 0 3.63536e-20 $X=1.35 $Y=1.31
r70 46 49 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=2.21
+ $X2=0.925 $Y2=2.21
r71 41 44 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=1.37
+ $X2=0.925 $Y2=1.37
r72 37 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r73 35 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.375
+ $X2=0.69 $Y2=2.21
r74 35 37 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=0.69 $Y=2.375
+ $X2=0.69 $Y2=2.955
r75 34 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=2.045
+ $X2=0.69 $Y2=2.21
r76 33 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.535
+ $X2=0.69 $Y2=1.37
r77 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.69 $Y=1.535
+ $X2=0.69 $Y2=2.045
r78 29 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.205
+ $X2=0.69 $Y2=1.37
r79 29 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=1.205
+ $X2=0.69 $Y2=0.755
r80 26 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.21 $X2=0.925 $Y2=2.21
r81 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.21
+ $X2=1.09 $Y2=2.21
r82 22 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.37 $X2=0.925 $Y2=1.37
r83 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.37
+ $X2=1.09 $Y2=1.37
r84 17 19 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.855 $Y=2.225
+ $X2=1.855 $Y2=3.235
r85 13 15 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.425 $Y=1.235
+ $X2=1.425 $Y2=0.835
r86 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=2.15
+ $X2=1.855 $Y2=2.225
r87 11 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.78 $Y=2.15
+ $X2=1.09 $Y2=2.15
r88 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=1.31
+ $X2=1.425 $Y2=1.235
r89 9 24 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.35 $Y=1.31 $X2=1.09
+ $Y2=1.31
r90 3 39 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r91 3 37 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r92 1 31 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%S0 3 8 9 11 12 13 15 18 24 26 32
c65 8 0 1.8854e-20 $X=0.475 $Y=3.235
r66 29 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.85
+ $X2=0.27 $Y2=2.85
r67 26 29 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.27 $Y=1.825
+ $X2=0.27 $Y2=2.85
r68 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.825
+ $X2=0.55 $Y2=1.825
r69 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.825 $X2=0.27 $Y2=1.825
r70 21 23 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.825
+ $X2=0.475 $Y2=1.825
r71 16 18 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.855 $Y=1.715
+ $X2=1.855 $Y2=0.835
r72 13 15 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.425 $Y=3.94
+ $X2=1.425 $Y2=3.235
r73 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=4.015
+ $X2=1.425 $Y2=3.94
r74 11 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.35 $Y=4.015 $X2=0.55
+ $Y2=4.015
r75 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=1.79
+ $X2=1.855 $Y2=1.715
r76 9 24 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.78 $Y=1.79
+ $X2=0.55 $Y2=1.79
r77 6 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=3.94
+ $X2=0.55 $Y2=4.015
r78 6 8 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=3.94 $X2=0.475
+ $Y2=3.235
r79 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=1.825
r80 5 8 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=3.235
r81 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.66
+ $X2=0.475 $Y2=1.825
r82 1 3 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=0.475 $Y=1.66
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%A0 1 3 11 15 22 24 26 28
c42 28 0 1.8854e-20 $X=1.265 $Y=2.48
r43 25 26 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=2.635
+ $X2=1.237 $Y2=2.805
r44 23 24 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.237 $Y=0.855
+ $X2=1.237 $Y2=1.025
r45 22 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.265 $Y=2.48
+ $X2=1.265 $Y2=2.48
r46 22 25 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.265 $Y=2.48
+ $X2=1.265 $Y2=2.635
r47 22 24 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=1.265 $Y=2.48
+ $X2=1.265 $Y2=1.025
r48 15 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.21 $Y=2.955
+ $X2=1.21 $Y2=3.635
r49 15 26 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.21 $Y=2.955
+ $X2=1.21 $Y2=2.805
r50 11 23 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.21 $Y=0.755 $X2=1.21
+ $Y2=0.855
r51 3 17 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=2.605 $X2=1.21 $Y2=3.635
r52 3 15 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=2.605 $X2=1.21 $Y2=2.955
r53 1 11 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%Y 1 3 10 16 24 26 29
c37 29 0 3.63536e-20 $X=1.64 $Y=1.74
r38 24 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=1.625
+ $X2=1.64 $Y2=1.74
r39 23 26 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.64 $Y=1.115
+ $X2=1.64 $Y2=1
r40 23 24 0.49107 $w=1.7e-07 $l=5.1e-07 $layer=MET1_cond $X=1.64 $Y=1.115
+ $X2=1.64 $Y2=1.625
r41 19 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.64 $Y=2.955
+ $X2=1.64 $Y2=3.635
r42 16 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.74
+ $X2=1.64 $Y2=1.74
r43 16 19 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=1.64 $Y=1.74
+ $X2=1.64 $Y2=2.955
r44 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1 $X2=1.64
+ $Y2=1
r45 10 13 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.64 $Y=0.755
+ $X2=1.64 $Y2=1
r46 3 21 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=2.605 $X2=1.64 $Y2=3.635
r47 3 19 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=2.605 $X2=1.64 $Y2=2.955
r48 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.5 $Y=0.575
+ $X2=1.64 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__MUX2_1%A1 1 3 10 20
r17 15 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.07 $Y=2.955
+ $X2=2.07 $Y2=3.635
r18 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.11
+ $X2=2.07 $Y2=2.11
r19 13 15 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.07 $Y=2.11
+ $X2=2.07 $Y2=2.955
r20 10 13 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=2.07 $Y=0.755
+ $X2=2.07 $Y2=2.11
r21 3 17 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.605 $X2=2.07 $Y2=3.635
r22 3 15 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.605 $X2=2.07 $Y2=2.955
r23 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.93 $Y=0.575
+ $X2=2.07 $Y2=0.755
.ends

