* File: sky130_osu_sc_18T_hs__aoi21_l.pxi.spice
* Created: Fri Nov 12 13:47:32 2021
* 
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%GND N_GND_M1004_s N_GND_M1005_d N_GND_M1004_b
+ N_GND_c_3_p N_GND_c_4_p N_GND_c_20_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_18T_HS__AOI21_L%GND
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%VDD N_VDD_M1003_d N_VDD_M1003_b N_VDD_c_42_p
+ N_VDD_c_43_p N_VDD_c_49_p VDD N_VDD_c_44_p
+ PM_SKY130_OSU_SC_18T_HS__AOI21_L%VDD
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%A0 N_A0_c_67_n N_A0_c_68_n N_A0_M1004_g
+ N_A0_M1003_g N_A0_c_72_n N_A0_c_74_n N_A0_c_75_n A0
+ PM_SKY130_OSU_SC_18T_HS__AOI21_L%A0
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%A1 N_A1_M1002_g N_A1_M1000_g N_A1_c_108_n
+ N_A1_c_109_n N_A1_c_110_n A1 PM_SKY130_OSU_SC_18T_HS__AOI21_L%A1
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%B0 N_B0_M1005_g N_B0_M1001_g N_B0_c_159_n
+ N_B0_c_160_n N_B0_c_161_n N_B0_c_163_n N_B0_c_164_n N_B0_c_165_n B0
+ PM_SKY130_OSU_SC_18T_HS__AOI21_L%B0
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%A_27_617# N_A_27_617#_M1003_s
+ N_A_27_617#_M1000_d N_A_27_617#_c_207_n N_A_27_617#_c_210_n
+ N_A_27_617#_c_220_n N_A_27_617#_c_212_n
+ PM_SKY130_OSU_SC_18T_HS__AOI21_L%A_27_617#
x_PM_SKY130_OSU_SC_18T_HS__AOI21_L%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_223_n
+ N_Y_c_226_n N_Y_c_227_n N_Y_c_229_n Y N_Y_c_232_n
+ PM_SKY130_OSU_SC_18T_HS__AOI21_L%Y
cc_1 N_GND_M1004_b N_A0_c_67_n 0.0660236f $X=-0.045 $Y=0 $X2=0.295 $Y2=2.63
cc_2 N_GND_M1004_b N_A0_c_68_n 0.0198745f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.69
cc_3 N_GND_c_3_p N_A0_c_68_n 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.69
cc_4 N_GND_c_4_p N_A0_c_68_n 0.00606474f $X=1.455 $Y=0.152 $X2=0.475 $Y2=1.69
cc_5 N_GND_c_5_p N_A0_c_68_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.69
cc_6 N_GND_M1004_b N_A0_c_72_n 0.0324933f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.77
cc_7 N_GND_c_3_p N_A0_c_72_n 0.00534003f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.77
cc_8 N_GND_M1004_b N_A0_c_74_n 0.0421132f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_9 N_GND_M1004_b N_A0_c_75_n 0.00438599f $X=-0.045 $Y=0 $X2=0.385 $Y2=2.765
cc_10 N_GND_M1004_b N_A1_M1002_g 0.0407759f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_11 N_GND_c_4_p N_A1_M1002_g 0.00606474f $X=1.455 $Y=0.152 $X2=0.835 $Y2=1.075
cc_12 N_GND_c_5_p N_A1_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=1.075
cc_13 N_GND_M1004_b N_A1_M1000_g 0.0273376f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_14 N_GND_M1004_b N_A1_c_108_n 0.0355308f $X=-0.045 $Y=0 $X2=0.815 $Y2=2.255
cc_15 N_GND_M1004_b N_A1_c_109_n 0.00889603f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.96
cc_16 N_GND_M1004_b N_A1_c_110_n 0.00478352f $X=-0.045 $Y=0 $X2=0.815 $Y2=2.255
cc_17 N_GND_M1004_b A1 0.00323672f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.96
cc_18 N_GND_M1004_b N_B0_M1005_g 0.0384502f $X=-0.045 $Y=0 $X2=1.325 $Y2=0.945
cc_19 N_GND_c_4_p N_B0_M1005_g 0.00606474f $X=1.455 $Y=0.152 $X2=1.325 $Y2=0.945
cc_20 N_GND_c_20_p N_B0_M1005_g 0.00713292f $X=1.54 $Y=0.825 $X2=1.325 $Y2=0.945
cc_21 N_GND_c_5_p N_B0_M1005_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.325 $Y2=0.945
cc_22 N_GND_M1004_b N_B0_M1001_g 5.06723e-19 $X=-0.045 $Y=0 $X2=1.335 $Y2=4.585
cc_23 N_GND_M1004_b N_B0_c_159_n 0.0493362f $X=-0.045 $Y=0 $X2=1.47 $Y2=2.745
cc_24 N_GND_M1004_b N_B0_c_160_n 0.0237317f $X=-0.045 $Y=0 $X2=1.47 $Y2=2.82
cc_25 N_GND_M1004_b N_B0_c_161_n 0.0498222f $X=-0.045 $Y=0 $X2=1.47 $Y2=1.86
cc_26 N_GND_c_20_p N_B0_c_161_n 0.00379395f $X=1.54 $Y=0.825 $X2=1.47 $Y2=1.86
cc_27 N_GND_M1004_b N_B0_c_163_n 0.0141127f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.59
cc_28 N_GND_M1004_b N_B0_c_164_n 0.00387834f $X=-0.045 $Y=0 $X2=1.25 $Y2=1.86
cc_29 N_GND_M1004_b N_B0_c_165_n 0.011995f $X=-0.045 $Y=0 $X2=1.53 $Y2=1.86
cc_30 N_GND_M1004_b B0 0.0176529f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.59
cc_31 N_GND_M1004_b N_Y_c_223_n 0.00156053f $X=-0.045 $Y=0 $X2=1.05 $Y2=0.825
cc_32 N_GND_c_4_p N_Y_c_223_n 0.00736239f $X=1.455 $Y=0.152 $X2=1.05 $Y2=0.825
cc_33 N_GND_c_5_p N_Y_c_223_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.05 $Y2=0.825
cc_34 N_GND_M1004_b N_Y_c_226_n 0.0225607f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.22
cc_35 N_GND_M1004_b N_Y_c_227_n 0.0138131f $X=-0.045 $Y=0 $X2=1.465 $Y2=1.48
cc_36 N_GND_c_20_p N_Y_c_227_n 0.00869812f $X=1.54 $Y=0.825 $X2=1.465 $Y2=1.48
cc_37 N_GND_M1004_b N_Y_c_229_n 0.00701376f $X=-0.045 $Y=0 $X2=1.195 $Y2=1.48
cc_38 N_GND_c_3_p N_Y_c_229_n 0.00100286f $X=0.26 $Y=0.825 $X2=1.195 $Y2=1.48
cc_39 N_GND_M1004_b Y 0.0092181f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.07
cc_40 N_GND_M1004_b N_Y_c_232_n 0.0114144f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.22
cc_41 N_VDD_M1003_b N_A0_M1003_g 0.0258897f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_42 N_VDD_c_42_p N_A0_M1003_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_43 N_VDD_c_43_p N_A0_M1003_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.475 $Y2=4.585
cc_44 N_VDD_c_44_p N_A0_M1003_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=4.585
cc_45 N_VDD_M1003_b N_A0_c_75_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.385
+ $Y2=2.765
cc_46 N_VDD_M1003_d A0 0.00612249f $X=0.55 $Y=3.085 $X2=0.385 $Y2=3.33
cc_47 N_VDD_M1003_b N_A1_M1000_g 0.0189802f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_48 N_VDD_c_43_p N_A1_M1000_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.905 $Y2=4.585
cc_49 N_VDD_c_49_p N_A1_M1000_g 0.00606474f $X=1.02 $Y=6.44 $X2=0.905 $Y2=4.585
cc_50 N_VDD_c_44_p N_A1_M1000_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.905 $Y2=4.585
cc_51 N_VDD_M1003_b N_A1_c_109_n 0.00476834f $X=-0.045 $Y=2.905 $X2=0.725
+ $Y2=2.96
cc_52 N_VDD_M1003_b A1 0.0103281f $X=-0.045 $Y=2.905 $X2=0.725 $Y2=2.96
cc_53 N_VDD_M1003_b N_B0_M1001_g 0.0246768f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=4.585
cc_54 N_VDD_c_49_p N_B0_M1001_g 0.00606474f $X=1.02 $Y=6.44 $X2=1.335 $Y2=4.585
cc_55 N_VDD_c_44_p N_B0_M1001_g 0.00468827f $X=1.02 $Y=6.47 $X2=1.335 $Y2=4.585
cc_56 N_VDD_M1003_b N_A_27_617#_c_207_n 0.00156053f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.135
cc_57 N_VDD_c_42_p N_A_27_617#_c_207_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=4.135
cc_58 N_VDD_c_44_p N_A_27_617#_c_207_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26
+ $Y2=4.135
cc_59 N_VDD_M1003_d N_A_27_617#_c_210_n 0.00743028f $X=0.55 $Y=3.085 $X2=1.035
+ $Y2=3.97
cc_60 N_VDD_c_43_p N_A_27_617#_c_210_n 0.0135055f $X=0.69 $Y=4.475 $X2=1.035
+ $Y2=3.97
cc_61 N_VDD_M1003_b N_A_27_617#_c_212_n 0.00155118f $X=-0.045 $Y=2.905 $X2=1.12
+ $Y2=4.135
cc_62 N_VDD_c_49_p N_A_27_617#_c_212_n 0.00734006f $X=1.02 $Y=6.44 $X2=1.12
+ $Y2=4.135
cc_63 N_VDD_c_44_p N_A_27_617#_c_212_n 0.00475776f $X=1.02 $Y=6.47 $X2=1.12
+ $Y2=4.135
cc_64 N_VDD_M1003_b N_Y_c_226_n 0.00917206f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.22
cc_65 N_VDD_c_49_p N_Y_c_226_n 0.00757793f $X=1.02 $Y=6.44 $X2=1.55 $Y2=2.22
cc_66 N_VDD_c_44_p N_Y_c_226_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.55 $Y2=2.22
cc_67 N_A0_c_67_n N_A1_M1002_g 0.00899556f $X=0.295 $Y=2.63 $X2=0.835 $Y2=1.075
cc_68 N_A0_c_68_n N_A1_M1002_g 0.0854438f $X=0.475 $Y=1.69 $X2=0.835 $Y2=1.075
cc_69 N_A0_c_67_n N_A1_M1000_g 0.00367405f $X=0.295 $Y=2.63 $X2=0.905 $Y2=4.585
cc_70 N_A0_c_74_n N_A1_M1000_g 0.0804191f $X=0.475 $Y=2.765 $X2=0.905 $Y2=4.585
cc_71 N_A0_c_75_n N_A1_M1000_g 0.00277246f $X=0.385 $Y=2.765 $X2=0.905 $Y2=4.585
cc_72 A0 N_A1_M1000_g 0.00309207f $X=0.385 $Y=3.33 $X2=0.905 $Y2=4.585
cc_73 N_A0_c_67_n N_A1_c_108_n 0.0125472f $X=0.295 $Y=2.63 $X2=0.815 $Y2=2.255
cc_74 N_A0_c_67_n N_A1_c_109_n 0.00365573f $X=0.295 $Y=2.63 $X2=0.725 $Y2=2.96
cc_75 N_A0_c_74_n N_A1_c_109_n 0.00281397f $X=0.475 $Y=2.765 $X2=0.725 $Y2=2.96
cc_76 N_A0_c_75_n N_A1_c_109_n 0.0297299f $X=0.385 $Y=2.765 $X2=0.725 $Y2=2.96
cc_77 N_A0_c_67_n N_A1_c_110_n 0.00661569f $X=0.295 $Y=2.63 $X2=0.815 $Y2=2.255
cc_78 N_A0_c_74_n A1 0.00417236f $X=0.475 $Y=2.765 $X2=0.725 $Y2=2.96
cc_79 N_A0_c_75_n A1 0.00775911f $X=0.385 $Y=2.765 $X2=0.725 $Y2=2.96
cc_80 A0 A1 0.00560453f $X=0.385 $Y=3.33 $X2=0.725 $Y2=2.96
cc_81 N_A0_c_75_n N_A_27_617#_M1003_s 0.00882571f $X=0.385 $Y=2.765 $X2=0.135
+ $Y2=3.085
cc_82 A0 N_A_27_617#_M1003_s 0.0124771f $X=0.385 $Y=3.33 $X2=0.135 $Y2=3.085
cc_83 N_A0_M1003_g N_A_27_617#_c_210_n 0.0152354f $X=0.475 $Y=4.585 $X2=1.035
+ $Y2=3.97
cc_84 N_A0_c_75_n N_A_27_617#_c_210_n 0.00155918f $X=0.385 $Y=2.765 $X2=1.035
+ $Y2=3.97
cc_85 A0 N_A_27_617#_c_210_n 0.00806826f $X=0.385 $Y=3.33 $X2=1.035 $Y2=3.97
cc_86 N_A0_c_75_n N_A_27_617#_c_220_n 0.00100283f $X=0.385 $Y=2.765 $X2=0.345
+ $Y2=3.97
cc_87 A0 N_A_27_617#_c_220_n 0.00366477f $X=0.385 $Y=3.33 $X2=0.345 $Y2=3.97
cc_88 N_A0_c_68_n N_Y_c_229_n 0.00104729f $X=0.475 $Y=1.69 $X2=1.195 $Y2=1.48
cc_89 N_A1_M1002_g N_B0_M1005_g 0.035383f $X=0.835 $Y=1.075 $X2=1.325 $Y2=0.945
cc_90 N_A1_c_108_n N_B0_c_159_n 0.0147459f $X=0.815 $Y=2.255 $X2=1.47 $Y2=2.745
cc_91 N_A1_M1000_g N_B0_c_160_n 0.0622722f $X=0.905 $Y=4.585 $X2=1.47 $Y2=2.82
cc_92 A1 N_B0_c_160_n 0.00105858f $X=0.725 $Y=2.96 $X2=1.47 $Y2=2.82
cc_93 N_A1_M1002_g N_B0_c_161_n 0.0039494f $X=0.835 $Y=1.075 $X2=1.47 $Y2=1.86
cc_94 N_A1_M1002_g N_B0_c_163_n 0.00326852f $X=0.835 $Y=1.075 $X2=1.165 $Y2=2.59
cc_95 N_A1_c_108_n N_B0_c_163_n 0.00506769f $X=0.815 $Y=2.255 $X2=1.165 $Y2=2.59
cc_96 N_A1_c_109_n N_B0_c_163_n 0.0109205f $X=0.725 $Y=2.96 $X2=1.165 $Y2=2.59
cc_97 N_A1_c_110_n N_B0_c_163_n 0.0226306f $X=0.815 $Y=2.255 $X2=1.165 $Y2=2.59
cc_98 N_A1_M1002_g N_B0_c_164_n 0.00477017f $X=0.835 $Y=1.075 $X2=1.25 $Y2=1.86
cc_99 N_A1_M1000_g B0 0.00717682f $X=0.905 $Y=4.585 $X2=1.165 $Y2=2.59
cc_100 N_A1_c_109_n B0 0.00705035f $X=0.725 $Y=2.96 $X2=1.165 $Y2=2.59
cc_101 A1 B0 0.00582284f $X=0.725 $Y=2.96 $X2=1.165 $Y2=2.59
cc_102 N_A1_M1000_g N_A_27_617#_c_210_n 0.0180368f $X=0.905 $Y=4.585 $X2=1.035
+ $Y2=3.97
cc_103 N_A1_M1002_g N_Y_c_223_n 0.00258639f $X=0.835 $Y=1.075 $X2=1.05 $Y2=0.825
cc_104 N_A1_c_108_n N_Y_c_223_n 3.56057e-19 $X=0.815 $Y=2.255 $X2=1.05 $Y2=0.825
cc_105 N_A1_M1000_g N_Y_c_226_n 8.50177e-19 $X=0.905 $Y=4.585 $X2=1.55 $Y2=2.22
cc_106 N_A1_c_109_n N_Y_c_226_n 0.00666053f $X=0.725 $Y=2.96 $X2=1.55 $Y2=2.22
cc_107 A1 N_Y_c_226_n 0.00511095f $X=0.725 $Y=2.96 $X2=1.55 $Y2=2.22
cc_108 N_A1_M1002_g N_Y_c_229_n 0.00584309f $X=0.835 $Y=1.075 $X2=1.195 $Y2=1.48
cc_109 N_A1_c_108_n N_Y_c_229_n 0.00171207f $X=0.815 $Y=2.255 $X2=1.195 $Y2=1.48
cc_110 N_A1_M1002_g Y 3.27704e-19 $X=0.835 $Y=1.075 $X2=1.55 $Y2=2.07
cc_111 N_B0_M1005_g N_Y_c_223_n 0.0147465f $X=1.325 $Y=0.945 $X2=1.05 $Y2=0.825
cc_112 N_B0_c_164_n N_Y_c_223_n 0.00317724f $X=1.25 $Y=1.86 $X2=1.05 $Y2=0.825
cc_113 N_B0_M1001_g N_Y_c_226_n 0.0166065f $X=1.335 $Y=4.585 $X2=1.55 $Y2=2.22
cc_114 N_B0_c_159_n N_Y_c_226_n 0.0192649f $X=1.47 $Y=2.745 $X2=1.55 $Y2=2.22
cc_115 N_B0_c_160_n N_Y_c_226_n 0.00834782f $X=1.47 $Y=2.82 $X2=1.55 $Y2=2.22
cc_116 N_B0_c_161_n N_Y_c_226_n 0.00170788f $X=1.47 $Y=1.86 $X2=1.55 $Y2=2.22
cc_117 N_B0_c_163_n N_Y_c_226_n 0.027719f $X=1.165 $Y=2.59 $X2=1.55 $Y2=2.22
cc_118 N_B0_c_165_n N_Y_c_226_n 0.0101032f $X=1.53 $Y=1.86 $X2=1.55 $Y2=2.22
cc_119 B0 N_Y_c_226_n 0.00715529f $X=1.165 $Y=2.59 $X2=1.55 $Y2=2.22
cc_120 N_B0_M1005_g N_Y_c_227_n 0.0119364f $X=1.325 $Y=0.945 $X2=1.465 $Y2=1.48
cc_121 N_B0_c_161_n N_Y_c_227_n 0.00145385f $X=1.47 $Y=1.86 $X2=1.465 $Y2=1.48
cc_122 N_B0_c_164_n N_Y_c_227_n 0.0028071f $X=1.25 $Y=1.86 $X2=1.465 $Y2=1.48
cc_123 N_B0_c_165_n N_Y_c_227_n 0.00728929f $X=1.53 $Y=1.86 $X2=1.465 $Y2=1.48
cc_124 N_B0_M1005_g N_Y_c_229_n 6.90188e-19 $X=1.325 $Y=0.945 $X2=1.195 $Y2=1.48
cc_125 N_B0_c_164_n N_Y_c_229_n 0.00487807f $X=1.25 $Y=1.86 $X2=1.195 $Y2=1.48
cc_126 N_B0_M1005_g Y 0.00272607f $X=1.325 $Y=0.945 $X2=1.55 $Y2=2.07
cc_127 N_B0_c_159_n Y 0.00138242f $X=1.47 $Y=2.745 $X2=1.55 $Y2=2.07
cc_128 N_B0_c_161_n Y 0.01116f $X=1.47 $Y=1.86 $X2=1.55 $Y2=2.07
cc_129 N_B0_c_163_n Y 0.00642461f $X=1.165 $Y=2.59 $X2=1.55 $Y2=2.07
cc_130 N_B0_c_165_n Y 0.0205824f $X=1.53 $Y=1.86 $X2=1.55 $Y2=2.07
cc_131 N_B0_c_159_n N_Y_c_232_n 0.00517151f $X=1.47 $Y=2.745 $X2=1.55 $Y2=2.22
cc_132 N_B0_c_161_n N_Y_c_232_n 8.18646e-19 $X=1.47 $Y=1.86 $X2=1.55 $Y2=2.22
cc_133 N_B0_c_163_n N_Y_c_232_n 0.00655582f $X=1.165 $Y=2.59 $X2=1.55 $Y2=2.22
cc_134 N_B0_c_165_n N_Y_c_232_n 0.00439213f $X=1.53 $Y=1.86 $X2=1.55 $Y2=2.22
