* File: sky130_osu_sc_12T_hs__or2_l.spice
* Created: Fri Nov 12 15:13:08 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__or2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_l  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_A_27_605#_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_GND_M1000_d N_A_M1000_g N_A_27_605#_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_27_605#_M1001_g N_GND_M1000_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_110_605# N_B_M1002_g N_A_27_605#_M1002_s N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=19.9167 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_VDD_M1004_d N_A_M1004_g A_110_605# N_VDD_M1002_b PSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=19.9167 M=1 R=5.6 SA=75000.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_27_605#_M1005_g N_VDD_M1004_d N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=3.23635 P=7.21
pX7_noxref noxref_8 B B PROBETYPE=1
pX8_noxref noxref_9 A A PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_l.pxi.spice"
*
.ends
*
*
