* File: sky130_osu_sc_15T_ls__dffr_l.spice
* Created: Fri Nov 12 14:55:59 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__dffr_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__dffr_l  GND VDD RN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* RN	RN
* VDD	VDD
* GND	GND
MM1013 N_A_110_115#_M1013_d N_RN_M1013_g N_GND_M1013_s N_GND_M1013_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_217_713#_M1009_d N_A_110_115#_M1009_g N_GND_M1009_s N_GND_M1013_b
+ NSHORT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_A_342_466#_M1001_g N_A_217_713#_M1009_d N_GND_M1013_b
+ NSHORT L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1002 A_576_115# N_D_M1002_g N_GND_M1002_s N_GND_M1013_b NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1028 N_A_342_466#_M1028_d N_A_618_89#_M1028_g A_576_115# N_GND_M1013_b NSHORT
+ L=0.15 W=0.74 AD=0.1665 AS=0.0777 PD=1.19 PS=0.95 NRD=13.776 NRS=8.1 M=1
+ R=4.93333 SA=75000.6 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1024 A_768_115# N_CK_M1024_g N_A_342_466#_M1028_d N_GND_M1013_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1665 PD=0.95 PS=1.19 NRD=8.1 NRS=13.776 M=1 R=4.93333
+ SA=75001.1 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1026 N_GND_M1026_d N_A_217_713#_M1026_g A_768_115# N_GND_M1013_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.0777 PD=1.02 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.5 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1020 A_926_115# N_A_217_713#_M1020_g N_GND_M1026_d N_GND_M1013_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1036 PD=0.95 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1010 N_A_998_115#_M1010_d N_CK_M1010_g A_926_115# N_GND_M1013_b NSHORT L=0.15
+ W=0.74 AD=0.1665 AS=0.0777 PD=1.19 PS=0.95 NRD=13.776 NRS=8.1 M=1 R=4.93333
+ SA=75002.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1011 A_1118_115# N_A_618_89#_M1011_g N_A_998_115#_M1010_d N_GND_M1013_b NSHORT
+ L=0.15 W=0.74 AD=0.0777 AS=0.1665 PD=0.95 PS=1.19 NRD=8.1 NRS=13.776 M=1
+ R=4.93333 SA=75002.9 SB=75001 A=0.111 P=1.78 MULT=1
MM1016 N_GND_M1016_d N_A_1160_89#_M1016_g A_1118_115# N_GND_M1013_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.0777 PD=1.02 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75003.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_618_89#_M1004_d N_CK_M1004_g N_GND_M1016_d N_GND_M1013_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_1160_89#_M1005_d N_A_998_115#_M1005_g N_GND_M1005_s N_GND_M1013_b
+ NSHORT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1006 N_GND_M1006_d N_A_110_115#_M1006_g N_A_1160_89#_M1005_d N_GND_M1013_b
+ NSHORT L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_A_1160_89#_M1007_g N_QN_M1007_s N_GND_M1013_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1003 N_Q_M1003_d N_QN_M1003_g N_GND_M1007_d N_GND_M1013_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_A_110_115#_M1000_d N_RN_M1000_g N_VDD_M1000_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1018 A_300_713# N_A_110_115#_M1018_g N_A_217_713#_M1018_s N_VDD_M1000_b
+ PHIGHVT L=0.15 W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1
+ R=8.4 SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1022 N_VDD_M1022_d N_A_342_466#_M1022_g A_300_713# N_VDD_M1000_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 A_576_565# N_D_M1008_g N_VDD_M1008_s N_VDD_M1000_b PHIGHVT L=0.15 W=2
+ AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75003.7 A=0.3 P=4.3 MULT=1
MM1015 N_A_342_466#_M1015_d N_CK_M1015_g A_576_565# N_VDD_M1000_b PHIGHVT L=0.15
+ W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75000.5 SB=75003.3 A=0.3 P=4.3 MULT=1
MM1021 A_768_565# N_A_618_89#_M1021_g N_A_342_466#_M1015_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75001.1 SB=75002.7 A=0.3 P=4.3 MULT=1
MM1019 N_VDD_M1019_d N_A_217_713#_M1019_g A_768_565# N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333
+ SA=75001.5 SB=75002.4 A=0.3 P=4.3 MULT=1
MM1027 A_926_565# N_A_217_713#_M1027_g N_VDD_M1019_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333
+ SA=75001.9 SB=75001.9 A=0.3 P=4.3 MULT=1
MM1029 N_A_998_115#_M1029_d N_A_618_89#_M1029_g A_926_565# N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75002.3 SB=75001.6 A=0.3 P=4.3 MULT=1
MM1030 A_1118_565# N_CK_M1030_g N_A_998_115#_M1029_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75002.9 SB=75001 A=0.3 P=4.3 MULT=1
MM1031 N_VDD_M1031_d N_A_1160_89#_M1031_g A_1118_565# N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333
+ SA=75003.3 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1023 N_A_618_89#_M1023_d N_CK_M1023_g N_VDD_M1031_d N_VDD_M1000_b PHIGHVT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.7 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1012 A_1466_713# N_A_998_115#_M1012_g N_A_1160_89#_M1012_s N_VDD_M1000_b
+ PHIGHVT L=0.15 W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1
+ R=8.4 SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_VDD_M1017_d N_A_110_115#_M1017_g A_1466_713# N_VDD_M1000_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1014 N_VDD_M1014_d N_A_1160_89#_M1014_g N_QN_M1014_s N_VDD_M1000_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_Q_M1025_d N_QN_M1025_g N_VDD_M1014_d N_VDD_M1000_b PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref N_GND_M1013_b N_VDD_M1000_b NWDIODE A=28.4232 P=25.17
pX33_noxref noxref_24 RN RN PROBETYPE=1
pX34_noxref noxref_25 D D PROBETYPE=1
pX35_noxref noxref_26 CK CK PROBETYPE=1
pX36_noxref noxref_27 QN QN PROBETYPE=1
pX37_noxref noxref_28 Q Q PROBETYPE=1
c_1607 A_926_565# 0 1.57671e-19 $X=4.63 $Y=2.825
*
.include "sky130_osu_sc_15T_ls__dffr_l.pxi.spice"
*
.ends
*
*
