* File: sky130_osu_sc_15T_hs__addh_1.pex.spice
* Created: Fri Nov 12 14:26:25 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%GND 1 2 45 47 55 57 70 86 88
c95 45 0 1.81192e-19 $X=-0.045 $Y=0
r96 86 88 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r97 72 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r98 68 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r99 68 70 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.74
r100 58 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r101 57 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r102 53 81 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r103 53 55 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.885
r104 47 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r105 45 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r106 45 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r107 45 72 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r108 45 57 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r109 45 58 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r110 45 47 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r111 2 70 91 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.74
r112 1 55 182 $w=1.7e-07 $l=3.97618e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.885
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%VDD 1 2 3 37 39 46 50 56 60 68 74 82 86
r56 82 86 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=3.74 $Y2=5.397
r57 74 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=5.36
+ $X2=3.74 $Y2=5.36
r58 72 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=5.397
+ $X2=3.05 $Y2=5.397
r59 72 74 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=5.397
+ $X2=3.74 $Y2=5.397
r60 68 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.05 $Y=3.215
+ $X2=3.05 $Y2=4.575
r61 66 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=5.245
+ $X2=3.05 $Y2=5.397
r62 66 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=5.245
+ $X2=3.05 $Y2=4.575
r63 63 65 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=5.397
+ $X2=2.38 $Y2=5.397
r64 61 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=5.397
+ $X2=1.61 $Y2=5.397
r65 61 63 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=5.397
+ $X2=1.7 $Y2=5.397
r66 60 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=5.397
+ $X2=3.05 $Y2=5.397
r67 60 65 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=5.397
+ $X2=2.38 $Y2=5.397
r68 56 59 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.61 $Y=3.555
+ $X2=1.61 $Y2=4.575
r69 54 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=5.245
+ $X2=1.61 $Y2=5.397
r70 54 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.61 $Y=5.245
+ $X2=1.61 $Y2=4.575
r71 51 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=5.397
+ $X2=0.75 $Y2=5.397
r72 51 53 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=5.397
+ $X2=1.02 $Y2=5.397
r73 50 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=5.397
+ $X2=1.61 $Y2=5.397
r74 50 53 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=5.397
+ $X2=1.02 $Y2=5.397
r75 46 49 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.75 $Y=3.215
+ $X2=0.75 $Y2=4.575
r76 44 77 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=5.245
+ $X2=0.75 $Y2=5.397
r77 44 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.75 $Y=5.245
+ $X2=0.75 $Y2=4.575
r78 41 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r79 39 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=5.397
+ $X2=0.75 $Y2=5.397
r80 39 41 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=5.397
+ $X2=0.34 $Y2=5.397
r81 37 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=5.245 $X2=3.74 $Y2=5.33
r82 37 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r83 37 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r84 37 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r85 37 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r86 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r87 3 71 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=2.825 $X2=3.05 $Y2=4.575
r88 3 68 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=2.825 $X2=3.05 $Y2=3.215
r89 2 59 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.825 $X2=1.61 $Y2=4.575
r90 2 56 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=2.825 $X2=1.61 $Y2=3.555
r91 1 49 240 $w=1.7e-07 $l=1.8473e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.75 $Y2=4.575
r92 1 46 240 $w=1.7e-07 $l=4.79687e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.75 $Y2=3.215
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%CON 1 3 4 15 19 22 29 31 32 35 39 41 43
+ 45 49 55 58 59 64 67
c129 67 0 2.55765e-19 $X=3.42 $Y=1.59
c130 59 0 1.57622e-19 $X=0.78 $Y=1.59
c131 43 0 1.92558e-19 $X=3.42 $Y=1.505
c132 31 0 1.81192e-19 $X=2.62 $Y=1.675
r133 59 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.59
+ $X2=0.635 $Y2=1.59
r134 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.59
+ $X2=2.62 $Y2=1.59
r135 58 59 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.59
+ $X2=0.78 $Y2=1.59
r136 57 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.59
+ $X2=3.42 $Y2=1.59
r137 54 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.59
+ $X2=2.62 $Y2=1.59
r138 49 51 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.84 $Y=3.215
+ $X2=3.84 $Y2=4.575
r139 47 49 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.84 $Y=2.775
+ $X2=3.84 $Y2=3.215
r140 43 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.505
+ $X2=3.42 $Y2=1.59
r141 43 45 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.42 $Y=1.505
+ $X2=3.42 $Y2=1.065
r142 42 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.69
+ $X2=2.62 $Y2=2.69
r143 41 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.69
+ $X2=3.84 $Y2=2.775
r144 41 42 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.69
+ $X2=2.705 $Y2=2.69
r145 40 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.59
+ $X2=2.62 $Y2=1.59
r146 39 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.59
+ $X2=3.42 $Y2=1.59
r147 39 40 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.59
+ $X2=2.705 $Y2=1.59
r148 35 37 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.62 $Y=3.215
+ $X2=2.62 $Y2=4.575
r149 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.775
+ $X2=2.62 $Y2=2.69
r150 33 35 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.62 $Y=2.775
+ $X2=2.62 $Y2=3.215
r151 32 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.605
+ $X2=2.62 $Y2=2.69
r152 31 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.675
+ $X2=2.62 $Y2=1.59
r153 31 32 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.675
+ $X2=2.62 $Y2=2.605
r154 29 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.59
+ $X2=0.635 $Y2=1.59
r155 26 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.35 $Y=1.59
+ $X2=0.635 $Y2=1.59
r156 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.59 $X2=0.35 $Y2=1.59
r157 22 24 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.59
+ $X2=0.382 $Y2=1.755
r158 22 23 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.59
+ $X2=0.382 $Y2=1.425
r159 19 24 1061.43 $w=1.5e-07 $l=2.07e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=1.755
r160 15 23 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=1.425
r161 4 51 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=2.825 $X2=3.84 $Y2=4.575
r162 4 49 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=2.825 $X2=3.84 $Y2=3.215
r163 3 37 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=2.825 $X2=2.62 $Y2=4.575
r164 3 35 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=2.825 $X2=2.62 $Y2=3.215
r165 1 45 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=1.065
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%B 3 7 11 15 18 22 25 30 39 42 44
c102 44 0 4.99902e-20 $X=3.21 $Y=1.96
c103 22 0 1.42567e-19 $X=3.205 $Y=1.96
c104 18 0 1.57622e-19 $X=0.905 $Y=1.96
c105 7 0 4.43035e-20 $X=0.965 $Y=3.825
r106 41 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=3.205 $Y=1.96
+ $X2=3.21 $Y2=1.96
r107 41 42 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.205 $Y=1.96
+ $X2=3.06 $Y2=1.96
r108 39 42 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=1.962
+ $X2=3.06 $Y2=1.962
r109 37 39 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=1.96
+ $X2=1.05 $Y2=1.96
r110 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=1.96
+ $X2=3.205 $Y2=1.96
r111 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=1.96
r112 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.96 $X2=3.205 $Y2=1.96
r113 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.96
+ $X2=3.205 $Y2=2.125
r114 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.96 $X2=0.905 $Y2=1.96
r115 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=2.125
r116 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.96
+ $X2=0.905 $Y2=1.795
r117 15 23 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=3.265 $Y=3.825
+ $X2=3.265 $Y2=2.125
r118 9 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.795
+ $X2=3.205 $Y2=1.96
r119 9 11 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.205 $Y=1.795
+ $X2=3.205 $Y2=0.995
r120 7 20 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=0.965 $Y=3.825
+ $X2=0.965 $Y2=2.125
r121 3 19 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.965 $Y=0.895
+ $X2=0.965 $Y2=1.795
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%A 3 7 11 15 18 22 26 31 40 42 43
c87 22 0 1.74252e-19 $X=3.685 $Y=2.33
r88 42 43 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.33
+ $X2=3.54 $Y2=2.33
r89 40 43 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.327
+ $X2=3.54 $Y2=2.327
r90 38 40 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.33
+ $X2=1.53 $Y2=2.33
r91 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.33
+ $X2=3.685 $Y2=2.33
r92 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.33
+ $X2=1.385 $Y2=2.33
r93 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.33 $X2=3.685 $Y2=2.33
r94 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.33
+ $X2=3.685 $Y2=2.495
r95 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.33
+ $X2=3.685 $Y2=2.165
r96 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.33 $X2=1.385 $Y2=2.33
r97 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.33
+ $X2=1.385 $Y2=2.495
r98 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.33
+ $X2=1.385 $Y2=2.165
r99 15 23 599.936 $w=1.5e-07 $l=1.17e-06 $layer=POLY_cond $X=3.635 $Y=0.995
+ $X2=3.635 $Y2=2.165
r100 11 24 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.625 $Y=3.825
+ $X2=3.625 $Y2=2.495
r101 7 20 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.395 $Y=3.825
+ $X2=1.395 $Y2=2.495
r102 3 19 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.325 $Y=0.895
+ $X2=1.325 $Y2=2.165
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%A_208_565# 1 3 9 10 13 15 17 19 21 22 24
+ 26 29 31 35 38 42 43 46 49 51
c116 29 0 2.52869e-20 $X=2.835 $Y=3.825
c117 24 0 8.1513e-20 $X=2.775 $Y=1.49
r118 51 53 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.695
+ $X2=1.825 $Y2=1.695
r119 50 51 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.695
+ $X2=1.725 $Y2=1.695
r120 48 51 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.86
+ $X2=1.725 $Y2=1.695
r121 48 49 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=1.86
+ $X2=1.725 $Y2=2.665
r122 44 50 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.53
+ $X2=1.54 $Y2=1.695
r123 44 46 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.54 $Y=1.53
+ $X2=1.54 $Y2=0.885
r124 42 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=2.75
+ $X2=1.725 $Y2=2.665
r125 42 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=2.75
+ $X2=1.265 $Y2=2.75
r126 38 40 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.18 $Y=3.555
+ $X2=1.18 $Y2=4.575
r127 36 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=2.835
+ $X2=1.265 $Y2=2.75
r128 36 38 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.18 $Y=2.835
+ $X2=1.18 $Y2=3.555
r129 34 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.695 $X2=1.825 $Y2=1.695
r130 32 34 23.6453 $w=2.65e-07 $l=1.3e-07 $layer=POLY_cond $X=1.825 $Y=1.565
+ $X2=1.825 $Y2=1.695
r131 27 29 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=2.835 $Y=2.485
+ $X2=2.835 $Y2=3.825
r132 24 26 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.775 $Y=1.49
+ $X2=2.775 $Y2=0.995
r133 23 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.565
+ $X2=2.285 $Y2=1.565
r134 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.565
+ $X2=2.775 $Y2=1.49
r135 22 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.565
+ $X2=2.36 $Y2=1.565
r136 19 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.49
+ $X2=2.285 $Y2=1.565
r137 19 21 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.285 $Y=1.49
+ $X2=2.285 $Y2=0.995
r138 18 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.41
+ $X2=1.885 $Y2=2.41
r139 17 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.41
+ $X2=2.835 $Y2=2.485
r140 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.41 $X2=1.96
+ $Y2=2.41
r141 16 32 16.0701 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.565
+ $X2=1.825 $Y2=1.565
r142 15 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.565
+ $X2=2.285 $Y2=1.565
r143 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.565
+ $X2=1.96 $Y2=1.565
r144 11 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.485
+ $X2=1.885 $Y2=2.41
r145 11 13 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=1.885 $Y=2.485
+ $X2=1.885 $Y2=3.825
r146 10 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.335
+ $X2=1.885 $Y2=2.41
r147 9 34 39.0139 $w=2.65e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.885 $Y=1.86
+ $X2=1.825 $Y2=1.695
r148 9 10 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=1.86
+ $X2=1.885 $Y2=2.335
r149 3 40 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.825 $X2=1.18 $Y2=4.575
r150 3 38 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.825 $X2=1.18 $Y2=3.555
r151 1 46 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.885
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%S 1 3 10 16 26 29 32
c31 32 0 4.43035e-20 $X=0.26 $Y=3.07
r32 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.07
r33 24 26 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=2.125
r34 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.33
+ $X2=0.26 $Y2=1.215
r35 23 26 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.33
+ $X2=0.26 $Y2=2.125
r36 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=4.575
r37 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.07
+ $X2=0.26 $Y2=3.07
r38 16 19 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.26 $Y=3.07
+ $X2=0.26 $Y2=3.215
r39 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.215
+ $X2=0.26 $Y2=1.215
r40 10 13 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.26 $Y=0.885
+ $X2=0.26 $Y2=1.215
r41 3 21 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r42 3 19 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.215
r43 1 10 182 $w=1.7e-07 $l=3.67219e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.885
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%CO 1 3 11 15 23 26 27 30
c51 26 0 2.52869e-20 $X=2.175 $Y=2.7
r52 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.7
+ $X2=2.175 $Y2=2.7
r53 26 28 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.7
+ $X2=2.137 $Y2=2.785
r54 26 27 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.7
+ $X2=2.137 $Y2=2.615
r55 21 23 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.25
+ $X2=2.175 $Y2=1.25
r56 19 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=1.335
+ $X2=2.175 $Y2=1.25
r57 19 27 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=2.175 $Y=1.335
+ $X2=2.175 $Y2=2.615
r58 15 17 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.1 $Y=3.215
+ $X2=2.1 $Y2=4.575
r59 15 28 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.1 $Y=3.215 $X2=2.1
+ $Y2=2.785
r60 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.165
+ $X2=2.07 $Y2=1.25
r61 9 11 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.07 $Y=1.165
+ $X2=2.07 $Y2=0.74
r62 3 17 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=2.825 $X2=2.1 $Y2=4.575
r63 3 15 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=2.825 $X2=2.1 $Y2=3.215
r64 1 11 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_HS__ADDH_1%A_570_115# 1 2 11 13 14
r11 15 17 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.85 $Y=0.645
+ $X2=3.85 $Y2=0.74
r12 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.56
+ $X2=3.85 $Y2=0.645
r13 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.56
+ $X2=3.075 $Y2=0.56
r14 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.645
+ $X2=3.075 $Y2=0.56
r15 9 11 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.99 $Y=0.645
+ $X2=2.99 $Y2=0.74
r16 2 17 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.74
r17 1 11 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.74
.ends

