magic
tech sky130A
magscale 1 2
timestamp 1606864602
<< checkpaint >>
rect -1209 -1243 1345 2575
<< nwell >>
rect -9 581 199 1341
<< nmos >>
rect 80 115 110 451
<< pmos >>
rect 80 817 110 1217
<< ndiff >>
rect 27 403 80 451
rect 27 131 35 403
rect 69 131 80 403
rect 27 115 80 131
rect 110 403 163 451
rect 110 131 121 403
rect 155 131 163 403
rect 110 115 163 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 861 35 1201
rect 69 861 80 1201
rect 27 817 80 861
rect 110 1201 163 1217
rect 110 861 121 1201
rect 155 861 163 1201
rect 110 817 163 861
<< ndiffc >>
rect 35 131 69 403
rect 121 131 155 403
<< pdiffc >>
rect 35 861 69 1201
rect 121 861 155 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1271 85 1305
<< poly >>
rect 80 1217 110 1243
rect 80 451 110 817
rect 80 80 110 115
<< locali >>
rect 0 1311 198 1332
rect 0 1271 51 1311
rect 85 1271 198 1311
rect 35 1201 69 1271
rect 35 845 69 861
rect 121 1201 155 1271
rect 121 845 155 861
rect 35 403 69 419
rect 35 61 69 131
rect 121 403 155 419
rect 121 61 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1311 198 1332
rect 0 1277 51 1311
rect 85 1277 198 1311
rect 0 1271 198 1277
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
