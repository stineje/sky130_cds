* File: sky130_osu_sc_15T_ls__and2_6.pex.spice
* Created: Fri Nov 12 14:53:48 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__AND2_6%GND 1 2 3 4 47 49 57 59 66 68 75 77 85
+ 95 97
r105 95 97 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.06 $Y2=0.152
r106 83 85 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.7 $Y=0.305
+ $X2=3.7 $Y2=0.74
r107 78 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.152
+ $X2=2.84 $Y2=0.152
r108 77 83 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=3.615 $Y=0.152
+ $X2=3.7 $Y2=0.305
r109 73 91 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.152
r110 73 75 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.74
r111 69 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r112 68 91 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.152
r113 64 90 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r114 64 66 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.74
r115 59 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r116 55 57 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r117 47 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=0.19
+ $X2=3.06 $Y2=0.19
r118 47 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r119 47 55 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r120 47 49 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r121 47 60 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r122 47 77 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.615 $Y2=0.152
r123 47 78 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.925 $Y2=0.152
r124 47 68 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r125 47 69 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r126 47 59 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r127 47 60 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r128 47 49 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r129 4 85 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.74
r130 3 75 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.74
r131 2 66 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.74
r132 1 57 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_6%VDD 1 2 3 4 5 41 45 49 55 59 65 69 75 79
+ 86 97 101
r70 97 101 1.26676 $w=3.05e-07 $l=2.72e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=3.06 $Y2=5.397
r71 91 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r72 86 89 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.7 $Y=3.215
+ $X2=3.7 $Y2=4.575
r73 84 89 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.7 $Y=5.245 $X2=3.7
+ $Y2=4.575
r74 82 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.06 $Y=5.36
+ $X2=3.06 $Y2=5.36
r75 80 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=2.84 $Y2=5.397
r76 80 82 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.925 $Y=5.397
+ $X2=3.06 $Y2=5.397
r77 79 84 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.7 $Y2=5.245
r78 79 82 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=3.615 $Y=5.397
+ $X2=3.06 $Y2=5.397
r79 75 78 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.215
+ $X2=2.84 $Y2=4.575
r80 73 95 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=5.397
r81 73 78 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.575
r82 70 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r83 70 72 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r84 69 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.397
r85 69 72 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r86 65 68 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.215
+ $X2=1.98 $Y2=4.575
r87 63 94 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r88 63 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.575
r89 60 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r90 60 62 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r91 59 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r92 59 62 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r93 55 58 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=3.555
+ $X2=1.12 $Y2=4.575
r94 53 93 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r95 53 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.575
r96 50 91 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r97 50 52 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r98 49 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r99 49 52 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r100 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.895
+ $X2=0.26 $Y2=4.575
r101 43 91 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r102 43 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.575
r103 41 82 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=5.245 $X2=3.06 $Y2=5.33
r104 41 72 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r105 41 62 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r106 41 52 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r107 41 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r108 5 89 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=4.575
r109 5 86 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=2.825 $X2=3.7 $Y2=3.215
r110 4 78 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.575
r111 4 75 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.215
r112 3 68 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.575
r113 3 65 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.215
r114 2 58 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r115 2 55 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.555
r116 1 48 400 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r117 1 45 400 $w=1.7e-07 $l=1.13077e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_6%A 3 7 12 15 23
r29 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=3.07
+ $X2=0.24 $Y2=3.07
r30 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=3.07
+ $X2=0.235 $Y2=3.07
r31 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.235 $Y=2.505
+ $X2=0.235 $Y2=3.07
r32 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.235
+ $Y=2.505 $X2=0.235 $Y2=2.505
r33 10 12 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.235 $Y=2.505
+ $X2=0.475 $Y2=2.505
r34 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=2.505
r35 5 7 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=3.825
r36 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=2.505
r37 1 3 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_6%B 3 7 10 13 21
c38 7 0 1.42883e-19 $X=0.905 $Y=3.825
r39 19 21 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.915 $Y=2.7
+ $X2=0.92 $Y2=2.7
r40 16 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.915 $Y=2.7
+ $X2=0.915 $Y2=2.7
r41 13 16 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.915 $Y=2.165
+ $X2=0.915 $Y2=2.7
r42 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=2.165 $X2=0.915 $Y2=2.165
r43 10 11 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.165
+ $X2=0.905 $Y2=2
r44 5 10 49.0931 $w=2.9e-07 $l=1.7e-07 $layer=POLY_cond $X=0.905 $Y=2.335
+ $X2=0.905 $Y2=2.165
r45 5 7 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=0.905 $Y=2.335
+ $X2=0.905 $Y2=3.825
r46 3 11 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=2
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_6%A_27_115# 1 3 11 14 15 17 18 20 24 26 28
+ 29 31 35 37 39 40 42 46 48 50 51 53 57 60 61 63 64 66 70 72 74 75 80 81 82 83
+ 84 85 86 87 88 91 94 97 101 103 110
c188 57 0 1.33323e-19 $X=3.055 $Y=0.945
c189 46 0 1.33323e-19 $X=2.625 $Y=0.945
c190 35 0 1.33323e-19 $X=2.195 $Y=0.945
c191 24 0 1.33323e-19 $X=1.765 $Y=0.945
r192 108 110 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.575 $Y=3.39
+ $X2=0.69 $Y2=3.39
r193 105 107 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=1.675
+ $X2=0.575 $Y2=1.675
r194 101 107 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=1.675
+ $X2=0.575 $Y2=1.675
r195 101 103 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.66 $Y=1.675
+ $X2=1.395 $Y2=1.675
r196 97 99 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=3.555
+ $X2=0.69 $Y2=4.575
r197 95 110 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.475
+ $X2=0.69 $Y2=3.39
r198 95 97 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.475
+ $X2=0.69 $Y2=3.555
r199 94 108 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.575 $Y=3.305
+ $X2=0.575 $Y2=3.39
r200 93 107 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.575 $Y=1.76
+ $X2=0.575 $Y2=1.675
r201 93 94 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=0.575 $Y=1.76
+ $X2=0.575 $Y2=3.305
r202 89 105 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=1.675
r203 89 91 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.74
r204 78 103 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.675 $X2=1.395 $Y2=1.675
r205 78 79 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.675
+ $X2=1.395 $Y2=1.84
r206 75 78 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.395 $Y=1.585
+ $X2=1.395 $Y2=1.675
r207 75 76 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=1.585
+ $X2=1.395 $Y2=1.51
r208 72 74 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.485 $Y=2.7
+ $X2=3.485 $Y2=3.825
r209 68 70 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.485 $Y=1.51
+ $X2=3.485 $Y2=0.945
r210 67 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.625
+ $X2=3.055 $Y2=2.625
r211 66 72 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.485 $Y2=2.7
r212 66 67 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.625
+ $X2=3.13 $Y2=2.625
r213 65 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.585
+ $X2=3.055 $Y2=1.585
r214 64 68 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.585
+ $X2=3.485 $Y2=1.51
r215 64 65 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.585
+ $X2=3.13 $Y2=1.585
r216 61 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.7 $X2=3.055
+ $Y2=2.625
r217 61 63 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.055 $Y=2.7
+ $X2=3.055 $Y2=3.825
r218 60 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=2.55
+ $X2=3.055 $Y2=2.625
r219 59 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.66
+ $X2=3.055 $Y2=1.585
r220 59 60 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.055 $Y=1.66
+ $X2=3.055 $Y2=2.55
r221 55 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.51
+ $X2=3.055 $Y2=1.585
r222 55 57 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.055 $Y=1.51
+ $X2=3.055 $Y2=0.945
r223 54 86 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.625
+ $X2=2.625 $Y2=2.625
r224 53 88 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=3.055 $Y2=2.625
r225 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.625
+ $X2=2.7 $Y2=2.625
r226 52 85 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.585
+ $X2=2.625 $Y2=1.585
r227 51 87 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.585
+ $X2=3.055 $Y2=1.585
r228 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.585
+ $X2=2.7 $Y2=1.585
r229 48 86 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=2.625
r230 48 50 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r231 44 85 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.625 $Y2=1.585
r232 44 46 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.625 $Y2=0.945
r233 43 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r234 42 86 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.625
r235 42 43 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r236 41 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.585
+ $X2=2.195 $Y2=1.585
r237 40 85 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.625 $Y2=1.585
r238 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.27 $Y2=1.585
r239 37 84 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=2.625
r240 37 39 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r241 33 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=1.585
r242 33 35 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=0.945
r243 32 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r244 31 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r245 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r246 30 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.585
+ $X2=1.765 $Y2=1.585
r247 29 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=2.195 $Y2=1.585
r248 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=1.84 $Y2=1.585
r249 26 82 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r250 26 28 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r251 22 81 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=1.585
r252 22 24 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=0.945
r253 21 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.53 $Y=1.585
+ $X2=1.395 $Y2=1.585
r254 20 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.585
+ $X2=1.765 $Y2=1.585
r255 20 21 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.69 $Y=1.585
+ $X2=1.53 $Y2=1.585
r256 19 80 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.625
+ $X2=1.335 $Y2=2.625
r257 18 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r258 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.41 $Y2=2.625
r259 15 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=2.625
r260 15 17 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r261 14 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.55
+ $X2=1.335 $Y2=2.625
r262 14 79 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.335 $Y=2.55
+ $X2=1.335 $Y2=1.84
r263 11 76 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.335 $Y=0.945
+ $X2=1.335 $Y2=1.51
r264 3 99 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.575
r265 3 97 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.555
r266 1 91 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_6%Y 1 2 3 7 8 9 26 32 40 46 54 60 67 68 70
+ 72 74 77 78 79 80 81 82 83
c124 82 0 1.33323e-19 $X=3.27 $Y=1.335
c125 79 0 2.66647e-19 $X=2.555 $Y=1.22
c126 67 0 1.33323e-19 $X=1.55 $Y=1.335
c127 32 0 1.42883e-19 $X=1.55 $Y=2.33
r128 83 95 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=2.215
+ $X2=3.27 $Y2=2.33
r129 82 93 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=1.22
r130 82 83 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=3.27 $Y=1.335
+ $X2=3.27 $Y2=2.215
r131 81 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=2.33
+ $X2=2.41 $Y2=2.33
r132 80 95 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=2.33
+ $X2=3.27 $Y2=2.33
r133 80 81 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=2.33
+ $X2=2.555 $Y2=2.33
r134 79 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.555 $Y=1.22
+ $X2=2.41 $Y2=1.22
r135 78 93 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=3.27 $Y2=1.22
r136 78 79 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.125 $Y=1.22
+ $X2=2.555 $Y2=1.22
r137 77 91 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.215
+ $X2=2.41 $Y2=2.33
r138 76 89 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r139 76 77 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.215
r140 75 87 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.33
+ $X2=1.55 $Y2=2.33
r141 74 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=2.41 $Y2=2.33
r142 74 75 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=1.695 $Y2=2.33
r143 73 85 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r144 72 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r145 72 73 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r146 68 87 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r147 68 70 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r148 67 85 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r149 67 70 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r150 63 65 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.27 $Y=3.215
+ $X2=3.27 $Y2=4.575
r151 60 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=2.33
+ $X2=3.27 $Y2=2.33
r152 60 63 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.27 $Y=2.33
+ $X2=3.27 $Y2=3.215
r153 57 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.27 $Y=1.22
+ $X2=3.27 $Y2=1.22
r154 54 57 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.27 $Y=0.74
+ $X2=3.27 $Y2=1.22
r155 49 51 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.215
+ $X2=2.41 $Y2=4.575
r156 46 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=2.33
r157 46 49 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=3.215
r158 43 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r159 40 43 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.41 $Y=0.74
+ $X2=2.41 $Y2=1.22
r160 35 37 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.215
+ $X2=1.55 $Y2=4.575
r161 32 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r162 32 35 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=3.215
r163 29 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r164 26 29 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.22
r165 9 65 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=4.575
r166 9 63 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.825 $X2=3.27 $Y2=3.215
r167 8 51 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.575
r168 8 49 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.215
r169 7 37 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.575
r170 7 35 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.215
r171 3 54 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.74
r172 2 40 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.74
r173 1 26 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

