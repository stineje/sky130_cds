* File: sky130_osu_sc_18T_ms__xnor2_l.pxi.spice
* Created: Fri Nov 12 14:07:33 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%GND N_GND_M1002_d N_GND_M1008_d N_GND_M1002_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_14_p N_GND_c_50_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_MS__XNOR2_L%GND
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%VDD N_VDD_M1004_d N_VDD_M1009_d N_VDD_M1004_b
+ N_VDD_c_74_p N_VDD_c_75_p N_VDD_c_71_p N_VDD_c_89_p N_VDD_c_91_p VDD
+ N_VDD_c_72_p PM_SKY130_OSU_SC_18T_MS__XNOR2_L%VDD
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%A N_A_c_110_n N_A_M1002_g N_A_M1004_g
+ N_A_c_114_n N_A_M1000_g N_A_M1007_g N_A_c_117_n N_A_c_118_n N_A_c_119_n
+ N_A_c_120_n N_A_c_121_n N_A_c_125_n N_A_c_126_n N_A_c_129_n N_A_c_130_n
+ N_A_c_145_p N_A_c_131_n A N_A_c_134_n PM_SKY130_OSU_SC_18T_MS__XNOR2_L%A
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1004_s N_A_27_115#_M1001_g N_A_27_115#_c_225_n
+ N_A_27_115#_M1006_g N_A_27_115#_c_228_n N_A_27_115#_c_229_n
+ N_A_27_115#_c_230_n N_A_27_115#_c_233_n N_A_27_115#_c_234_n
+ N_A_27_115#_c_235_n N_A_27_115#_c_236_n
+ PM_SKY130_OSU_SC_18T_MS__XNOR2_L%A_27_115#
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%A_238_89# N_A_238_89#_M1003_d
+ N_A_238_89#_M1005_d N_A_238_89#_M1010_g N_A_238_89#_M1011_g
+ N_A_238_89#_c_305_n N_A_238_89#_c_306_n N_A_238_89#_c_307_n
+ N_A_238_89#_c_309_n N_A_238_89#_c_310_n
+ PM_SKY130_OSU_SC_18T_MS__XNOR2_L%A_238_89#
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%B N_B_c_362_n N_B_M1008_g N_B_c_378_n
+ N_B_M1009_g N_B_c_366_n N_B_c_367_n N_B_c_368_n N_B_M1003_g N_B_c_371_n
+ N_B_c_385_n N_B_M1005_g N_B_c_372_n N_B_c_374_n N_B_c_375_n B
+ PM_SKY130_OSU_SC_18T_MS__XNOR2_L%B
x_PM_SKY130_OSU_SC_18T_MS__XNOR2_L%Y N_Y_M1010_d N_Y_M1011_d N_Y_c_418_n
+ N_Y_c_419_n N_Y_c_450_n N_Y_c_424_n N_Y_c_434_n Y N_Y_c_423_n N_Y_c_428_n
+ PM_SKY130_OSU_SC_18T_MS__XNOR2_L%Y
cc_1 N_GND_M1002_b N_A_c_110_n 0.0183137f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.65
cc_2 N_GND_c_2_p N_A_c_110_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.65
cc_3 N_GND_c_3_p N_A_c_110_n 0.00354579f $X=0.69 $Y=0.825 $X2=0.475 $Y2=1.65
cc_4 N_GND_c_4_p N_A_c_110_n 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=1.65
cc_5 N_GND_M1002_b N_A_c_114_n 0.00591749f $X=-0.045 $Y=0 $X2=0.71 $Y2=1.725
cc_6 N_GND_c_3_p N_A_c_114_n 0.00308996f $X=0.69 $Y=0.825 $X2=0.71 $Y2=1.725
cc_7 N_GND_M1002_b N_A_M1007_g 0.0214281f $X=-0.045 $Y=0 $X2=1.865 $Y2=4.585
cc_8 N_GND_M1002_b N_A_c_117_n 0.00962022f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.725
cc_9 N_GND_M1002_b N_A_c_118_n 0.0608283f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.86
cc_10 N_GND_M1002_b N_A_c_119_n 0.00432809f $X=-0.045 $Y=0 $X2=0.45 $Y2=3.01
cc_11 N_GND_M1002_b N_A_c_120_n 0.0240752f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.725
cc_12 N_GND_M1002_b N_A_c_121_n 0.0135251f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.65
cc_13 N_GND_c_3_p N_A_c_121_n 0.00354579f $X=0.69 $Y=0.825 $X2=0.845 $Y2=1.65
cc_14 N_GND_c_14_p N_A_c_121_n 0.00606474f $X=2.355 $Y=0.152 $X2=0.845 $Y2=1.65
cc_15 N_GND_c_4_p N_A_c_121_n 0.00468827f $X=2.38 $Y=0.19 $X2=0.845 $Y2=1.65
cc_16 N_GND_M1002_b N_A_c_125_n 0.052624f $X=-0.045 $Y=0 $X2=1.865 $Y2=2.405
cc_17 N_GND_M1002_d N_A_c_126_n 0.00190776f $X=0.55 $Y=0.575 $X2=0.845 $Y2=1.48
cc_18 N_GND_M1002_b N_A_c_126_n 0.00185864f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.48
cc_19 N_GND_c_3_p N_A_c_126_n 4.48624e-19 $X=0.69 $Y=0.825 $X2=0.845 $Y2=1.48
cc_20 N_GND_M1002_b N_A_c_129_n 0.00983735f $X=-0.045 $Y=0 $X2=2.145 $Y2=1.48
cc_21 N_GND_M1002_b N_A_c_130_n 0.00276199f $X=-0.045 $Y=0 $X2=2.225 $Y2=2.39
cc_22 N_GND_M1002_d N_A_c_131_n 0.00527794f $X=0.55 $Y=0.575 $X2=0.99 $Y2=1.48
cc_23 N_GND_M1002_b N_A_c_131_n 0.00167452f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.48
cc_24 N_GND_c_3_p N_A_c_131_n 0.00332581f $X=0.69 $Y=0.825 $X2=0.99 $Y2=1.48
cc_25 N_GND_M1002_b N_A_c_134_n 0.0024881f $X=-0.045 $Y=0 $X2=2.145 $Y2=1.48
cc_26 N_GND_M1002_b N_A_27_115#_M1001_g 0.0184711f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=4.585
cc_27 N_GND_M1002_b N_A_27_115#_c_225_n 0.0174779f $X=-0.045 $Y=0 $X2=1.865
+ $Y2=1.685
cc_28 N_GND_c_14_p N_A_27_115#_c_225_n 0.00606474f $X=2.355 $Y=0.152 $X2=1.865
+ $Y2=1.685
cc_29 N_GND_c_4_p N_A_27_115#_c_225_n 0.00468827f $X=2.38 $Y=0.19 $X2=1.865
+ $Y2=1.685
cc_30 N_GND_M1002_b N_A_27_115#_c_228_n 0.0277923f $X=-0.045 $Y=0 $X2=0.845
+ $Y2=2.39
cc_31 N_GND_M1002_b N_A_27_115#_c_229_n 0.0362346f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.85
cc_32 N_GND_M1002_b N_A_27_115#_c_230_n 0.0360665f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_33 N_GND_c_2_p N_A_27_115#_c_230_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_34 N_GND_c_4_p N_A_27_115#_c_230_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_35 N_GND_M1002_b N_A_27_115#_c_233_n 0.0201658f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.455
cc_36 N_GND_M1002_b N_A_27_115#_c_234_n 0.0354732f $X=-0.045 $Y=0 $X2=1.68
+ $Y2=2.39
cc_37 N_GND_M1002_b N_A_27_115#_c_235_n 0.00497247f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.85
cc_38 N_GND_M1002_b N_A_27_115#_c_236_n 0.00692367f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.39
cc_39 N_GND_M1002_b N_A_238_89#_M1010_g 0.0703714f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=1.075
cc_40 N_GND_c_14_p N_A_238_89#_M1010_g 0.00606474f $X=2.355 $Y=0.152 $X2=1.265
+ $Y2=1.075
cc_41 N_GND_c_4_p N_A_238_89#_M1010_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.265
+ $Y2=1.075
cc_42 N_GND_M1002_b N_A_238_89#_c_305_n 0.021482f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=2.765
cc_43 N_GND_M1002_b N_A_238_89#_c_306_n 0.0330247f $X=-0.045 $Y=0 $X2=2.785
+ $Y2=2.765
cc_44 N_GND_M1002_b N_A_238_89#_c_307_n 0.0612319f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=0.825
cc_45 N_GND_c_4_p N_A_238_89#_c_307_n 0.00476261f $X=2.38 $Y=0.19 $X2=2.87
+ $Y2=0.825
cc_46 N_GND_M1002_b N_A_238_89#_c_309_n 0.00243339f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=3.455
cc_47 N_GND_M1002_b N_A_238_89#_c_310_n 0.00720662f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=2.765
cc_48 N_GND_M1002_b N_B_c_362_n 0.0134938f $X=-0.045 $Y=0 $X2=2.225 $Y2=1.65
cc_49 N_GND_c_14_p N_B_c_362_n 0.00606474f $X=2.355 $Y=0.152 $X2=2.225 $Y2=1.65
cc_50 N_GND_c_50_p N_B_c_362_n 0.00354579f $X=2.44 $Y=0.825 $X2=2.225 $Y2=1.65
cc_51 N_GND_c_4_p N_B_c_362_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.225 $Y2=1.65
cc_52 N_GND_M1002_b N_B_c_366_n 0.00761231f $X=-0.045 $Y=0 $X2=2.58 $Y2=2.935
cc_53 N_GND_M1002_b N_B_c_367_n 0.00457156f $X=-0.045 $Y=0 $X2=2.3 $Y2=2.935
cc_54 N_GND_M1002_b N_B_c_368_n 0.0243862f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.65
cc_55 N_GND_c_50_p N_B_c_368_n 0.00354579f $X=2.44 $Y=0.825 $X2=2.655 $Y2=1.65
cc_56 N_GND_c_4_p N_B_c_368_n 0.00468827f $X=2.38 $Y=0.19 $X2=2.655 $Y2=1.65
cc_57 N_GND_M1002_b N_B_c_371_n 0.0472661f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.86
cc_58 N_GND_M1002_b N_B_c_372_n 0.0459817f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.832
cc_59 N_GND_c_50_p N_B_c_372_n 0.00243878f $X=2.44 $Y=0.825 $X2=2.655 $Y2=1.832
cc_60 N_GND_M1002_b N_B_c_374_n 0.00181559f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.935
cc_61 N_GND_M1002_b N_B_c_375_n 0.00227638f $X=-0.045 $Y=0 $X2=2.53 $Y2=1.85
cc_62 N_GND_c_50_p N_B_c_375_n 0.00234562f $X=2.44 $Y=0.825 $X2=2.53 $Y2=1.85
cc_63 N_GND_M1002_b B 0.00236483f $X=-0.045 $Y=0 $X2=2.53 $Y2=1.85
cc_64 N_GND_M1002_b N_Y_c_418_n 0.00785776f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.85
cc_65 N_GND_M1002_b N_Y_c_419_n 0.00313975f $X=-0.045 $Y=0 $X2=1.565 $Y2=0.825
cc_66 N_GND_c_14_p N_Y_c_419_n 0.0149397f $X=2.355 $Y=0.152 $X2=1.565 $Y2=0.825
cc_67 N_GND_c_4_p N_Y_c_419_n 0.00958198f $X=2.38 $Y=0.19 $X2=1.565 $Y2=0.825
cc_68 N_GND_M1002_b Y 0.00698114f $X=-0.045 $Y=0 $X2=1.42 $Y2=2.135
cc_69 N_GND_M1002_b N_Y_c_423_n 0.00238374f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.85
cc_70 N_VDD_M1004_b N_A_M1007_g 0.0215143f $X=-0.045 $Y=2.905 $X2=1.865
+ $Y2=4.585
cc_71 N_VDD_c_71_p N_A_M1007_g 0.00606474f $X=2.355 $Y=6.507 $X2=1.865 $Y2=4.585
cc_72 N_VDD_c_72_p N_A_M1007_g 0.00468827f $X=2.38 $Y=6.47 $X2=1.865 $Y2=4.585
cc_73 N_VDD_M1004_b N_A_c_119_n 0.0279802f $X=-0.045 $Y=2.905 $X2=0.45 $Y2=3.01
cc_74 N_VDD_c_74_p N_A_c_119_n 0.00606474f $X=0.605 $Y=6.507 $X2=0.45 $Y2=3.01
cc_75 N_VDD_c_75_p N_A_c_119_n 0.00354579f $X=0.69 $Y=3.455 $X2=0.45 $Y2=3.01
cc_76 N_VDD_c_72_p N_A_c_119_n 0.00468827f $X=2.38 $Y=6.47 $X2=0.45 $Y2=3.01
cc_77 N_VDD_M1004_b N_A_27_115#_M1001_g 0.0197604f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_78 N_VDD_c_75_p N_A_27_115#_M1001_g 0.00354579f $X=0.69 $Y=3.455 $X2=0.905
+ $Y2=4.585
cc_79 N_VDD_c_71_p N_A_27_115#_M1001_g 0.00606474f $X=2.355 $Y=6.507 $X2=0.905
+ $Y2=4.585
cc_80 N_VDD_c_72_p N_A_27_115#_M1001_g 0.00468827f $X=2.38 $Y=6.47 $X2=0.905
+ $Y2=4.585
cc_81 N_VDD_c_75_p N_A_27_115#_c_228_n 0.0017177f $X=0.69 $Y=3.455 $X2=0.845
+ $Y2=2.39
cc_82 N_VDD_M1004_b N_A_27_115#_c_233_n 0.0104815f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.455
cc_83 N_VDD_c_74_p N_A_27_115#_c_233_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=3.455
cc_84 N_VDD_c_72_p N_A_27_115#_c_233_n 0.00476261f $X=2.38 $Y=6.47 $X2=0.26
+ $Y2=3.455
cc_85 N_VDD_M1004_b N_A_238_89#_M1011_g 0.0192967f $X=-0.045 $Y=2.905 $X2=1.265
+ $Y2=4.585
cc_86 N_VDD_c_71_p N_A_238_89#_M1011_g 0.00606474f $X=2.355 $Y=6.507 $X2=1.265
+ $Y2=4.585
cc_87 N_VDD_c_72_p N_A_238_89#_M1011_g 0.00468827f $X=2.38 $Y=6.47 $X2=1.265
+ $Y2=4.585
cc_88 N_VDD_M1004_b N_A_238_89#_c_305_n 0.00559382f $X=-0.045 $Y=2.905 $X2=1.325
+ $Y2=2.765
cc_89 N_VDD_c_89_p N_A_238_89#_c_306_n 0.00811678f $X=2.44 $Y=3.455 $X2=2.785
+ $Y2=2.765
cc_90 N_VDD_M1004_b N_A_238_89#_c_309_n 0.00991954f $X=-0.045 $Y=2.905 $X2=2.87
+ $Y2=3.455
cc_91 N_VDD_c_91_p N_A_238_89#_c_309_n 0.00757793f $X=2.38 $Y=6.47 $X2=2.87
+ $Y2=3.455
cc_92 N_VDD_c_72_p N_A_238_89#_c_309_n 0.00476261f $X=2.38 $Y=6.47 $X2=2.87
+ $Y2=3.455
cc_93 N_VDD_M1004_b N_B_c_378_n 0.0139689f $X=-0.045 $Y=2.905 $X2=2.225 $Y2=3.01
cc_94 N_VDD_c_71_p N_B_c_378_n 0.00606474f $X=2.355 $Y=6.507 $X2=2.225 $Y2=3.01
cc_95 N_VDD_c_89_p N_B_c_378_n 0.00354579f $X=2.44 $Y=3.455 $X2=2.225 $Y2=3.01
cc_96 N_VDD_c_72_p N_B_c_378_n 0.00468827f $X=2.38 $Y=6.47 $X2=2.225 $Y2=3.01
cc_97 N_VDD_M1004_b N_B_c_366_n 0.00535962f $X=-0.045 $Y=2.905 $X2=2.58
+ $Y2=2.935
cc_98 N_VDD_c_89_p N_B_c_366_n 0.00221017f $X=2.44 $Y=3.455 $X2=2.58 $Y2=2.935
cc_99 N_VDD_M1004_b N_B_c_367_n 0.00345657f $X=-0.045 $Y=2.905 $X2=2.3 $Y2=2.935
cc_100 N_VDD_M1004_b N_B_c_385_n 0.0183291f $X=-0.045 $Y=2.905 $X2=2.655
+ $Y2=3.01
cc_101 N_VDD_c_89_p N_B_c_385_n 0.00354579f $X=2.44 $Y=3.455 $X2=2.655 $Y2=3.01
cc_102 N_VDD_c_91_p N_B_c_385_n 0.00606474f $X=2.38 $Y=6.47 $X2=2.655 $Y2=3.01
cc_103 N_VDD_c_72_p N_B_c_385_n 0.00468827f $X=2.38 $Y=6.47 $X2=2.655 $Y2=3.01
cc_104 N_VDD_M1004_b N_B_c_374_n 0.00423637f $X=-0.045 $Y=2.905 $X2=2.655
+ $Y2=2.935
cc_105 N_VDD_M1004_b N_Y_c_424_n 0.00313975f $X=-0.045 $Y=2.905 $X2=1.565
+ $Y2=3.455
cc_106 N_VDD_c_71_p N_Y_c_424_n 0.0149397f $X=2.355 $Y=6.507 $X2=1.565 $Y2=3.455
cc_107 N_VDD_c_72_p N_Y_c_424_n 0.00958198f $X=2.38 $Y=6.47 $X2=1.565 $Y2=3.455
cc_108 N_VDD_M1004_b Y 0.00321849f $X=-0.045 $Y=2.905 $X2=1.42 $Y2=2.135
cc_109 N_VDD_c_75_p N_Y_c_428_n 0.0045586f $X=0.69 $Y=3.455 $X2=1.425 $Y2=3.33
cc_110 N_A_c_118_n N_A_27_115#_M1001_g 0.0111858f $X=0.45 $Y=2.86 $X2=0.905
+ $Y2=4.585
cc_111 N_A_c_119_n N_A_27_115#_M1001_g 0.0245263f $X=0.45 $Y=3.01 $X2=0.905
+ $Y2=4.585
cc_112 N_A_c_129_n N_A_27_115#_c_225_n 0.00311835f $X=2.145 $Y=1.48 $X2=1.865
+ $Y2=1.685
cc_113 N_A_c_145_p N_A_27_115#_c_225_n 0.0134125f $X=2 $Y=1.48 $X2=1.865
+ $Y2=1.685
cc_114 N_A_c_134_n N_A_27_115#_c_225_n 9.56269e-19 $X=2.145 $Y=1.48 $X2=1.865
+ $Y2=1.685
cc_115 N_A_c_118_n N_A_27_115#_c_228_n 0.0212638f $X=0.45 $Y=2.86 $X2=0.845
+ $Y2=2.39
cc_116 N_A_c_120_n N_A_27_115#_c_228_n 0.0184269f $X=0.845 $Y=1.725 $X2=0.845
+ $Y2=2.39
cc_117 N_A_c_126_n N_A_27_115#_c_228_n 6.74966e-19 $X=0.845 $Y=1.48 $X2=0.845
+ $Y2=2.39
cc_118 N_A_c_131_n N_A_27_115#_c_228_n 4.48459e-19 $X=0.99 $Y=1.48 $X2=0.845
+ $Y2=2.39
cc_119 N_A_c_125_n N_A_27_115#_c_229_n 0.00515091f $X=1.865 $Y=2.405 $X2=1.765
+ $Y2=1.85
cc_120 N_A_c_129_n N_A_27_115#_c_229_n 0.00194908f $X=2.145 $Y=1.48 $X2=1.765
+ $Y2=1.85
cc_121 N_A_c_145_p N_A_27_115#_c_229_n 0.00130191f $X=2 $Y=1.48 $X2=1.765
+ $Y2=1.85
cc_122 N_A_c_110_n N_A_27_115#_c_230_n 0.00703867f $X=0.475 $Y=1.65 $X2=0.26
+ $Y2=0.825
cc_123 N_A_c_117_n N_A_27_115#_c_230_n 0.022872f $X=0.45 $Y=1.725 $X2=0.26
+ $Y2=0.825
cc_124 N_A_c_126_n N_A_27_115#_c_230_n 0.0184292f $X=0.845 $Y=1.48 $X2=0.26
+ $Y2=0.825
cc_125 N_A_c_131_n N_A_27_115#_c_230_n 0.00710152f $X=0.99 $Y=1.48 $X2=0.26
+ $Y2=0.825
cc_126 N_A_c_118_n N_A_27_115#_c_233_n 0.0221084f $X=0.45 $Y=2.86 $X2=0.26
+ $Y2=3.455
cc_127 N_A_c_119_n N_A_27_115#_c_233_n 0.00727773f $X=0.45 $Y=3.01 $X2=0.26
+ $Y2=3.455
cc_128 N_A_c_114_n N_A_27_115#_c_234_n 8.76512e-19 $X=0.71 $Y=1.725 $X2=1.68
+ $Y2=2.39
cc_129 N_A_c_118_n N_A_27_115#_c_234_n 0.0199699f $X=0.45 $Y=2.86 $X2=1.68
+ $Y2=2.39
cc_130 N_A_c_119_n N_A_27_115#_c_234_n 0.00165231f $X=0.45 $Y=3.01 $X2=1.68
+ $Y2=2.39
cc_131 N_A_c_120_n N_A_27_115#_c_234_n 8.34298e-19 $X=0.845 $Y=1.725 $X2=1.68
+ $Y2=2.39
cc_132 N_A_c_125_n N_A_27_115#_c_234_n 0.00528869f $X=1.865 $Y=2.405 $X2=1.68
+ $Y2=2.39
cc_133 N_A_c_126_n N_A_27_115#_c_234_n 0.00826927f $X=0.845 $Y=1.48 $X2=1.68
+ $Y2=2.39
cc_134 N_A_c_130_n N_A_27_115#_c_234_n 0.0116688f $X=2.225 $Y=2.39 $X2=1.68
+ $Y2=2.39
cc_135 N_A_c_125_n N_A_27_115#_c_235_n 5.00447e-19 $X=1.865 $Y=2.405 $X2=1.765
+ $Y2=1.85
cc_136 N_A_c_129_n N_A_27_115#_c_235_n 0.0360591f $X=2.145 $Y=1.48 $X2=1.765
+ $Y2=1.85
cc_137 N_A_c_145_p N_A_27_115#_c_235_n 0.00737704f $X=2 $Y=1.48 $X2=1.765
+ $Y2=1.85
cc_138 N_A_c_118_n N_A_238_89#_M1010_g 0.00462097f $X=0.45 $Y=2.86 $X2=1.265
+ $Y2=1.075
cc_139 N_A_c_121_n N_A_238_89#_M1010_g 0.0961644f $X=0.845 $Y=1.65 $X2=1.265
+ $Y2=1.075
cc_140 N_A_c_125_n N_A_238_89#_M1010_g 0.00525031f $X=1.865 $Y=2.405 $X2=1.265
+ $Y2=1.075
cc_141 N_A_c_126_n N_A_238_89#_M1010_g 0.00228168f $X=0.845 $Y=1.48 $X2=1.265
+ $Y2=1.075
cc_142 N_A_c_145_p N_A_238_89#_M1010_g 0.0133678f $X=2 $Y=1.48 $X2=1.265
+ $Y2=1.075
cc_143 N_A_c_131_n N_A_238_89#_M1010_g 8.6716e-19 $X=0.99 $Y=1.48 $X2=1.265
+ $Y2=1.075
cc_144 N_A_M1007_g N_A_238_89#_M1011_g 0.0616724f $X=1.865 $Y=4.585 $X2=1.265
+ $Y2=4.585
cc_145 N_A_M1007_g N_A_238_89#_c_305_n 0.0126871f $X=1.865 $Y=4.585 $X2=1.325
+ $Y2=2.765
cc_146 N_A_M1007_g N_A_238_89#_c_306_n 0.018341f $X=1.865 $Y=4.585 $X2=2.785
+ $Y2=2.765
cc_147 N_A_c_125_n N_A_238_89#_c_306_n 0.00796541f $X=1.865 $Y=2.405 $X2=2.785
+ $Y2=2.765
cc_148 N_A_c_130_n N_A_238_89#_c_306_n 0.0206305f $X=2.225 $Y=2.39 $X2=2.785
+ $Y2=2.765
cc_149 N_A_c_129_n N_A_238_89#_c_307_n 0.0132855f $X=2.145 $Y=1.48 $X2=2.87
+ $Y2=0.825
cc_150 N_A_c_130_n N_A_238_89#_c_307_n 0.00742262f $X=2.225 $Y=2.39 $X2=2.87
+ $Y2=0.825
cc_151 N_A_c_134_n N_A_238_89#_c_307_n 0.00547471f $X=2.145 $Y=1.48 $X2=2.87
+ $Y2=0.825
cc_152 N_A_c_129_n N_B_c_362_n 0.00753906f $X=2.145 $Y=1.48 $X2=2.225 $Y2=1.65
cc_153 N_A_c_134_n N_B_c_362_n 0.00991486f $X=2.145 $Y=1.48 $X2=2.225 $Y2=1.65
cc_154 N_A_M1007_g N_B_c_367_n 0.199321f $X=1.865 $Y=4.585 $X2=2.3 $Y2=2.935
cc_155 N_A_c_125_n N_B_c_367_n 0.00779298f $X=1.865 $Y=2.405 $X2=2.3 $Y2=2.935
cc_156 N_A_c_129_n N_B_c_368_n 0.00106222f $X=2.145 $Y=1.48 $X2=2.655 $Y2=1.65
cc_157 N_A_c_134_n N_B_c_368_n 0.00122438f $X=2.145 $Y=1.48 $X2=2.655 $Y2=1.65
cc_158 N_A_M1007_g N_B_c_371_n 0.00402444f $X=1.865 $Y=4.585 $X2=2.655 $Y2=2.86
cc_159 N_A_c_125_n N_B_c_371_n 0.0193201f $X=1.865 $Y=2.405 $X2=2.655 $Y2=2.86
cc_160 N_A_c_129_n N_B_c_371_n 0.00243832f $X=2.145 $Y=1.48 $X2=2.655 $Y2=2.86
cc_161 N_A_c_130_n N_B_c_371_n 0.00131152f $X=2.225 $Y=2.39 $X2=2.655 $Y2=2.86
cc_162 N_A_c_125_n N_B_c_372_n 0.00620704f $X=1.865 $Y=2.405 $X2=2.655 $Y2=1.832
cc_163 N_A_c_129_n N_B_c_372_n 0.00728935f $X=2.145 $Y=1.48 $X2=2.655 $Y2=1.832
cc_164 N_A_c_130_n N_B_c_372_n 0.00132282f $X=2.225 $Y=2.39 $X2=2.655 $Y2=1.832
cc_165 N_A_c_129_n N_B_c_375_n 0.0165474f $X=2.145 $Y=1.48 $X2=2.53 $Y2=1.85
cc_166 N_A_c_125_n B 0.00116112f $X=1.865 $Y=2.405 $X2=2.53 $Y2=1.85
cc_167 N_A_c_129_n B 0.007568f $X=2.145 $Y=1.48 $X2=2.53 $Y2=1.85
cc_168 N_A_c_130_n B 0.00408329f $X=2.225 $Y=2.39 $X2=2.53 $Y2=1.85
cc_169 N_A_c_134_n B 0.00136805f $X=2.145 $Y=1.48 $X2=2.53 $Y2=1.85
cc_170 N_A_c_145_p N_Y_M1010_d 0.00659511f $X=2 $Y=1.48 $X2=1.34 $Y2=0.575
cc_171 N_A_c_129_n N_Y_c_418_n 0.00604346f $X=2.145 $Y=1.48 $X2=1.425 $Y2=1.85
cc_172 N_A_c_145_p N_Y_c_418_n 0.0114959f $X=2 $Y=1.48 $X2=1.425 $Y2=1.85
cc_173 N_A_c_131_n N_Y_c_418_n 7.8621e-19 $X=0.99 $Y=1.48 $X2=1.425 $Y2=1.85
cc_174 N_A_c_134_n N_Y_c_418_n 7.10974e-19 $X=2.145 $Y=1.48 $X2=1.425 $Y2=1.85
cc_175 N_A_c_126_n N_Y_c_434_n 0.0136175f $X=0.845 $Y=1.48 $X2=1.537 $Y2=1.415
cc_176 N_A_c_129_n N_Y_c_434_n 5.37889e-19 $X=2.145 $Y=1.48 $X2=1.537 $Y2=1.415
cc_177 N_A_c_145_p N_Y_c_434_n 0.027218f $X=2 $Y=1.48 $X2=1.537 $Y2=1.415
cc_178 N_A_c_131_n N_Y_c_434_n 0.00133183f $X=0.99 $Y=1.48 $X2=1.537 $Y2=1.415
cc_179 N_A_c_134_n N_Y_c_434_n 0.00144576f $X=2.145 $Y=1.48 $X2=1.537 $Y2=1.415
cc_180 N_A_c_120_n Y 2.24638e-19 $X=0.845 $Y=1.725 $X2=1.42 $Y2=2.135
cc_181 N_A_c_125_n Y 0.00743805f $X=1.865 $Y=2.405 $X2=1.42 $Y2=2.135
cc_182 N_A_c_126_n Y 0.00146257f $X=0.845 $Y=1.48 $X2=1.42 $Y2=2.135
cc_183 N_A_c_130_n Y 6.70937e-19 $X=2.225 $Y=2.39 $X2=1.42 $Y2=2.135
cc_184 N_A_c_120_n N_Y_c_423_n 0.0011785f $X=0.845 $Y=1.725 $X2=1.425 $Y2=1.85
cc_185 N_A_c_126_n N_Y_c_423_n 0.00531647f $X=0.845 $Y=1.48 $X2=1.425 $Y2=1.85
cc_186 N_A_c_145_p N_Y_c_423_n 0.0259322f $X=2 $Y=1.48 $X2=1.425 $Y2=1.85
cc_187 N_A_c_145_p A_196_115# 0.015419f $X=2 $Y=1.48 $X2=0.98 $Y2=0.575
cc_188 N_A_c_131_n A_196_115# 8.19673e-19 $X=0.99 $Y=1.48 $X2=0.98 $Y2=0.575
cc_189 N_A_c_129_n A_388_115# 0.00262479f $X=2.145 $Y=1.48 $X2=1.94 $Y2=0.575
cc_190 N_A_c_145_p A_388_115# 0.00457146f $X=2 $Y=1.48 $X2=1.94 $Y2=0.575
cc_191 N_A_c_134_n A_388_115# 0.00638831f $X=2.145 $Y=1.48 $X2=1.94 $Y2=0.575
cc_192 N_A_27_115#_c_225_n N_A_238_89#_M1010_g 0.0253069f $X=1.865 $Y=1.685
+ $X2=1.265 $Y2=1.075
cc_193 N_A_27_115#_c_228_n N_A_238_89#_M1010_g 0.119517f $X=0.845 $Y=2.39
+ $X2=1.265 $Y2=1.075
cc_194 N_A_27_115#_c_229_n N_A_238_89#_M1010_g 0.0141925f $X=1.765 $Y=1.85
+ $X2=1.265 $Y2=1.075
cc_195 N_A_27_115#_c_234_n N_A_238_89#_M1010_g 0.0146245f $X=1.68 $Y=2.39
+ $X2=1.265 $Y2=1.075
cc_196 N_A_27_115#_c_235_n N_A_238_89#_M1010_g 0.00755502f $X=1.765 $Y=1.85
+ $X2=1.265 $Y2=1.075
cc_197 N_A_27_115#_M1001_g N_A_238_89#_c_305_n 0.119517f $X=0.905 $Y=4.585
+ $X2=1.325 $Y2=2.765
cc_198 N_A_27_115#_c_234_n N_A_238_89#_c_305_n 0.00220335f $X=1.68 $Y=2.39
+ $X2=1.325 $Y2=2.765
cc_199 N_A_27_115#_M1001_g N_A_238_89#_c_306_n 0.00444529f $X=0.905 $Y=4.585
+ $X2=2.785 $Y2=2.765
cc_200 N_A_27_115#_c_229_n N_A_238_89#_c_306_n 6.30959e-19 $X=1.765 $Y=1.85
+ $X2=2.785 $Y2=2.765
cc_201 N_A_27_115#_c_234_n N_A_238_89#_c_306_n 0.0436145f $X=1.68 $Y=2.39
+ $X2=2.785 $Y2=2.765
cc_202 N_A_27_115#_c_225_n N_B_c_362_n 0.0413157f $X=1.865 $Y=1.685 $X2=2.225
+ $Y2=1.65
cc_203 N_A_27_115#_c_229_n N_B_c_372_n 0.0456843f $X=1.765 $Y=1.85 $X2=2.655
+ $Y2=1.832
cc_204 N_A_27_115#_c_225_n N_Y_c_418_n 0.00208671f $X=1.865 $Y=1.685 $X2=1.425
+ $Y2=1.85
cc_205 N_A_27_115#_c_229_n N_Y_c_418_n 0.00161977f $X=1.765 $Y=1.85 $X2=1.425
+ $Y2=1.85
cc_206 N_A_27_115#_c_234_n N_Y_c_418_n 0.00556015f $X=1.68 $Y=2.39 $X2=1.425
+ $Y2=1.85
cc_207 N_A_27_115#_c_235_n N_Y_c_418_n 0.0159901f $X=1.765 $Y=1.85 $X2=1.425
+ $Y2=1.85
cc_208 N_A_27_115#_M1001_g N_Y_c_450_n 7.92921e-19 $X=0.905 $Y=4.585 $X2=1.565
+ $Y2=3.445
cc_209 N_A_27_115#_c_225_n N_Y_c_434_n 0.00531991f $X=1.865 $Y=1.685 $X2=1.537
+ $Y2=1.415
cc_210 N_A_27_115#_c_229_n N_Y_c_434_n 0.00194835f $X=1.765 $Y=1.85 $X2=1.537
+ $Y2=1.415
cc_211 N_A_27_115#_c_235_n N_Y_c_434_n 0.00214832f $X=1.765 $Y=1.85 $X2=1.537
+ $Y2=1.415
cc_212 N_A_27_115#_M1001_g Y 0.00191867f $X=0.905 $Y=4.585 $X2=1.42 $Y2=2.135
cc_213 N_A_27_115#_c_228_n Y 9.27207e-19 $X=0.845 $Y=2.39 $X2=1.42 $Y2=2.135
cc_214 N_A_27_115#_c_229_n Y 7.0267e-19 $X=1.765 $Y=1.85 $X2=1.42 $Y2=2.135
cc_215 N_A_27_115#_c_234_n Y 0.0160336f $X=1.68 $Y=2.39 $X2=1.42 $Y2=2.135
cc_216 N_A_27_115#_c_235_n Y 0.015499f $X=1.765 $Y=1.85 $X2=1.42 $Y2=2.135
cc_217 N_A_27_115#_c_229_n N_Y_c_423_n 0.00394131f $X=1.765 $Y=1.85 $X2=1.425
+ $Y2=1.85
cc_218 N_A_27_115#_c_234_n N_Y_c_423_n 0.00440188f $X=1.68 $Y=2.39 $X2=1.425
+ $Y2=1.85
cc_219 N_A_27_115#_c_235_n N_Y_c_423_n 0.00746221f $X=1.765 $Y=1.85 $X2=1.425
+ $Y2=1.85
cc_220 N_A_27_115#_M1001_g N_Y_c_428_n 0.00108503f $X=0.905 $Y=4.585 $X2=1.425
+ $Y2=3.33
cc_221 N_A_238_89#_c_306_n N_B_c_367_n 0.0133212f $X=2.785 $Y=2.765 $X2=2.3
+ $Y2=2.935
cc_222 N_A_238_89#_c_307_n N_B_c_368_n 0.0378987f $X=2.87 $Y=0.825 $X2=2.655
+ $Y2=1.65
cc_223 N_A_238_89#_c_306_n N_B_c_371_n 0.020054f $X=2.785 $Y=2.765 $X2=2.655
+ $Y2=2.86
cc_224 N_A_238_89#_c_309_n N_B_c_371_n 0.0145613f $X=2.87 $Y=3.455 $X2=2.655
+ $Y2=2.86
cc_225 N_A_238_89#_c_306_n N_B_c_372_n 0.00180943f $X=2.785 $Y=2.765 $X2=2.655
+ $Y2=1.832
cc_226 N_A_238_89#_c_306_n N_B_c_375_n 0.00433845f $X=2.785 $Y=2.765 $X2=2.53
+ $Y2=1.85
cc_227 N_A_238_89#_c_307_n N_B_c_375_n 0.0214571f $X=2.87 $Y=0.825 $X2=2.53
+ $Y2=1.85
cc_228 N_A_238_89#_c_307_n B 0.00642833f $X=2.87 $Y=0.825 $X2=2.53 $Y2=1.85
cc_229 N_A_238_89#_M1011_g N_Y_c_450_n 0.0034761f $X=1.265 $Y=4.585 $X2=1.565
+ $Y2=3.445
cc_230 N_A_238_89#_c_305_n N_Y_c_450_n 0.00170549f $X=1.325 $Y=2.765 $X2=1.565
+ $Y2=3.445
cc_231 N_A_238_89#_c_306_n N_Y_c_450_n 0.015078f $X=2.785 $Y=2.765 $X2=1.565
+ $Y2=3.445
cc_232 N_A_238_89#_M1010_g N_Y_c_434_n 0.00684302f $X=1.265 $Y=1.075 $X2=1.537
+ $Y2=1.415
cc_233 N_A_238_89#_M1010_g Y 0.00982251f $X=1.265 $Y=1.075 $X2=1.42 $Y2=2.135
cc_234 N_A_238_89#_M1011_g Y 0.00464698f $X=1.265 $Y=4.585 $X2=1.42 $Y2=2.135
cc_235 N_A_238_89#_c_305_n Y 0.00651733f $X=1.325 $Y=2.765 $X2=1.42 $Y2=2.135
cc_236 N_A_238_89#_c_306_n Y 0.0165306f $X=2.785 $Y=2.765 $X2=1.42 $Y2=2.135
cc_237 N_A_238_89#_M1010_g N_Y_c_423_n 0.00425916f $X=1.265 $Y=1.075 $X2=1.425
+ $Y2=1.85
cc_238 N_A_238_89#_M1011_g N_Y_c_428_n 0.00624758f $X=1.265 $Y=4.585 $X2=1.425
+ $Y2=3.33
cc_239 N_A_238_89#_c_306_n N_Y_c_428_n 0.00233457f $X=2.785 $Y=2.765 $X2=1.425
+ $Y2=3.33
