magic
tech sky130A
magscale 1 2
timestamp 1606864608
<< checkpaint >>
rect -1209 -1243 1617 2575
<< nwell >>
rect -9 581 462 1341
<< nmos >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
rect 338 115 368 315
<< pmos >>
rect 80 617 110 1217
rect 152 617 182 1217
rect 252 617 282 1217
rect 324 617 354 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 199 166 315
rect 110 131 121 199
rect 155 131 166 199
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 267 338 315
rect 282 199 293 267
rect 327 199 338 267
rect 282 115 338 199
rect 368 199 421 315
rect 368 131 379 199
rect 413 131 421 199
rect 368 115 421 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 617 152 1217
rect 182 1201 252 1217
rect 182 725 200 1201
rect 234 725 252 1201
rect 182 617 252 725
rect 282 617 324 1217
rect 354 1201 407 1217
rect 354 793 365 1201
rect 399 793 407 1201
rect 354 617 407 793
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 199
rect 207 131 241 267
rect 293 199 327 267
rect 379 131 413 199
<< pdiffc >>
rect 35 793 69 1201
rect 200 725 234 1201
rect 365 793 399 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
<< poly >>
rect 80 1217 110 1243
rect 152 1217 182 1243
rect 252 1217 282 1243
rect 324 1217 354 1243
rect 80 585 110 617
rect 56 569 110 585
rect 56 535 66 569
rect 100 535 110 569
rect 56 519 110 535
rect 56 370 86 519
rect 152 471 182 617
rect 130 461 196 471
rect 130 427 146 461
rect 180 427 196 461
rect 130 417 196 427
rect 56 340 110 370
rect 80 315 110 340
rect 166 315 196 417
rect 252 409 282 617
rect 324 592 354 617
rect 324 562 368 592
rect 338 478 368 562
rect 338 462 430 478
rect 338 428 384 462
rect 418 428 430 462
rect 338 412 430 428
rect 238 393 292 409
rect 238 359 248 393
rect 282 359 292 393
rect 238 343 292 359
rect 252 315 282 343
rect 338 315 368 412
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
rect 338 89 368 115
<< polycont >>
rect 66 535 100 569
rect 146 427 180 461
rect 384 428 418 462
rect 248 359 282 393
<< locali >>
rect 0 1311 462 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 462 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 200 1201 234 1217
rect 365 1201 399 1271
rect 365 777 399 793
rect 200 700 234 725
rect 200 666 350 700
rect 66 569 100 649
rect 66 519 100 535
rect 146 575 162 609
rect 146 461 180 575
rect 146 411 180 427
rect 223 409 257 501
rect 223 393 282 409
rect 223 359 248 393
rect 223 343 282 359
rect 316 387 350 666
rect 384 462 418 478
rect 384 412 418 428
rect 35 267 241 301
rect 35 115 69 131
rect 121 199 155 215
rect 121 61 155 131
rect 293 279 316 283
rect 293 267 350 279
rect 327 249 350 267
rect 293 183 327 199
rect 379 199 413 215
rect 241 131 379 149
rect 207 115 413 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 462 61
rect 0 0 462 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 66 649 100 683
rect 162 575 196 609
rect 223 501 257 535
rect 384 428 418 462
rect 316 353 350 387
rect 316 279 350 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
<< metal1 >>
rect 0 1311 462 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 462 1311
rect 0 1271 462 1277
rect 54 683 112 689
rect 54 649 66 683
rect 100 649 134 683
rect 54 643 112 649
rect 150 609 208 615
rect 150 575 162 609
rect 196 575 230 609
rect 150 569 208 575
rect 211 535 269 541
rect 189 501 223 535
rect 257 501 269 535
rect 211 495 269 501
rect 372 462 430 468
rect 350 428 384 462
rect 418 428 430 462
rect 372 422 430 428
rect 304 387 362 393
rect 304 353 316 387
rect 350 353 362 387
rect 304 347 362 353
rect 316 319 350 347
rect 304 313 362 319
rect 304 279 316 313
rect 350 279 362 313
rect 304 273 362 279
rect 0 55 462 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 462 55
rect 0 0 462 21
<< labels >>
rlabel metal1 240 518 240 518 1 B0
port 4 n
rlabel viali 179 592 179 592 1 A1
port 2 n
rlabel viali 83 666 83 666 1 A0
port 1 n
rlabel viali 333 370 333 370 1 Y
port 3 n
rlabel viali 401 445 401 445 1 B1
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
