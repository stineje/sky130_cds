* File: sky130_osu_sc_18T_ms__and2_6.pxi.spice
* Created: Thu Oct 29 17:27:33 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__AND2_6%noxref_1 N_noxref_1_M1002_d N_noxref_1_M1006_s
+ N_noxref_1_M1010_s N_noxref_1_M1014_s N_noxref_1_M1004_b N_noxref_1_c_2_p
+ N_noxref_1_c_7_p N_noxref_1_c_14_p N_noxref_1_c_20_p N_noxref_1_c_26_p
+ N_noxref_1_c_31_p N_noxref_1_c_37_p N_noxref_1_c_43_p N_noxref_1_c_99_p
+ N_noxref_1_c_100_p PM_SKY130_OSU_SC_18T_MS__AND2_6%noxref_1
x_PM_SKY130_OSU_SC_18T_MS__AND2_6%noxref_2 N_noxref_2_M1005_s N_noxref_2_M1000_d
+ N_noxref_2_M1007_s N_noxref_2_M1011_s N_noxref_2_M1015_s N_noxref_2_M1005_b
+ N_noxref_2_c_160_p N_noxref_2_c_102_p N_noxref_2_c_103_p N_noxref_2_c_113_p
+ N_noxref_2_c_119_p N_noxref_2_c_124_p N_noxref_2_c_129_p N_noxref_2_c_133_p
+ N_noxref_2_c_138_p N_noxref_2_c_142_p N_noxref_2_c_165_p N_noxref_2_c_166_p
+ N_noxref_2_c_167_p PM_SKY130_OSU_SC_18T_MS__AND2_6%noxref_2
x_PM_SKY130_OSU_SC_18T_MS__AND2_6%A N_A_M1004_g N_A_M1005_g A N_A_c_170_n
+ N_A_c_171_n PM_SKY130_OSU_SC_18T_MS__AND2_6%A
x_PM_SKY130_OSU_SC_18T_MS__AND2_6%B N_B_M1002_g N_B_M1000_g B N_B_c_202_n
+ N_B_c_203_n PM_SKY130_OSU_SC_18T_MS__AND2_6%B
x_PM_SKY130_OSU_SC_18T_MS__AND2_6%A_27_115# N_A_27_115#_M1004_s
+ N_A_27_115#_M1005_d N_A_27_115#_M1001_g N_A_27_115#_c_238_n
+ N_A_27_115#_c_283_n N_A_27_115#_M1003_g N_A_27_115#_c_239_n
+ N_A_27_115#_c_240_n N_A_27_115#_M1006_g N_A_27_115#_c_287_n
+ N_A_27_115#_M1007_g N_A_27_115#_c_244_n N_A_27_115#_c_246_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_293_n N_A_27_115#_M1009_g
+ N_A_27_115#_c_250_n N_A_27_115#_c_251_n N_A_27_115#_M1010_g
+ N_A_27_115#_c_297_n N_A_27_115#_M1011_g N_A_27_115#_c_255_n
+ N_A_27_115#_c_257_n N_A_27_115#_M1012_g N_A_27_115#_c_261_n
+ N_A_27_115#_c_302_n N_A_27_115#_M1013_g N_A_27_115#_c_262_n
+ N_A_27_115#_c_263_n N_A_27_115#_M1014_g N_A_27_115#_c_306_n
+ N_A_27_115#_M1015_g N_A_27_115#_c_267_n N_A_27_115#_c_268_n
+ N_A_27_115#_c_269_n N_A_27_115#_c_270_n N_A_27_115#_c_271_n
+ N_A_27_115#_c_272_n N_A_27_115#_c_273_n N_A_27_115#_c_274_n
+ N_A_27_115#_c_275_n N_A_27_115#_c_276_n N_A_27_115#_c_278_n
+ N_A_27_115#_c_315_n N_A_27_115#_c_279_n N_A_27_115#_c_280_n
+ N_A_27_115#_c_326_n N_A_27_115#_c_282_n
+ PM_SKY130_OSU_SC_18T_MS__AND2_6%A_27_115#
x_PM_SKY130_OSU_SC_18T_MS__AND2_6%Y N_Y_M1001_d N_Y_M1008_d N_Y_M1012_d
+ N_Y_M1003_d N_Y_M1009_d N_Y_M1013_d N_Y_c_423_n N_Y_c_426_n Y N_Y_c_428_n
+ N_Y_c_430_n N_Y_c_431_n N_Y_c_432_n N_Y_c_434_n N_Y_c_437_n N_Y_c_438_n
+ N_Y_c_439_n N_Y_c_442_n N_Y_c_443_n N_Y_c_444_n N_Y_c_445_n N_Y_c_446_n
+ N_Y_c_450_n N_Y_c_454_n PM_SKY130_OSU_SC_18T_MS__AND2_6%Y
cc_1 N_noxref_1_M1004_b N_A_M1004_g 0.0805447f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=1.075
cc_2 N_noxref_1_c_2_p N_A_M1004_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475
+ $Y2=1.075
cc_3 N_noxref_1_M1004_b N_A_c_170_n 0.00329519f $X=-0.045 $Y=0 $X2=0.235
+ $Y2=2.765
cc_4 N_noxref_1_M1004_b N_A_c_171_n 0.0447183f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=2.765
cc_5 N_noxref_1_M1004_b N_B_M1002_g 0.0456699f $X=-0.045 $Y=0 $X2=0.835
+ $Y2=1.075
cc_6 N_noxref_1_c_2_p N_B_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835
+ $Y2=1.075
cc_7 N_noxref_1_c_7_p N_B_M1002_g 0.00376152f $X=1.05 $Y=0.825 $X2=0.835
+ $Y2=1.075
cc_8 N_noxref_1_M1004_b N_B_M1000_g 0.0145087f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=4.585
cc_9 N_noxref_1_M1004_b B 0.00685421f $X=-0.045 $Y=0 $X2=0.92 $Y2=2.96
cc_10 N_noxref_1_M1004_b N_B_c_202_n 0.00352155f $X=-0.045 $Y=0 $X2=0.915
+ $Y2=2.425
cc_11 N_noxref_1_M1004_b N_B_c_203_n 0.0304191f $X=-0.045 $Y=0 $X2=0.915
+ $Y2=2.425
cc_12 N_noxref_1_M1004_b N_A_27_115#_M1001_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_13 N_noxref_1_c_7_p N_A_27_115#_M1001_g 0.0103278f $X=1.05 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_14 N_noxref_1_c_14_p N_A_27_115#_M1001_g 0.00606474f $X=1.895 $Y=0.152
+ $X2=1.335 $Y2=1.075
cc_15 N_noxref_1_M1004_b N_A_27_115#_c_238_n 0.0465667f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=2.81
cc_16 N_noxref_1_M1004_b N_A_27_115#_c_239_n 0.00863342f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.885
cc_17 N_noxref_1_M1004_b N_A_27_115#_c_240_n 0.0104564f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.845
cc_18 N_noxref_1_M1004_b N_A_27_115#_M1006_g 0.0202142f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_19 N_noxref_1_c_14_p N_A_27_115#_M1006_g 0.00606474f $X=1.895 $Y=0.152
+ $X2=1.765 $Y2=1.075
cc_20 N_noxref_1_c_20_p N_A_27_115#_M1006_g 0.00356864f $X=1.98 $Y=0.825
+ $X2=1.765 $Y2=1.075
cc_21 N_noxref_1_M1004_b N_A_27_115#_c_244_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.845
cc_22 N_noxref_1_c_20_p N_A_27_115#_c_244_n 0.00256938f $X=1.98 $Y=0.825
+ $X2=2.12 $Y2=1.845
cc_23 N_noxref_1_M1004_b N_A_27_115#_c_246_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.885
cc_24 N_noxref_1_M1004_b N_A_27_115#_M1008_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.075
cc_25 N_noxref_1_c_20_p N_A_27_115#_M1008_g 0.00356864f $X=1.98 $Y=0.825
+ $X2=2.195 $Y2=1.075
cc_26 N_noxref_1_c_26_p N_A_27_115#_M1008_g 0.00606474f $X=2.755 $Y=0.152
+ $X2=2.195 $Y2=1.075
cc_27 N_noxref_1_M1004_b N_A_27_115#_c_250_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.845
cc_28 N_noxref_1_M1004_b N_A_27_115#_c_251_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.885
cc_29 N_noxref_1_M1004_b N_A_27_115#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.075
cc_30 N_noxref_1_c_26_p N_A_27_115#_M1010_g 0.00606474f $X=2.755 $Y=0.152
+ $X2=2.625 $Y2=1.075
cc_31 N_noxref_1_c_31_p N_A_27_115#_M1010_g 0.00356864f $X=2.84 $Y=0.825
+ $X2=2.625 $Y2=1.075
cc_32 N_noxref_1_M1004_b N_A_27_115#_c_255_n 0.0181078f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.845
cc_33 N_noxref_1_c_31_p N_A_27_115#_c_255_n 0.00256938f $X=2.84 $Y=0.825
+ $X2=2.98 $Y2=1.845
cc_34 N_noxref_1_M1004_b N_A_27_115#_c_257_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.885
cc_35 N_noxref_1_M1004_b N_A_27_115#_M1012_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.075
cc_36 N_noxref_1_c_31_p N_A_27_115#_M1012_g 0.00356864f $X=2.84 $Y=0.825
+ $X2=3.055 $Y2=1.075
cc_37 N_noxref_1_c_37_p N_A_27_115#_M1012_g 0.00606474f $X=3.615 $Y=0.152
+ $X2=3.055 $Y2=1.075
cc_38 N_noxref_1_M1004_b N_A_27_115#_c_261_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.81
cc_39 N_noxref_1_M1004_b N_A_27_115#_c_262_n 0.0369419f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.845
cc_40 N_noxref_1_M1004_b N_A_27_115#_c_263_n 0.0268552f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.885
cc_41 N_noxref_1_M1004_b N_A_27_115#_M1014_g 0.0264941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.075
cc_42 N_noxref_1_c_37_p N_A_27_115#_M1014_g 0.00606474f $X=3.615 $Y=0.152
+ $X2=3.485 $Y2=1.075
cc_43 N_noxref_1_c_43_p N_A_27_115#_M1014_g 0.00713292f $X=3.7 $Y=0.825
+ $X2=3.485 $Y2=1.075
cc_44 N_noxref_1_M1004_b N_A_27_115#_c_267_n 0.00339913f $X=-0.045 $Y=0
+ $X2=1.335 $Y2=2.885
cc_45 N_noxref_1_M1004_b N_A_27_115#_c_268_n 0.00873941f $X=-0.045 $Y=0
+ $X2=1.765 $Y2=1.845
cc_46 N_noxref_1_M1004_b N_A_27_115#_c_269_n 0.00735657f $X=-0.045 $Y=0
+ $X2=1.765 $Y2=2.885
cc_47 N_noxref_1_M1004_b N_A_27_115#_c_270_n 0.00873941f $X=-0.045 $Y=0
+ $X2=2.195 $Y2=1.845
cc_48 N_noxref_1_M1004_b N_A_27_115#_c_271_n 0.00735657f $X=-0.045 $Y=0
+ $X2=2.195 $Y2=2.885
cc_49 N_noxref_1_M1004_b N_A_27_115#_c_272_n 0.00873941f $X=-0.045 $Y=0
+ $X2=2.625 $Y2=1.845
cc_50 N_noxref_1_M1004_b N_A_27_115#_c_273_n 0.00735657f $X=-0.045 $Y=0
+ $X2=2.625 $Y2=2.885
cc_51 N_noxref_1_M1004_b N_A_27_115#_c_274_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.845
cc_52 N_noxref_1_M1004_b N_A_27_115#_c_275_n 0.00151234f $X=-0.045 $Y=0
+ $X2=3.055 $Y2=2.885
cc_53 N_noxref_1_M1004_b N_A_27_115#_c_276_n 0.0148636f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_54 N_noxref_1_c_2_p N_A_27_115#_c_276_n 0.00736239f $X=0.965 $Y=0.152
+ $X2=0.26 $Y2=0.825
cc_55 N_noxref_1_M1004_b N_A_27_115#_c_278_n 0.00626966f $X=-0.045 $Y=0
+ $X2=0.575 $Y2=3.545
cc_56 N_noxref_1_M1004_b N_A_27_115#_c_279_n 0.0164401f $X=-0.045 $Y=0 $X2=0.66
+ $Y2=1.935
cc_57 N_noxref_1_M1004_b N_A_27_115#_c_280_n 0.0251886f $X=-0.045 $Y=0 $X2=1.395
+ $Y2=1.935
cc_58 N_noxref_1_c_7_p N_A_27_115#_c_280_n 0.00704977f $X=1.05 $Y=0.825
+ $X2=1.395 $Y2=1.935
cc_59 N_noxref_1_M1004_b N_A_27_115#_c_282_n 0.0264756f $X=-0.045 $Y=0 $X2=1.395
+ $Y2=1.845
cc_60 N_noxref_1_M1004_b N_Y_c_423_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55
+ $Y2=1.595
cc_61 N_noxref_1_c_7_p N_Y_c_423_n 0.00127231f $X=1.05 $Y=0.825 $X2=1.55
+ $Y2=1.595
cc_62 N_noxref_1_c_20_p N_Y_c_423_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=1.55
+ $Y2=1.595
cc_63 N_noxref_1_M1004_b N_Y_c_426_n 0.00675046f $X=-0.045 $Y=0 $X2=1.55
+ $Y2=2.475
cc_64 N_noxref_1_M1004_b Y 0.030773f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_65 N_noxref_1_M1006_s N_Y_c_428_n 0.0127884f $X=1.84 $Y=0.575 $X2=2.265
+ $Y2=1.48
cc_66 N_noxref_1_c_20_p N_Y_c_428_n 0.0142303f $X=1.98 $Y=0.825 $X2=2.265
+ $Y2=1.48
cc_67 N_noxref_1_M1004_b N_Y_c_430_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.59
cc_68 N_noxref_1_M1004_b N_Y_c_431_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41
+ $Y2=2.475
cc_69 N_noxref_1_M1010_s N_Y_c_432_n 0.0127884f $X=2.7 $Y=0.575 $X2=3.125
+ $Y2=1.48
cc_70 N_noxref_1_c_31_p N_Y_c_432_n 0.0142303f $X=2.84 $Y=0.825 $X2=3.125
+ $Y2=1.48
cc_71 N_noxref_1_M1004_b N_Y_c_434_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555
+ $Y2=1.48
cc_72 N_noxref_1_c_20_p N_Y_c_434_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=2.555
+ $Y2=1.48
cc_73 N_noxref_1_c_31_p N_Y_c_434_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=2.555
+ $Y2=1.48
cc_74 N_noxref_1_M1004_b N_Y_c_437_n 0.0144211f $X=-0.045 $Y=0 $X2=3.125
+ $Y2=2.59
cc_75 N_noxref_1_M1004_b N_Y_c_438_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555
+ $Y2=2.59
cc_76 N_noxref_1_M1004_b N_Y_c_439_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27
+ $Y2=1.595
cc_77 N_noxref_1_c_31_p N_Y_c_439_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=3.27
+ $Y2=1.595
cc_78 N_noxref_1_c_43_p N_Y_c_439_n 0.00134236f $X=3.7 $Y=0.825 $X2=3.27
+ $Y2=1.595
cc_79 N_noxref_1_M1004_b N_Y_c_442_n 0.0485933f $X=-0.045 $Y=0 $X2=3.27
+ $Y2=2.475
cc_80 N_noxref_1_M1004_b N_Y_c_443_n 0.0110121f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_81 N_noxref_1_M1004_b N_Y_c_444_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.59
cc_82 N_noxref_1_M1004_b N_Y_c_445_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.59
cc_83 N_noxref_1_M1004_b N_Y_c_446_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55
+ $Y2=0.825
cc_84 N_noxref_1_c_7_p N_Y_c_446_n 0.0187614f $X=1.05 $Y=0.825 $X2=1.55
+ $Y2=0.825
cc_85 N_noxref_1_c_14_p N_Y_c_446_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55
+ $Y2=0.825
cc_86 N_noxref_1_c_20_p N_Y_c_446_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=1.55
+ $Y2=0.825
cc_87 N_noxref_1_M1004_b N_Y_c_450_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41
+ $Y2=0.825
cc_88 N_noxref_1_c_20_p N_Y_c_450_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=2.41
+ $Y2=0.825
cc_89 N_noxref_1_c_26_p N_Y_c_450_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41
+ $Y2=0.825
cc_90 N_noxref_1_c_31_p N_Y_c_450_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=2.41
+ $Y2=0.825
cc_91 N_noxref_1_M1004_b N_Y_c_454_n 0.00155118f $X=-0.045 $Y=0 $X2=3.27
+ $Y2=0.825
cc_92 N_noxref_1_c_31_p N_Y_c_454_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=3.27
+ $Y2=0.825
cc_93 N_noxref_1_c_37_p N_Y_c_454_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27
+ $Y2=0.825
cc_94 N_noxref_1_M1004_b GND 0.271923f $X=-0.045 $Y=0 $X2=0.34 $Y2=0.22
cc_95 N_noxref_1_c_2_p GND 0.0679129f $X=0.965 $Y=0.152 $X2=0.34 $Y2=0.22
cc_96 N_noxref_1_c_14_p GND 0.0478817f $X=1.895 $Y=0.152 $X2=0.34 $Y2=0.22
cc_97 N_noxref_1_c_26_p GND 0.0435303f $X=2.755 $Y=0.152 $X2=0.34 $Y2=0.22
cc_98 N_noxref_1_c_37_p GND 0.0898764f $X=3.615 $Y=0.152 $X2=0.34 $Y2=0.22
cc_99 N_noxref_1_c_99_p GND 0.0189324f $X=1.98 $Y=0.152 $X2=0.34 $Y2=0.22
cc_100 N_noxref_1_c_100_p GND 0.0189324f $X=2.84 $Y=0.152 $X2=0.34 $Y2=0.22
cc_101 N_noxref_2_M1005_b N_A_M1005_g 0.0189715f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_102 N_noxref_2_c_102_p N_A_M1005_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475
+ $Y2=4.585
cc_103 N_noxref_2_c_103_p N_A_M1005_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_104 N_noxref_2_M1005_s A 0.00790556f $X=0.135 $Y=3.085 $X2=0.24 $Y2=3.33
cc_105 N_noxref_2_M1005_b A 0.0115315f $X=-0.045 $Y=2.905 $X2=0.24 $Y2=3.33
cc_106 N_noxref_2_c_102_p A 0.00459217f $X=0.26 $Y=4.135 $X2=0.24 $Y2=3.33
cc_107 N_noxref_2_M1005_s N_A_c_170_n 0.0150633f $X=0.135 $Y=3.085 $X2=0.235
+ $Y2=2.765
cc_108 N_noxref_2_M1005_b N_A_c_170_n 0.00613107f $X=-0.045 $Y=2.905 $X2=0.235
+ $Y2=2.765
cc_109 N_noxref_2_c_102_p N_A_c_170_n 0.00337102f $X=0.26 $Y=4.135 $X2=0.235
+ $Y2=2.765
cc_110 N_noxref_2_M1005_b N_A_c_171_n 0.0124943f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.765
cc_111 N_noxref_2_M1005_b N_B_M1000_g 0.0187479f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_112 N_noxref_2_c_103_p N_B_M1000_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905
+ $Y2=4.585
cc_113 N_noxref_2_c_113_p N_B_M1000_g 0.00354579f $X=1.12 $Y=3.795 $X2=0.905
+ $Y2=4.585
cc_114 N_noxref_2_M1005_b B 0.00872506f $X=-0.045 $Y=2.905 $X2=0.92 $Y2=2.96
cc_115 N_noxref_2_c_113_p B 9.65504e-19 $X=1.12 $Y=3.795 $X2=0.92 $Y2=2.96
cc_116 N_noxref_2_M1005_b N_B_c_202_n 0.00130234f $X=-0.045 $Y=2.905 $X2=0.915
+ $Y2=2.425
cc_117 N_noxref_2_M1005_b N_A_27_115#_c_283_n 0.0171069f $X=-0.045 $Y=2.905
+ $X2=1.335 $Y2=2.96
cc_118 N_noxref_2_c_113_p N_A_27_115#_c_283_n 0.00354579f $X=1.12 $Y=3.795
+ $X2=1.335 $Y2=2.96
cc_119 N_noxref_2_c_119_p N_A_27_115#_c_283_n 0.00606474f $X=1.895 $Y=6.507
+ $X2=1.335 $Y2=2.96
cc_120 N_noxref_2_M1005_b N_A_27_115#_c_239_n 0.00448664f $X=-0.045 $Y=2.905
+ $X2=1.69 $Y2=2.885
cc_121 N_noxref_2_M1005_b N_A_27_115#_c_287_n 0.017006f $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.96
cc_122 N_noxref_2_c_113_p N_A_27_115#_c_287_n 3.67508e-19 $X=1.12 $Y=3.795
+ $X2=1.765 $Y2=2.96
cc_123 N_noxref_2_c_119_p N_A_27_115#_c_287_n 0.00610567f $X=1.895 $Y=6.507
+ $X2=1.765 $Y2=2.96
cc_124 N_noxref_2_c_124_p N_A_27_115#_c_287_n 0.00373985f $X=1.98 $Y=3.455
+ $X2=1.765 $Y2=2.96
cc_125 N_noxref_2_M1005_b N_A_27_115#_c_246_n 0.00396043f $X=-0.045 $Y=2.905
+ $X2=2.12 $Y2=2.885
cc_126 N_noxref_2_c_124_p N_A_27_115#_c_246_n 0.00379272f $X=1.98 $Y=3.455
+ $X2=2.12 $Y2=2.885
cc_127 N_noxref_2_M1005_b N_A_27_115#_c_293_n 0.0166898f $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.96
cc_128 N_noxref_2_c_124_p N_A_27_115#_c_293_n 0.00354579f $X=1.98 $Y=3.455
+ $X2=2.195 $Y2=2.96
cc_129 N_noxref_2_c_129_p N_A_27_115#_c_293_n 0.00606474f $X=2.755 $Y=6.507
+ $X2=2.195 $Y2=2.96
cc_130 N_noxref_2_M1005_b N_A_27_115#_c_251_n 0.00448664f $X=-0.045 $Y=2.905
+ $X2=2.55 $Y2=2.885
cc_131 N_noxref_2_M1005_b N_A_27_115#_c_297_n 0.0166898f $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=2.96
cc_132 N_noxref_2_c_129_p N_A_27_115#_c_297_n 0.00606474f $X=2.755 $Y=6.507
+ $X2=2.625 $Y2=2.96
cc_133 N_noxref_2_c_133_p N_A_27_115#_c_297_n 0.00354579f $X=2.84 $Y=3.455
+ $X2=2.625 $Y2=2.96
cc_134 N_noxref_2_M1005_b N_A_27_115#_c_257_n 0.00396043f $X=-0.045 $Y=2.905
+ $X2=2.98 $Y2=2.885
cc_135 N_noxref_2_c_133_p N_A_27_115#_c_257_n 0.00379272f $X=2.84 $Y=3.455
+ $X2=2.98 $Y2=2.885
cc_136 N_noxref_2_M1005_b N_A_27_115#_c_302_n 0.0166898f $X=-0.045 $Y=2.905
+ $X2=3.055 $Y2=2.96
cc_137 N_noxref_2_c_133_p N_A_27_115#_c_302_n 0.00354579f $X=2.84 $Y=3.455
+ $X2=3.055 $Y2=2.96
cc_138 N_noxref_2_c_138_p N_A_27_115#_c_302_n 0.00606474f $X=3.615 $Y=6.507
+ $X2=3.055 $Y2=2.96
cc_139 N_noxref_2_M1005_b N_A_27_115#_c_263_n 0.00840215f $X=-0.045 $Y=2.905
+ $X2=3.41 $Y2=2.885
cc_140 N_noxref_2_M1005_b N_A_27_115#_c_306_n 0.0209036f $X=-0.045 $Y=2.905
+ $X2=3.485 $Y2=2.96
cc_141 N_noxref_2_c_138_p N_A_27_115#_c_306_n 0.00606474f $X=3.615 $Y=6.507
+ $X2=3.485 $Y2=2.96
cc_142 N_noxref_2_c_142_p N_A_27_115#_c_306_n 0.00713292f $X=3.7 $Y=3.455
+ $X2=3.485 $Y2=2.96
cc_143 N_noxref_2_M1005_b N_A_27_115#_c_267_n 0.00196792f $X=-0.045 $Y=2.905
+ $X2=1.335 $Y2=2.885
cc_144 N_noxref_2_M1005_b N_A_27_115#_c_269_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.885
cc_145 N_noxref_2_M1005_b N_A_27_115#_c_271_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.885
cc_146 N_noxref_2_M1005_b N_A_27_115#_c_273_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=2.885
cc_147 N_noxref_2_M1005_b N_A_27_115#_c_275_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=3.055 $Y2=2.885
cc_148 N_noxref_2_M1005_b N_A_27_115#_c_278_n 8.35397e-19 $X=-0.045 $Y=2.905
+ $X2=0.575 $Y2=3.545
cc_149 N_noxref_2_M1005_b N_A_27_115#_c_315_n 0.00155118f $X=-0.045 $Y=2.905
+ $X2=0.69 $Y2=3.795
cc_150 N_noxref_2_c_103_p N_A_27_115#_c_315_n 0.0075556f $X=1.035 $Y=6.507
+ $X2=0.69 $Y2=3.795
cc_151 N_noxref_2_c_124_p N_Y_c_430_n 0.00634153f $X=1.98 $Y=3.455 $X2=2.265
+ $Y2=2.59
cc_152 N_noxref_2_c_133_p N_Y_c_437_n 0.00634153f $X=2.84 $Y=3.455 $X2=3.125
+ $Y2=2.59
cc_153 N_noxref_2_M1005_b N_Y_c_443_n 0.00347838f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=2.59
cc_154 N_noxref_2_c_119_p N_Y_c_443_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55
+ $Y2=2.59
cc_155 N_noxref_2_M1005_b N_Y_c_444_n 0.00380347f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.59
cc_156 N_noxref_2_c_129_p N_Y_c_444_n 0.00734006f $X=2.755 $Y=6.507 $X2=2.41
+ $Y2=2.59
cc_157 N_noxref_2_M1005_b N_Y_c_445_n 0.00380347f $X=-0.045 $Y=2.905 $X2=3.27
+ $Y2=2.59
cc_158 N_noxref_2_c_138_p N_Y_c_445_n 0.00745425f $X=3.615 $Y=6.507 $X2=3.27
+ $Y2=2.59
cc_159 N_noxref_2_M1005_b VDD 0.278838f $X=-0.045 $Y=2.905 $X2=0.34 $Y2=6.44
cc_160 N_noxref_2_c_160_p VDD 0.0381711f $X=0.26 $Y=6.355 $X2=0.34 $Y2=6.44
cc_161 N_noxref_2_c_103_p VDD 0.0429496f $X=1.035 $Y=6.507 $X2=0.34 $Y2=6.44
cc_162 N_noxref_2_c_119_p VDD 0.0434027f $X=1.895 $Y=6.507 $X2=0.34 $Y2=6.44
cc_163 N_noxref_2_c_129_p VDD 0.0435303f $X=2.755 $Y=6.507 $X2=0.34 $Y2=6.44
cc_164 N_noxref_2_c_138_p VDD 0.0898764f $X=3.615 $Y=6.507 $X2=0.34 $Y2=6.44
cc_165 N_noxref_2_c_165_p VDD 0.0189324f $X=1.12 $Y=6.507 $X2=0.34 $Y2=6.44
cc_166 N_noxref_2_c_166_p VDD 0.0189324f $X=1.98 $Y=6.507 $X2=0.34 $Y2=6.44
cc_167 N_noxref_2_c_167_p VDD 0.0189324f $X=2.84 $Y=6.507 $X2=0.34 $Y2=6.44
cc_168 N_A_M1004_g N_B_M1002_g 0.129389f $X=0.475 $Y=1.075 $X2=0.835 $Y2=1.075
cc_169 N_A_M1004_g N_B_M1000_g 0.0497852f $X=0.475 $Y=1.075 $X2=0.905 $Y2=4.585
cc_170 N_A_M1004_g N_B_c_202_n 8.69605e-19 $X=0.475 $Y=1.075 $X2=0.915 $Y2=2.425
cc_171 N_A_M1004_g N_A_27_115#_c_276_n 0.0158254f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_172 N_A_M1004_g N_A_27_115#_c_278_n 0.0278506f $X=0.475 $Y=1.075 $X2=0.575
+ $Y2=3.545
cc_173 N_A_M1005_g N_A_27_115#_c_278_n 0.0152191f $X=0.475 $Y=4.585 $X2=0.575
+ $Y2=3.545
cc_174 A N_A_27_115#_c_278_n 0.00781918f $X=0.24 $Y=3.33 $X2=0.575 $Y2=3.545
cc_175 N_A_c_170_n N_A_27_115#_c_278_n 0.053763f $X=0.235 $Y=2.765 $X2=0.575
+ $Y2=3.545
cc_176 N_A_c_171_n N_A_27_115#_c_278_n 0.00844699f $X=0.475 $Y=2.765 $X2=0.575
+ $Y2=3.545
cc_177 N_A_M1004_g N_A_27_115#_c_279_n 0.0178909f $X=0.475 $Y=1.075 $X2=0.66
+ $Y2=1.935
cc_178 N_A_c_170_n N_A_27_115#_c_279_n 0.00451097f $X=0.235 $Y=2.765 $X2=0.66
+ $Y2=1.935
cc_179 N_A_c_171_n N_A_27_115#_c_279_n 0.00272689f $X=0.475 $Y=2.765 $X2=0.66
+ $Y2=1.935
cc_180 N_A_M1005_g N_A_27_115#_c_326_n 0.0109054f $X=0.475 $Y=4.585 $X2=0.69
+ $Y2=3.63
cc_181 N_A_M1004_g GND 0.00468827f $X=0.475 $Y=1.075 $X2=0.34 $Y2=0.22
cc_182 N_A_M1005_g VDD 0.00468827f $X=0.475 $Y=4.585 $X2=0.34 $Y2=6.44
cc_183 N_B_M1002_g N_A_27_115#_M1001_g 0.0468623f $X=0.835 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_184 N_B_M1000_g N_A_27_115#_c_238_n 0.0492452f $X=0.905 $Y=4.585 $X2=1.335
+ $Y2=2.81
cc_185 N_B_c_202_n N_A_27_115#_c_238_n 0.00498982f $X=0.915 $Y=2.425 $X2=1.335
+ $Y2=2.81
cc_186 N_B_c_203_n N_A_27_115#_c_238_n 0.0207593f $X=0.915 $Y=2.425 $X2=1.335
+ $Y2=2.81
cc_187 B N_A_27_115#_c_267_n 0.00380362f $X=0.92 $Y=2.96 $X2=1.335 $Y2=2.885
cc_188 N_B_M1002_g N_A_27_115#_c_278_n 0.00719886f $X=0.835 $Y=1.075 $X2=0.575
+ $Y2=3.545
cc_189 N_B_M1000_g N_A_27_115#_c_278_n 0.01267f $X=0.905 $Y=4.585 $X2=0.575
+ $Y2=3.545
cc_190 B N_A_27_115#_c_278_n 0.00871807f $X=0.92 $Y=2.96 $X2=0.575 $Y2=3.545
cc_191 N_B_c_202_n N_A_27_115#_c_278_n 0.0541394f $X=0.915 $Y=2.425 $X2=0.575
+ $Y2=3.545
cc_192 N_B_M1002_g N_A_27_115#_c_280_n 0.0171085f $X=0.835 $Y=1.075 $X2=1.395
+ $Y2=1.935
cc_193 N_B_c_202_n N_A_27_115#_c_280_n 0.0100447f $X=0.915 $Y=2.425 $X2=1.395
+ $Y2=1.935
cc_194 N_B_c_203_n N_A_27_115#_c_280_n 0.00235847f $X=0.915 $Y=2.425 $X2=1.395
+ $Y2=1.935
cc_195 B N_A_27_115#_c_326_n 0.00385574f $X=0.92 $Y=2.96 $X2=0.69 $Y2=3.63
cc_196 N_B_M1002_g N_Y_c_423_n 8.18972e-19 $X=0.835 $Y=1.075 $X2=1.55 $Y2=1.595
cc_197 N_B_c_202_n N_Y_c_426_n 0.00573285f $X=0.915 $Y=2.425 $X2=1.55 $Y2=2.475
cc_198 N_B_c_203_n N_Y_c_426_n 5.80618e-19 $X=0.915 $Y=2.425 $X2=1.55 $Y2=2.475
cc_199 N_B_M1002_g Y 6.5988e-19 $X=0.835 $Y=1.075 $X2=1.555 $Y2=2.22
cc_200 N_B_c_202_n Y 0.00671947f $X=0.915 $Y=2.425 $X2=1.555 $Y2=2.22
cc_201 B N_Y_c_443_n 0.00632423f $X=0.92 $Y=2.96 $X2=1.55 $Y2=2.59
cc_202 N_B_c_202_n N_Y_c_443_n 0.0138653f $X=0.915 $Y=2.425 $X2=1.55 $Y2=2.59
cc_203 N_B_M1002_g GND 0.00468827f $X=0.835 $Y=1.075 $X2=0.34 $Y2=0.22
cc_204 N_B_M1000_g VDD 0.00468827f $X=0.905 $Y=4.585 $X2=0.34 $Y2=6.44
cc_205 N_A_27_115#_M1001_g N_Y_c_423_n 0.00554705f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_206 N_A_27_115#_M1006_g N_Y_c_423_n 0.00259902f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_207 N_A_27_115#_c_280_n N_Y_c_423_n 0.00238892f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=1.595
cc_208 N_A_27_115#_c_238_n N_Y_c_426_n 0.00638728f $X=1.335 $Y=2.81 $X2=1.55
+ $Y2=2.475
cc_209 N_A_27_115#_c_239_n N_Y_c_426_n 0.00186325f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.475
cc_210 N_A_27_115#_c_240_n N_Y_c_426_n 0.00140336f $X=1.69 $Y=1.845 $X2=1.55
+ $Y2=2.475
cc_211 N_A_27_115#_c_280_n N_Y_c_426_n 0.00194461f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=2.475
cc_212 N_A_27_115#_c_282_n N_Y_c_426_n 0.00144278f $X=1.395 $Y=1.845 $X2=1.55
+ $Y2=2.475
cc_213 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_214 N_A_27_115#_c_238_n Y 0.00874077f $X=1.335 $Y=2.81 $X2=1.555 $Y2=2.22
cc_215 N_A_27_115#_c_240_n Y 0.00840707f $X=1.69 $Y=1.845 $X2=1.555 $Y2=2.22
cc_216 N_A_27_115#_M1006_g Y 0.00251111f $X=1.765 $Y=1.075 $X2=1.555 $Y2=2.22
cc_217 N_A_27_115#_c_280_n Y 0.0132141f $X=1.395 $Y=1.935 $X2=1.555 $Y2=2.22
cc_218 N_A_27_115#_c_282_n Y 0.00487273f $X=1.395 $Y=1.845 $X2=1.555 $Y2=2.22
cc_219 N_A_27_115#_M1006_g N_Y_c_428_n 0.0130095f $X=1.765 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_220 N_A_27_115#_c_244_n N_Y_c_428_n 0.00213861f $X=2.12 $Y=1.845 $X2=2.265
+ $Y2=1.48
cc_221 N_A_27_115#_M1008_g N_Y_c_428_n 0.0130095f $X=2.195 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_222 N_A_27_115#_c_268_n N_Y_c_430_n 0.0121767f $X=1.765 $Y=1.845 $X2=2.265
+ $Y2=2.59
cc_223 N_A_27_115#_c_269_n N_Y_c_430_n 0.0158479f $X=1.765 $Y=2.885 $X2=2.265
+ $Y2=2.59
cc_224 N_A_27_115#_M1008_g N_Y_c_431_n 0.00251111f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_225 N_A_27_115#_c_250_n N_Y_c_431_n 0.0177725f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.475
cc_226 N_A_27_115#_M1010_g N_Y_c_431_n 0.00251111f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_227 N_A_27_115#_c_261_n N_Y_c_431_n 0.00843025f $X=3.055 $Y=2.81 $X2=2.41
+ $Y2=2.475
cc_228 N_A_27_115#_M1010_g N_Y_c_432_n 0.0130095f $X=2.625 $Y=1.075 $X2=3.125
+ $Y2=1.48
cc_229 N_A_27_115#_c_255_n N_Y_c_432_n 0.00213861f $X=2.98 $Y=1.845 $X2=3.125
+ $Y2=1.48
cc_230 N_A_27_115#_M1012_g N_Y_c_432_n 0.0136594f $X=3.055 $Y=1.075 $X2=3.125
+ $Y2=1.48
cc_231 N_A_27_115#_M1008_g N_Y_c_434_n 0.00259902f $X=2.195 $Y=1.075 $X2=2.555
+ $Y2=1.48
cc_232 N_A_27_115#_M1010_g N_Y_c_434_n 0.00259902f $X=2.625 $Y=1.075 $X2=2.555
+ $Y2=1.48
cc_233 N_A_27_115#_c_261_n N_Y_c_437_n 0.0155956f $X=3.055 $Y=2.81 $X2=3.125
+ $Y2=2.59
cc_234 N_A_27_115#_c_272_n N_Y_c_437_n 0.00894336f $X=2.625 $Y=1.845 $X2=3.125
+ $Y2=2.59
cc_235 N_A_27_115#_c_273_n N_Y_c_437_n 0.00903839f $X=2.625 $Y=2.885 $X2=3.125
+ $Y2=2.59
cc_236 N_A_27_115#_c_250_n N_Y_c_438_n 0.00140336f $X=2.55 $Y=1.845 $X2=2.555
+ $Y2=2.59
cc_237 N_A_27_115#_c_261_n N_Y_c_438_n 0.0012308f $X=3.055 $Y=2.81 $X2=2.555
+ $Y2=2.59
cc_238 N_A_27_115#_c_270_n N_Y_c_438_n 0.00140336f $X=2.195 $Y=1.845 $X2=2.555
+ $Y2=2.59
cc_239 N_A_27_115#_c_271_n N_Y_c_438_n 0.00372651f $X=2.195 $Y=2.885 $X2=2.555
+ $Y2=2.59
cc_240 N_A_27_115#_M1012_g N_Y_c_439_n 0.00262362f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_241 N_A_27_115#_M1014_g N_Y_c_439_n 0.00939545f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_242 N_A_27_115#_M1012_g N_Y_c_442_n 0.00251111f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=2.475
cc_243 N_A_27_115#_c_261_n N_Y_c_442_n 0.0163934f $X=3.055 $Y=2.81 $X2=3.27
+ $Y2=2.475
cc_244 N_A_27_115#_c_262_n N_Y_c_442_n 0.0196907f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=2.475
cc_245 N_A_27_115#_c_263_n N_Y_c_442_n 0.00357274f $X=3.41 $Y=2.885 $X2=3.27
+ $Y2=2.475
cc_246 N_A_27_115#_M1014_g N_Y_c_442_n 0.00251111f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=2.475
cc_247 N_A_27_115#_c_238_n N_Y_c_443_n 0.00711959f $X=1.335 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_248 N_A_27_115#_c_283_n N_Y_c_443_n 0.00282264f $X=1.335 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_249 N_A_27_115#_c_239_n N_Y_c_443_n 0.0163883f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.59
cc_250 N_A_27_115#_c_240_n N_Y_c_443_n 0.00122399f $X=1.69 $Y=1.845 $X2=1.55
+ $Y2=2.59
cc_251 N_A_27_115#_c_287_n N_Y_c_443_n 0.00392729f $X=1.765 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_252 N_A_27_115#_c_280_n N_Y_c_443_n 0.00202105f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_253 N_A_27_115#_c_282_n N_Y_c_443_n 6.59752e-19 $X=1.395 $Y=1.845 $X2=1.55
+ $Y2=2.59
cc_254 N_A_27_115#_c_293_n N_Y_c_444_n 0.00392729f $X=2.195 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_255 N_A_27_115#_c_250_n N_Y_c_444_n 0.00250559f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.59
cc_256 N_A_27_115#_c_251_n N_Y_c_444_n 0.021445f $X=2.55 $Y=2.885 $X2=2.41
+ $Y2=2.59
cc_257 N_A_27_115#_c_297_n N_Y_c_444_n 0.00392729f $X=2.625 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_258 N_A_27_115#_c_261_n N_Y_c_444_n 0.00361281f $X=3.055 $Y=2.81 $X2=2.41
+ $Y2=2.59
cc_259 N_A_27_115#_c_261_n N_Y_c_445_n 0.00721971f $X=3.055 $Y=2.81 $X2=3.27
+ $Y2=2.59
cc_260 N_A_27_115#_c_302_n N_Y_c_445_n 0.00392729f $X=3.055 $Y=2.96 $X2=3.27
+ $Y2=2.59
cc_261 N_A_27_115#_c_262_n N_Y_c_445_n 0.00250559f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=2.59
cc_262 N_A_27_115#_c_263_n N_Y_c_445_n 0.0206674f $X=3.41 $Y=2.885 $X2=3.27
+ $Y2=2.59
cc_263 N_A_27_115#_c_306_n N_Y_c_445_n 0.00392729f $X=3.485 $Y=2.96 $X2=3.27
+ $Y2=2.59
cc_264 N_A_27_115#_M1001_g N_Y_c_446_n 0.00233629f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_265 N_A_27_115#_M1006_g N_Y_c_446_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_266 N_A_27_115#_c_280_n N_Y_c_446_n 0.00364905f $X=1.395 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_267 N_A_27_115#_c_282_n N_Y_c_446_n 0.00208849f $X=1.395 $Y=1.845 $X2=1.55
+ $Y2=0.825
cc_268 N_A_27_115#_M1008_g N_Y_c_450_n 0.00231637f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_269 N_A_27_115#_c_250_n N_Y_c_450_n 0.00280419f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=0.825
cc_270 N_A_27_115#_M1010_g N_Y_c_450_n 0.00231637f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_271 N_A_27_115#_M1012_g N_Y_c_454_n 0.00231637f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=0.825
cc_272 N_A_27_115#_c_262_n N_Y_c_454_n 0.00280419f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=0.825
cc_273 N_A_27_115#_M1014_g N_Y_c_454_n 0.00231637f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=0.825
cc_274 N_A_27_115#_M1001_g GND 0.00468827f $X=1.335 $Y=1.075 $X2=0.34 $Y2=0.22
cc_275 N_A_27_115#_M1006_g GND 0.00468827f $X=1.765 $Y=1.075 $X2=0.34 $Y2=0.22
cc_276 N_A_27_115#_M1008_g GND 0.00468827f $X=2.195 $Y=1.075 $X2=0.34 $Y2=0.22
cc_277 N_A_27_115#_M1010_g GND 0.00468827f $X=2.625 $Y=1.075 $X2=0.34 $Y2=0.22
cc_278 N_A_27_115#_M1012_g GND 0.00468827f $X=3.055 $Y=1.075 $X2=0.34 $Y2=0.22
cc_279 N_A_27_115#_M1014_g GND 0.00468827f $X=3.485 $Y=1.075 $X2=0.34 $Y2=0.22
cc_280 N_A_27_115#_c_276_n GND 0.00476261f $X=0.26 $Y=0.825 $X2=0.34 $Y2=0.22
cc_281 N_A_27_115#_c_283_n VDD 0.00468827f $X=1.335 $Y=2.96 $X2=0.34 $Y2=6.44
cc_282 N_A_27_115#_c_287_n VDD 0.00470215f $X=1.765 $Y=2.96 $X2=0.34 $Y2=6.44
cc_283 N_A_27_115#_c_293_n VDD 0.00468827f $X=2.195 $Y=2.96 $X2=0.34 $Y2=6.44
cc_284 N_A_27_115#_c_297_n VDD 0.00468827f $X=2.625 $Y=2.96 $X2=0.34 $Y2=6.44
cc_285 N_A_27_115#_c_302_n VDD 0.00468827f $X=3.055 $Y=2.96 $X2=0.34 $Y2=6.44
cc_286 N_A_27_115#_c_306_n VDD 0.00468827f $X=3.485 $Y=2.96 $X2=0.34 $Y2=6.44
cc_287 N_A_27_115#_c_315_n VDD 0.00475776f $X=0.69 $Y=3.795 $X2=0.34 $Y2=6.44
cc_288 N_Y_c_446_n GND 0.00475776f $X=1.55 $Y=0.825 $X2=0.34 $Y2=0.22
cc_289 N_Y_c_450_n GND 0.00475776f $X=2.41 $Y=0.825 $X2=0.34 $Y2=0.22
cc_290 N_Y_c_454_n GND 0.00475776f $X=3.27 $Y=0.825 $X2=0.34 $Y2=0.22
cc_291 N_Y_c_443_n VDD 0.00475776f $X=1.55 $Y=2.59 $X2=0.34 $Y2=6.44
cc_292 N_Y_c_444_n VDD 0.00475776f $X=2.41 $Y=2.59 $X2=0.34 $Y2=6.44
cc_293 N_Y_c_445_n VDD 0.00475776f $X=3.27 $Y=2.59 $X2=0.34 $Y2=6.44
