* File: sky130_osu_sc_12T_ls__dffs_1.pex.spice
* Created: Fri Nov 12 15:36:23 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%GND 1 2 3 4 5 6 97 99 107 109 113 115
+ 125 127 137 139 149 151 158 180 182
c216 137 0 3.34232e-19 $X=5.14 $Y=0.755
c217 113 0 3.14854e-19 $X=1.64 $Y=0.755
c218 97 0 1.27355e-19 $X=-0.055 $Y=0
r219 180 182 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=7.815 $Y2=0.152
r220 156 158 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.74
r221 152 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=0.152
+ $X2=6.88 $Y2=0.152
r222 147 172 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.152
r223 147 149 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.74
r224 139 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=0.152
+ $X2=6.88 $Y2=0.152
r225 135 137 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.14 $Y=0.305
+ $X2=5.14 $Y2=0.755
r226 128 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.152
+ $X2=3.39 $Y2=0.152
r227 123 168 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.152
r228 123 125 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.74
r229 115 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.152
+ $X2=3.39 $Y2=0.152
r230 111 113 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.64 $Y=0.305
+ $X2=1.64 $Y2=0.755
r231 109 110 15.8697 $w=3.03e-07 $l=4.2e-07 $layer=LI1_cond $X=1.555 $Y=0.152
+ $X2=1.135 $Y2=0.152
r232 105 107 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r233 97 182 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=0.19
+ $X2=7.815 $Y2=0.19
r234 97 180 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r235 97 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r236 97 151 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r237 97 135 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.14 $Y2=0.305
r238 97 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.055 $Y2=0.152
r239 97 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.225 $Y2=0.152
r240 97 111 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.64 $Y2=0.305
r241 97 109 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.555 $Y2=0.152
r242 97 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.725 $Y2=0.152
r243 97 105 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r244 97 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r245 97 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r246 97 151 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r247 97 152 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.965 $Y2=0.152
r248 97 139 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.795 $Y2=0.152
r249 97 140 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=5.225 $Y2=0.152
r250 97 127 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=5.055 $Y2=0.152
r251 97 128 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.475 $Y2=0.152
r252 97 115 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=3.305 $Y2=0.152
r253 97 116 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=1.725 $Y2=0.152
r254 97 99 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=0.335 $Y=0.152
+ $X2=0.965 $Y2=0.152
r255 6 158 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.74
r256 5 149 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.575 $X2=6.88 $Y2=0.74
r257 4 137 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5 $Y=0.575
+ $X2=5.14 $Y2=0.755
r258 3 125 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.575 $X2=3.39 $Y2=0.74
r259 2 113 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.575 $X2=1.64 $Y2=0.755
r260 1 107 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%VDD 1 2 3 4 5 6 7 8 81 85 87 93 99 101
+ 109 111 119 121 127 129 135 137 143 159 162 166
c113 143 0 1.98165e-19 $X=7.9 $Y=3.265
r114 162 166 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=4.287
+ $X2=7.815 $Y2=4.287
r115 159 166 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=4.25
+ $X2=7.815 $Y2=4.25
r116 148 162 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=4.25
+ $X2=0.335 $Y2=4.25
r117 141 159 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=4.287
r118 141 143 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=3.265
r119 138 157 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.035 $Y=4.287
+ $X2=6.95 $Y2=4.287
r120 138 140 3.7785 $w=3.03e-07 $l=1e-07 $layer=LI1_cond $X=7.035 $Y=4.287
+ $X2=7.135 $Y2=4.287
r121 137 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=4.287
+ $X2=7.9 $Y2=4.287
r122 137 140 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=4.287
+ $X2=7.135 $Y2=4.287
r123 133 157 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.95 $Y=4.135
+ $X2=6.95 $Y2=4.287
r124 133 135 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.95 $Y=4.135
+ $X2=6.95 $Y2=3.615
r125 130 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.09 $Y2=4.287
r126 130 132 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.455 $Y2=4.287
r127 129 157 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=4.287
+ $X2=6.95 $Y2=4.287
r128 129 132 15.4919 $w=3.03e-07 $l=4.1e-07 $layer=LI1_cond $X=6.865 $Y=4.287
+ $X2=6.455 $Y2=4.287
r129 125 156 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=4.287
r130 125 127 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=3.615
r131 122 155 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=4.287
+ $X2=5.14 $Y2=4.287
r132 122 124 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.225 $Y=4.287
+ $X2=5.775 $Y2=4.287
r133 121 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=6.09 $Y2=4.287
r134 121 124 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=5.775 $Y2=4.287
r135 117 155 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.14 $Y=4.135
+ $X2=5.14 $Y2=4.287
r136 117 119 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.14 $Y=4.135
+ $X2=5.14 $Y2=3.21
r137 114 116 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=4.287
+ $X2=4.415 $Y2=4.287
r138 112 153 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=4.287
+ $X2=3.39 $Y2=4.287
r139 112 114 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.475 $Y=4.287
+ $X2=3.735 $Y2=4.287
r140 111 155 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=4.287
+ $X2=5.14 $Y2=4.287
r141 111 116 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=5.055 $Y=4.287
+ $X2=4.415 $Y2=4.287
r142 107 153 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.39 $Y=4.135
+ $X2=3.39 $Y2=4.287
r143 107 109 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.39 $Y=4.135
+ $X2=3.39 $Y2=3.295
r144 104 106 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.375 $Y=4.287
+ $X2=3.055 $Y2=4.287
r145 102 152 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=4.287
+ $X2=1.64 $Y2=4.287
r146 102 104 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=1.725 $Y=4.287
+ $X2=2.375 $Y2=4.287
r147 101 153 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=4.287
+ $X2=3.39 $Y2=4.287
r148 101 106 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.305 $Y=4.287
+ $X2=3.055 $Y2=4.287
r149 97 152 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.64 $Y=4.135
+ $X2=1.64 $Y2=4.287
r150 97 99 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.64 $Y=4.135
+ $X2=1.64 $Y2=3.295
r151 96 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r152 95 152 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=4.287
+ $X2=1.64 $Y2=4.287
r153 95 96 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=1.555 $Y=4.287
+ $X2=1.205 $Y2=4.287
r154 91 150 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r155 91 93 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.615
r156 88 148 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r157 88 90 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.015 $Y2=4.287
r158 87 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r159 87 90 0.7557 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.015 $Y2=4.287
r160 83 148 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r161 83 85 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.615
r162 81 159 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=4.135 $X2=7.815 $Y2=4.22
r163 81 140 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=4.135 $X2=7.135 $Y2=4.22
r164 81 132 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=4.135 $X2=6.455 $Y2=4.22
r165 81 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=4.135 $X2=5.775 $Y2=4.22
r166 81 155 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=4.135 $X2=5.095 $Y2=4.22
r167 81 116 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=4.135 $X2=4.415 $Y2=4.22
r168 81 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=4.135 $X2=3.735 $Y2=4.22
r169 81 106 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=4.135 $X2=3.055 $Y2=4.22
r170 81 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=4.135 $X2=2.375 $Y2=4.22
r171 81 152 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=4.135 $X2=1.695 $Y2=4.22
r172 81 90 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=4.135 $X2=1.015 $Y2=4.22
r173 81 148 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=4.135 $X2=0.335 $Y2=4.22
r174 8 143 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=2.605 $X2=7.9 $Y2=3.265
r175 7 135 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=3.025 $X2=6.95 $Y2=3.615
r176 6 127 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=5.965
+ $Y=3.025 $X2=6.09 $Y2=3.615
r177 5 119 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=5
+ $Y=2.605 $X2=5.14 $Y2=3.21
r178 4 109 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=3.25
+ $Y=2.605 $X2=3.39 $Y2=3.295
r179 3 99 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=2.605 $X2=1.64 $Y2=3.295
r180 2 93 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=3.025 $X2=1.12 $Y2=3.615
r181 1 85 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.615
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%SN 3 7 9 11 14 17 21 25 31 35 36 37 39
c149 31 0 1.11496e-19 $X=6.94 $Y=1.165
c150 21 0 1.08672e-19 $X=6.735 $Y=1.232
c151 9 0 6.64688e-20 $X=6.665 $Y=1.04
r152 36 44 4.46514 $w=1.55e-07 $l=5.57237e-06 $layer=MET1_cond $X=1.405 $Y=0.985
+ $X2=6.94 $Y2=1.06
r153 36 37 1.23762 $w=1.4e-07 $l=1e-06 $layer=MET1_cond $X=1.405 $Y=0.985
+ $X2=0.405 $Y2=0.985
r154 35 39 0.0828968 $w=2.9e-07 $l=1.2e-07 $layer=MET1_cond $X=0.32 $Y=1.415
+ $X2=0.32 $Y2=1.535
r155 34 37 0.0706952 $w=1.4e-07 $l=1.14782e-07 $layer=MET1_cond $X=0.32 $Y=1.055
+ $X2=0.405 $Y2=0.985
r156 34 35 0.346638 $w=1.7e-07 $l=3.6e-07 $layer=MET1_cond $X=0.32 $Y=1.055
+ $X2=0.32 $Y2=1.415
r157 31 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.94 $Y=1.165
+ $X2=6.94 $Y2=1.165
r158 31 33 2.09542 $w=2.62e-07 $l=4.5e-08 $layer=LI1_cond $X=6.94 $Y=1.165
+ $X2=6.94 $Y2=1.21
r159 28 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=1.535
+ $X2=0.32 $Y2=1.535
r160 25 28 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.32 $Y=1.47
+ $X2=0.32 $Y2=1.535
r161 23 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.94
+ $Y=1.21 $X2=6.94 $Y2=1.21
r162 21 23 27.0712 $w=3.65e-07 $l=2.05e-07 $layer=POLY_cond $X=6.735 $Y=1.232
+ $X2=6.94 $Y2=1.232
r163 20 21 9.24384 $w=3.65e-07 $l=7e-08 $layer=POLY_cond $X=6.665 $Y=1.232
+ $X2=6.735 $Y2=1.232
r164 17 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.47 $X2=0.32 $Y2=1.47
r165 17 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.47
+ $X2=0.367 $Y2=1.635
r166 17 18 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.47
+ $X2=0.367 $Y2=1.305
r167 12 21 23.6381 $w=1.5e-07 $l=1.93e-07 $layer=POLY_cond $X=6.735 $Y=1.425
+ $X2=6.735 $Y2=1.232
r168 12 14 1035.79 $w=1.5e-07 $l=2.02e-06 $layer=POLY_cond $X=6.735 $Y=1.425
+ $X2=6.735 $Y2=3.445
r169 9 20 23.6381 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.665 $Y=1.04
+ $X2=6.665 $Y2=1.232
r170 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.665 $Y=1.04
+ $X2=6.665 $Y2=0.755
r171 7 19 928.106 $w=1.5e-07 $l=1.81e-06 $layer=POLY_cond $X=0.475 $Y=3.445
+ $X2=0.475 $Y2=1.635
r172 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.475 $Y=0.755
+ $X2=0.475 $Y2=1.305
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_152_89# 1 3 11 15 21 26 27 28 29 30 32
+ 35 39
c91 39 0 1.72079e-19 $X=2.415 $Y=0.755
c92 27 0 1.29912e-19 $X=2.33 $Y=1.285
c93 11 0 6.64688e-20 $X=0.835 $Y=0.755
r94 39 41 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=2.415 $Y=0.755
+ $X2=2.515 $Y2=0.755
r95 35 37 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=2.515 $Y=2.955
+ $X2=2.515 $Y2=3.635
r96 33 35 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=2.79
+ $X2=2.515 $Y2=2.955
r97 31 39 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.415 $Y=0.935
+ $X2=2.415 $Y2=0.755
r98 31 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.415 $Y=0.935
+ $X2=2.415 $Y2=1.2
r99 29 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.345 $Y=2.705
+ $X2=2.515 $Y2=2.79
r100 29 30 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.345 $Y=2.705
+ $X2=1.115 $Y2=2.705
r101 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=1.285
+ $X2=2.415 $Y2=1.2
r102 27 28 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.33 $Y=1.285
+ $X2=1.115 $Y2=1.285
r103 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=2.62
+ $X2=1.115 $Y2=2.705
r104 24 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.03 $Y=2.62
+ $X2=1.03 $Y2=1.925
r105 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=1.37
+ $X2=1.115 $Y2=1.285
r106 23 26 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.03 $Y=1.37
+ $X2=1.03 $Y2=1.925
r107 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.925 $X2=1.03 $Y2=1.925
r108 19 21 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.905 $Y=1.925
+ $X2=1.03 $Y2=1.925
r109 17 19 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.835 $Y=1.925
+ $X2=0.905 $Y2=1.925
r110 13 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.09
+ $X2=0.905 $Y2=1.925
r111 13 15 694.798 $w=1.5e-07 $l=1.355e-06 $layer=POLY_cond $X=0.905 $Y=2.09
+ $X2=0.905 $Y2=3.445
r112 9 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=1.76
+ $X2=0.835 $Y2=1.925
r113 9 11 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=0.835 $Y=1.76
+ $X2=0.835 $Y2=0.755
r114 3 37 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=2.605 $X2=2.515 $Y2=3.635
r115 3 35 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=2.605 $X2=2.515 $Y2=2.955
r116 1 41 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.575 $X2=2.515 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%D 3 7 10 14 19
c41 19 0 1.41836e-19 $X=1.915 $Y=1.74
c42 10 0 1.12321e-19 $X=1.915 $Y=1.74
r43 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.915 $Y=1.74
+ $X2=1.915 $Y2=1.74
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.74 $X2=1.915 $Y2=1.74
r45 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.74
+ $X2=1.915 $Y2=1.905
r46 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.74
+ $X2=1.915 $Y2=1.575
r47 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=1.855 $Y=3.235
+ $X2=1.855 $Y2=1.905
r48 3 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.855 $Y=0.835
+ $X2=1.855 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c233 76 0 1.65829e-19 $X=5.355 $Y=2.11
c234 74 0 1.97877e-19 $X=4.36 $Y=2.11
c235 55 0 6.79641e-20 $X=4.11 $Y=2.11
c236 54 0 1.70391e-19 $X=4.42 $Y=2.11
c237 52 0 1.80245e-19 $X=4.025 $Y=1.37
c238 48 0 1.98654e-19 $X=2.755 $Y=1.37
c239 44 0 1.86602e-19 $X=2.67 $Y=2.11
c240 37 0 4.60524e-20 $X=4.505 $Y=2.285
c241 33 0 9.70599e-20 $X=4.025 $Y=1.37
c242 30 0 1.29912e-19 $X=2.755 $Y=1.205
c243 25 0 1.41836e-19 $X=2.275 $Y=2.285
r244 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.65 $Y=2.11
+ $X2=4.505 $Y2=2.11
r245 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.355 $Y=2.11
+ $X2=5.5 $Y2=2.11
r246 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=5.355 $Y=2.11
+ $X2=4.65 $Y2=2.11
r247 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.42 $Y=2.11
+ $X2=2.275 $Y2=2.11
r248 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.36 $Y=2.11
+ $X2=4.505 $Y2=2.11
r249 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=4.36 $Y=2.11
+ $X2=2.42 $Y2=2.11
r250 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.505 $Y=2.11
+ $X2=4.505 $Y2=2.11
r251 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.505 $Y=2.11
+ $X2=4.505 $Y2=2.285
r252 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.275 $Y=2.11
+ $X2=2.275 $Y2=2.11
r253 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.275 $Y=2.11
+ $X2=2.275 $Y2=2.285
r254 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.5 $Y=2.11 $X2=5.5
+ $Y2=2.11
r255 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.5 $Y=2.11
+ $X2=5.5 $Y2=2.285
r256 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.11
+ $X2=4.505 $Y2=2.11
r257 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.42 $Y=2.11
+ $X2=4.11 $Y2=2.11
r258 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=2.025
+ $X2=4.11 $Y2=2.11
r259 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.025 $Y=2.025
+ $X2=4.025 $Y2=1.37
r260 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.755 $Y=2.025
+ $X2=2.755 $Y2=1.37
r261 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.11
+ $X2=2.275 $Y2=2.11
r262 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.67 $Y=2.11
+ $X2=2.755 $Y2=2.025
r263 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.67 $Y=2.11
+ $X2=2.36 $Y2=2.11
r264 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=2.285 $X2=5.5 $Y2=2.285
r265 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=5.382 $Y=1.205
+ $X2=5.382 $Y2=1.355
r266 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=2.285 $X2=4.505 $Y2=2.285
r267 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=2.285
+ $X2=4.505 $Y2=2.45
r268 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.37 $X2=4.025 $Y2=1.37
r269 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.37
+ $X2=4.025 $Y2=1.205
r270 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.37 $X2=2.755 $Y2=1.37
r271 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.37
+ $X2=2.755 $Y2=1.205
r272 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=2.285 $X2=2.275 $Y2=2.285
r273 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=2.285
+ $X2=2.275 $Y2=2.45
r274 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=5.41 $Y=2.12
+ $X2=5.457 $Y2=2.285
r275 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=5.41 $Y=2.12
+ $X2=5.41 $Y2=1.355
r276 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=5.355 $Y=2.45
+ $X2=5.457 $Y2=2.285
r277 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.355 $Y=2.45
+ $X2=5.355 $Y2=3.235
r278 17 40 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.355 $Y=0.835
+ $X2=5.355 $Y2=1.205
r279 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=4.565 $Y=3.235
+ $X2=4.565 $Y2=2.45
r280 10 34 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.965 $Y=0.835
+ $X2=3.965 $Y2=1.205
r281 7 30 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.815 $Y=0.835
+ $X2=2.815 $Y2=1.205
r282 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.215 $Y=3.235
+ $X2=2.215 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_27_115# 1 3 11 15 17 18 21 22 27 31 33
+ 37 43 46 53 55 56 57 59 62
c140 56 0 1.42775e-19 $X=3.11 $Y=1.37
c141 53 0 9.70599e-20 $X=3.345 $Y=1.37
c142 46 0 6.64688e-20 $X=0.26 $Y=0.74
c143 43 0 1.5821e-19 $X=3.345 $Y=2.285
c144 31 0 6.36774e-20 $X=3.605 $Y=3.235
c145 27 0 1.80245e-19 $X=3.605 $Y=0.835
c146 22 0 1.86602e-19 $X=3.25 $Y=2.285
c147 21 0 6.79641e-20 $X=3.53 $Y=2.285
c148 15 0 6.36774e-20 $X=3.175 $Y=3.235
r149 56 62 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.11 $Y=1.37
+ $X2=3.255 $Y2=1.37
r150 56 57 2.24833 $w=1.7e-07 $l=2.335e-06 $layer=MET1_cond $X=3.11 $Y=1.37
+ $X2=0.775 $Y2=1.37
r151 55 59 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.79
+ $X2=0.69 $Y2=1.905
r152 54 57 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.69 $Y=1.455
+ $X2=0.775 $Y2=1.37
r153 54 55 0.322566 $w=1.7e-07 $l=3.35e-07 $layer=MET1_cond $X=0.69 $Y=1.455
+ $X2=0.69 $Y2=1.79
r154 51 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.255 $Y=1.37
+ $X2=3.255 $Y2=1.37
r155 51 53 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=3.255 $Y=1.33
+ $X2=3.345 $Y2=1.33
r156 46 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.26 $Y=0.74
+ $X2=0.26 $Y2=0.91
r157 41 53 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=1.455
+ $X2=3.345 $Y2=1.33
r158 41 43 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.345 $Y=1.455
+ $X2=3.345 $Y2=2.285
r159 37 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.905
+ $X2=0.69 $Y2=1.905
r160 37 39 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=0.69 $Y=1.905
+ $X2=0.69 $Y2=3.615
r161 35 37 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.69 $Y=0.995
+ $X2=0.69 $Y2=1.905
r162 34 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.91
+ $X2=0.26 $Y2=0.91
r163 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=0.91
+ $X2=0.69 $Y2=0.995
r164 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.91
+ $X2=0.345 $Y2=0.91
r165 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.605 $Y=2.42
+ $X2=3.605 $Y2=3.235
r166 25 27 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.605 $Y=1.235
+ $X2=3.605 $Y2=0.835
r167 24 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=2.285 $X2=3.345 $Y2=2.285
r168 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=2.285
+ $X2=3.345 $Y2=2.285
r169 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.53 $Y=2.285
+ $X2=3.605 $Y2=2.42
r170 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=2.285
+ $X2=3.345 $Y2=2.285
r171 20 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.37 $X2=3.345 $Y2=1.37
r172 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=1.37
+ $X2=3.345 $Y2=1.37
r173 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.53 $Y=1.37
+ $X2=3.605 $Y2=1.235
r174 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=1.37
+ $X2=3.345 $Y2=1.37
r175 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=2.42
+ $X2=3.25 $Y2=2.285
r176 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.175 $Y=2.42
+ $X2=3.175 $Y2=3.235
r177 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=1.235
+ $X2=3.25 $Y2=1.37
r178 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.175 $Y=1.235
+ $X2=3.175 $Y2=0.835
r179 3 39 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=3.025 $X2=0.69 $Y2=3.615
r180 1 46 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_428_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 50 54 59 62 66 68 69 74
c196 69 0 2.16443e-19 $X=4.65 $Y=1.74
c197 44 0 3.63706e-19 $X=4.505 $Y=1.74
c198 39 0 1.56563e-19 $X=4.505 $Y=1.74
c199 34 0 1.98654e-19 $X=2.335 $Y=1.28
c200 18 0 1.12321e-19 $X=2.815 $Y=3.235
r201 69 71 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.65 $Y=1.74
+ $X2=4.505 $Y2=1.74
r202 68 74 0.0841272 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=5.405 $Y=1.74
+ $X2=5.52 $Y2=1.74
r203 68 69 0.726976 $w=1.7e-07 $l=7.55e-07 $layer=MET1_cond $X=5.405 $Y=1.74
+ $X2=4.65 $Y2=1.74
r204 66 67 19.0625 $w=1.76e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=1.755
+ $X2=5.845 $Y2=1.755
r205 65 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.74
+ $X2=5.52 $Y2=1.74
r206 65 66 3.46591 $w=1.76e-07 $l=5e-08 $layer=LI1_cond $X=5.52 $Y=1.755
+ $X2=5.57 $Y2=1.755
r207 60 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=2.705
+ $X2=5.845 $Y2=2.705
r208 59 62 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.62
+ $X2=5.845 $Y2=2.705
r209 58 67 0.578974 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=5.845 $Y=1.855
+ $X2=5.845 $Y2=1.755
r210 58 59 47.1364 $w=1.78e-07 $l=7.65e-07 $layer=LI1_cond $X=5.845 $Y=1.855
+ $X2=5.845 $Y2=2.62
r211 54 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.57 $Y=2.955
+ $X2=5.57 $Y2=3.635
r212 52 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=2.79
+ $X2=5.57 $Y2=2.705
r213 52 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=2.79
+ $X2=5.57 $Y2=2.955
r214 48 66 0.927112 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.57 $Y=1.655
+ $X2=5.57 $Y2=1.755
r215 48 50 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.57 $Y=1.655
+ $X2=5.57 $Y2=0.755
r216 44 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.505 $Y=1.74
+ $X2=4.505 $Y2=1.74
r217 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=1.74 $X2=4.505 $Y2=1.74
r218 39 41 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=4.505 $Y=1.74
+ $X2=4.505 $Y2=1.825
r219 39 40 50.6376 $w=2.7e-07 $l=1.75e-07 $layer=POLY_cond $X=4.505 $Y=1.74
+ $X2=4.505 $Y2=1.565
r220 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.215 $Y=1.28
+ $X2=2.335 $Y2=1.28
r221 30 40 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=4.565 $Y=0.835
+ $X2=4.565 $Y2=1.565
r222 27 37 19.8589 $w=1.55e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=1.825
+ $X2=3.965 $Y2=1.825
r223 26 41 15.0071 $w=1.6e-07 $l=1.35e-07 $layer=POLY_cond $X=4.37 $Y=1.825
+ $X2=4.505 $Y2=1.825
r224 26 27 152.942 $w=1.6e-07 $l=3.3e-07 $layer=POLY_cond $X=4.37 $Y=1.825
+ $X2=4.04 $Y2=1.825
r225 22 37 5.77175 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=3.965 $Y=1.905
+ $X2=3.965 $Y2=1.825
r226 22 24 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.965 $Y=1.905
+ $X2=3.965 $Y2=3.235
r227 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.89 $Y=1.82
+ $X2=2.815 $Y2=1.82
r228 20 37 19.8589 $w=1.55e-07 $l=7.74597e-08 $layer=POLY_cond $X=3.89 $Y=1.82
+ $X2=3.965 $Y2=1.825
r229 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.89 $Y=1.82 $X2=2.89
+ $Y2=1.82
r230 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.815 $Y=1.895
+ $X2=2.815 $Y2=1.82
r231 16 18 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=2.815 $Y=1.895
+ $X2=2.815 $Y2=3.235
r232 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.74 $Y=1.82
+ $X2=2.815 $Y2=1.82
r233 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.74 $Y=1.82
+ $X2=2.41 $Y2=1.82
r234 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.335 $Y=1.745
+ $X2=2.41 $Y2=1.82
r235 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.335 $Y=1.355
+ $X2=2.335 $Y2=1.28
r236 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.335 $Y=1.355
+ $X2=2.335 $Y2=1.745
r237 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.215 $Y=1.205
+ $X2=2.215 $Y2=1.28
r238 9 11 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.215 $Y=1.205
+ $X2=2.215 $Y2=0.835
r239 3 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=2.605 $X2=5.57 $Y2=3.635
r240 3 54 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=2.605 $X2=5.57 $Y2=2.955
r241 1 50 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.575 $X2=5.57 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_970_89# 1 3 11 15 23 26 28 32 33 35 36
+ 37 38 40 45 48 51 55 59 63 64 65 67 68 69 74
c198 59 0 6.64688e-20 $X=6.09 $Y=0.74
c199 40 0 1.6261e-19 $X=4.985 $Y=1.71
c200 37 0 8.77106e-20 $X=7.66 $Y=2.375
c201 36 0 1.11496e-19 $X=7.66 $Y=1.32
c202 32 0 2.20654e-19 $X=7.57 $Y=1.71
r203 68 74 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.425 $Y=1.71
+ $X2=7.57 $Y2=1.71
r204 68 69 1.41062 $w=1.7e-07 $l=1.465e-06 $layer=MET1_cond $X=7.425 $Y=1.71
+ $X2=5.96 $Y2=1.71
r205 66 69 0.0700348 $w=1.7e-07 $l=1.17707e-07 $layer=MET1_cond $X=5.882
+ $Y=1.795 $X2=5.96 $Y2=1.71
r206 66 67 0.628358 $w=1.55e-07 $l=5.95e-07 $layer=MET1_cond $X=5.882 $Y=1.795
+ $X2=5.882 $Y2=2.39
r207 65 71 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.13 $Y=2.48
+ $X2=4.985 $Y2=2.48
r208 64 67 0.0700348 $w=1.7e-07 $l=1.34681e-07 $layer=MET1_cond $X=5.785 $Y=2.48
+ $X2=5.882 $Y2=2.39
r209 64 65 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=5.785 $Y=2.48
+ $X2=5.13 $Y2=2.48
r210 59 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.09 $Y=0.74
+ $X2=6.09 $Y2=0.91
r211 55 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.57 $Y=1.71
+ $X2=7.57 $Y2=1.71
r212 53 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=1.71
+ $X2=6.52 $Y2=1.71
r213 53 55 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=6.605 $Y=1.71
+ $X2=7.57 $Y2=1.71
r214 49 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.795
+ $X2=6.52 $Y2=1.71
r215 49 51 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=6.52 $Y=1.795
+ $X2=6.52 $Y2=3.615
r216 48 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.625
+ $X2=6.52 $Y2=1.71
r217 47 48 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.52 $Y=0.995
+ $X2=6.52 $Y2=1.625
r218 46 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.91
+ $X2=6.09 $Y2=0.91
r219 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.435 $Y=0.91
+ $X2=6.52 $Y2=0.995
r220 45 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.435 $Y=0.91
+ $X2=6.175 $Y2=0.91
r221 43 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.985 $Y=2.48
+ $X2=4.985 $Y2=2.48
r222 40 43 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.985 $Y=1.71
+ $X2=4.985 $Y2=2.48
r223 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=2.375
+ $X2=7.66 $Y2=2.525
r224 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=1.17 $X2=7.66
+ $Y2=1.32
r225 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.635 $Y=1.875
+ $X2=7.635 $Y2=2.375
r226 33 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.635 $Y=1.545
+ $X2=7.635 $Y2=1.32
r227 32 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=1.71 $X2=7.57 $Y2=1.71
r228 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=1.71
+ $X2=7.572 $Y2=1.875
r229 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=1.71
+ $X2=7.572 $Y2=1.545
r230 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.71 $X2=4.985 $Y2=1.71
r231 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.71
+ $X2=4.985 $Y2=1.875
r232 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.71
+ $X2=4.985 $Y2=1.545
r233 26 38 228.147 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.685 $Y=3.235
+ $X2=7.685 $Y2=2.525
r234 23 35 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.685 $Y=0.835
+ $X2=7.685 $Y2=1.17
r235 15 30 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=4.925 $Y=3.235
+ $X2=4.925 $Y2=1.875
r236 11 29 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.925 $Y=0.835
+ $X2=4.925 $Y2=1.545
r237 3 51 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=3.025 $X2=6.52 $Y2=3.615
r238 1 59 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.965
+ $Y=0.575 $X2=6.09 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%A_808_115# 1 3 11 15 20 24 26 27 30 34
+ 37 42 45 46 47 48 55
c145 47 0 1.56563e-19 $X=5.955 $Y=1.37
c146 46 0 1.5821e-19 $X=3.83 $Y=1.37
c147 42 0 1.71621e-19 $X=4.265 $Y=0.755
c148 37 0 1.08672e-19 $X=6.1 $Y=1.37
c149 24 0 1.57671e-19 $X=3.685 $Y=1.37
r150 48 53 0.0841272 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.48 $Y=1.37
+ $X2=4.365 $Y2=1.37
r151 47 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.955 $Y=1.37
+ $X2=6.1 $Y2=1.37
r152 47 48 1.42025 $w=1.7e-07 $l=1.475e-06 $layer=MET1_cond $X=5.955 $Y=1.37
+ $X2=4.48 $Y2=1.37
r153 46 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.83 $Y=1.37
+ $X2=3.685 $Y2=1.37
r154 45 53 0.0873352 $w=2.3e-07 $l=1.2e-07 $layer=MET1_cond $X=4.245 $Y=1.37
+ $X2=4.365 $Y2=1.37
r155 45 46 0.399596 $w=1.7e-07 $l=4.15e-07 $layer=MET1_cond $X=4.245 $Y=1.37
+ $X2=3.83 $Y2=1.37
r156 42 44 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=4.272 $Y=0.755
+ $X2=4.272 $Y2=1.035
r157 37 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.1 $Y=1.37 $X2=6.1
+ $Y2=1.37
r158 34 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.365 $Y=1.37
+ $X2=4.365 $Y2=1.37
r159 34 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.365 $Y=1.37
+ $X2=4.365 $Y2=1.035
r160 28 30 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=4.265 $Y=2.79
+ $X2=4.265 $Y2=3.295
r161 26 28 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=2.705
+ $X2=4.265 $Y2=2.79
r162 26 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=2.705
+ $X2=3.77 $Y2=2.705
r163 24 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=1.37
+ $X2=3.685 $Y2=1.37
r164 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=2.62
+ $X2=3.77 $Y2=2.705
r165 22 24 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.685 $Y=2.62
+ $X2=3.685 $Y2=1.37
r166 18 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.1
+ $Y=1.37 $X2=6.1 $Y2=1.37
r167 18 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.1 $Y=1.37
+ $X2=6.305 $Y2=1.37
r168 13 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.535
+ $X2=6.305 $Y2=1.37
r169 13 15 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=6.305 $Y=1.535
+ $X2=6.305 $Y2=3.445
r170 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=1.37
r171 9 11 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=0.755
r172 3 30 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=4.04
+ $Y=2.605 $X2=4.265 $Y2=3.295
r173 1 42 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.575 $X2=4.265 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c83 42 0 8.77106e-20 $X=7.475 $Y=2.48
c84 33 0 9.99996e-20 $X=7.97 $Y=2.285
c85 31 0 1.20654e-19 $X=7.97 $Y=1.37
c86 18 0 1.98165e-19 $X=8.055 $Y=1.915
r87 40 42 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=7.47 $Y=2.48
+ $X2=7.475 $Y2=2.48
r88 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.055 $Y=2.2
+ $X2=8.055 $Y2=1.915
r89 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.055 $Y=1.455
+ $X2=8.055 $Y2=1.915
r90 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=2.285
+ $X2=8.055 $Y2=2.2
r91 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=2.285
+ $X2=7.555 $Y2=2.285
r92 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=1.37
+ $X2=8.055 $Y2=1.455
r93 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=1.37
+ $X2=7.555 $Y2=1.37
r94 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.47 $Y=2.48
+ $X2=7.47 $Y2=2.48
r95 27 29 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.47 $Y=2.48
+ $X2=7.47 $Y2=3.265
r96 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=2.37
+ $X2=7.555 $Y2=2.285
r97 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.47 $Y=2.37
+ $X2=7.47 $Y2=2.48
r98 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=1.285
+ $X2=7.555 $Y2=1.37
r99 21 23 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.47 $Y=1.285
+ $X2=7.47 $Y2=0.74
r100 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=1.915 $X2=8.055 $Y2=1.915
r101 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=1.915
+ $X2=8.055 $Y2=2.08
r102 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=1.915
+ $X2=8.055 $Y2=1.75
r103 15 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=8.115 $Y=3.235
+ $X2=8.115 $Y2=2.08
r104 11 19 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=8.115 $Y=0.835
+ $X2=8.115 $Y2=1.75
r105 3 29 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=2.605 $X2=7.47 $Y2=3.265
r106 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__DFFS_1%Q 1 3 11 15 18 21 25 28
r20 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=2.807
+ $X2=8.445 $Y2=2.807
r21 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.325 $Y=2.85
+ $X2=8.325 $Y2=2.85
r22 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=8.325 $Y=2.807
+ $X2=8.33 $Y2=2.807
r23 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=1.035
+ $X2=8.445 $Y2=1.035
r24 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.445 $Y=2.68
+ $X2=8.445 $Y2=2.807
r25 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=1.12
+ $X2=8.445 $Y2=1.035
r26 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=8.445 $Y=1.12
+ $X2=8.445 $Y2=2.68
r27 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.33 $Y=2.935
+ $X2=8.33 $Y2=2.807
r28 13 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.33 $Y=2.935
+ $X2=8.33 $Y2=3.265
r29 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=0.95 $X2=8.33
+ $Y2=1.035
r30 9 11 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.33 $Y=0.95 $X2=8.33
+ $Y2=0.74
r31 3 15 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=2.605 $X2=8.33 $Y2=3.265
r32 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.575 $X2=8.33 $Y2=0.74
.ends

