* File: sky130_osu_sc_18T_ls__dff_1.pex.spice
* Created: Thu Oct 29 17:35:21 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%GND 1 2 3 4 5 56 60 62 72 74 84 86 93 95
+ 102 106 119 121
c171 56 0 1.27355e-19 $X=-0.045 $Y=0
r172 119 121 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r173 106 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.152
+ $X2=0.715 $Y2=0.152
r174 100 102 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.545 $Y=0.305
+ $X2=6.545 $Y2=0.825
r175 91 93 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.165 $Y=0.305
+ $X2=5.165 $Y2=0.825
r176 87 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.152
+ $X2=4.215 $Y2=0.152
r177 82 111 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.152
r178 82 84 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.215 $Y=0.305
+ $X2=4.215 $Y2=0.825
r179 74 111 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.152
+ $X2=4.215 $Y2=0.152
r180 70 72 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.465 $Y=0.305
+ $X2=2.465 $Y2=0.825
r181 63 107 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.152
+ $X2=0.715 $Y2=0.152
r182 58 107 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.152
r183 58 60 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.715 $Y=0.305
+ $X2=0.715 $Y2=0.825
r184 56 100 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.545 $Y2=0.305
r185 56 95 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.152
+ $X2=6.46 $Y2=0.152
r186 56 106 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.63 $Y2=0.152
r187 56 121 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.17
+ $X2=6.46 $Y2=0.17
r188 56 119 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r189 56 91 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.165 $Y2=0.305
r190 56 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.08 $Y2=0.152
r191 56 96 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.152
+ $X2=5.25 $Y2=0.152
r192 56 70 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.465 $Y2=0.305
r193 56 62 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.38 $Y2=0.152
r194 56 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.152
+ $X2=2.55 $Y2=0.152
r195 56 95 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.46 $Y2=0.152
r196 56 96 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.25 $Y2=0.152
r197 56 86 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=5.08 $Y2=0.152
r198 56 87 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.42 $Y=0.152
+ $X2=4.3 $Y2=0.152
r199 56 74 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.13 $Y2=0.152
r200 56 75 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.55 $Y2=0.152
r201 56 62 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.38 $Y2=0.152
r202 56 63 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.8 $Y2=0.152
r203 5 102 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.405
+ $Y=0.575 $X2=6.545 $Y2=0.825
r204 4 93 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=5.04
+ $Y=0.575 $X2=5.165 $Y2=0.825
r205 3 84 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.075
+ $Y=0.575 $X2=4.215 $Y2=0.825
r206 2 72 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.575 $X2=2.465 $Y2=0.825
r207 1 60 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.575 $X2=0.715 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%VDD 1 2 3 4 5 46 50 54 62 66 74 78 84 88
+ 94 100 108 113 114
c99 94 0 1.98165e-19 $X=6.545 $Y=3.455
c100 50 0 5.41559e-20 $X=0.715 $Y=3.795
c101 1 0 1.59851e-19 $X=0.575 $Y=3.085
r102 113 114 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=6.49
+ $X2=6.46 $Y2=6.49
r103 108 113 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=6.46 $Y2=6.507
r104 108 117 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r105 100 117 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=0.63 $Y=6.507
+ $X2=0.34 $Y2=6.507
r106 100 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=6.507
+ $X2=0.715 $Y2=6.507
r107 94 97 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.545 $Y=3.455
+ $X2=6.545 $Y2=5.835
r108 92 114 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=6.355
+ $X2=6.545 $Y2=6.507
r109 92 97 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.545 $Y=6.355
+ $X2=6.545 $Y2=5.835
r110 89 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.25 $Y=6.507
+ $X2=5.165 $Y2=6.507
r111 89 91 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=5.25 $Y=6.507
+ $X2=5.78 $Y2=6.507
r112 88 114 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=6.507
+ $X2=6.545 $Y2=6.507
r113 88 91 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.46 $Y=6.507
+ $X2=5.78 $Y2=6.507
r114 84 87 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=5.165 $Y=3.795
+ $X2=5.165 $Y2=5.835
r115 82 106 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.165 $Y=6.355
+ $X2=5.165 $Y2=6.507
r116 82 87 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.165 $Y=6.355
+ $X2=5.165 $Y2=5.835
r117 79 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=6.507
+ $X2=4.215 $Y2=6.507
r118 79 81 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=4.3 $Y=6.507
+ $X2=4.42 $Y2=6.507
r119 78 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=6.507
+ $X2=5.165 $Y2=6.507
r120 78 81 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.08 $Y=6.507
+ $X2=4.42 $Y2=6.507
r121 74 77 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.215 $Y=3.455
+ $X2=4.215 $Y2=5.835
r122 72 104 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.215 $Y=6.355
+ $X2=4.215 $Y2=6.507
r123 72 77 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.215 $Y=6.355
+ $X2=4.215 $Y2=5.835
r124 69 71 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=6.507
+ $X2=3.74 $Y2=6.507
r125 67 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=6.507
+ $X2=2.465 $Y2=6.507
r126 67 69 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=2.55 $Y=6.507
+ $X2=3.06 $Y2=6.507
r127 66 104 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=6.507
+ $X2=4.215 $Y2=6.507
r128 66 71 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=4.13 $Y=6.507
+ $X2=3.74 $Y2=6.507
r129 62 65 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.465 $Y=3.795
+ $X2=2.465 $Y2=5.835
r130 60 103 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.465 $Y=6.355
+ $X2=2.465 $Y2=6.507
r131 60 65 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.465 $Y=6.355
+ $X2=2.465 $Y2=5.835
r132 57 59 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r133 55 101 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=6.507
+ $X2=0.715 $Y2=6.507
r134 55 57 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=0.8 $Y=6.507
+ $X2=1.02 $Y2=6.507
r135 54 103 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=6.507
+ $X2=2.465 $Y2=6.507
r136 54 59 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=6.507
+ $X2=1.7 $Y2=6.507
r137 50 53 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.715 $Y=3.795
+ $X2=0.715 $Y2=5.835
r138 48 101 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.715 $Y=6.355
+ $X2=0.715 $Y2=6.507
r139 48 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.715 $Y=6.355
+ $X2=0.715 $Y2=5.835
r140 46 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=6.355 $X2=6.46 $Y2=6.44
r141 46 117 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r142 46 106 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=6.355 $X2=5.1 $Y2=6.44
r143 46 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r144 46 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=6.355 $X2=5.78 $Y2=6.44
r145 46 81 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r146 46 71 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r147 46 69 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r148 46 59 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r149 46 57 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r150 5 97 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.405
+ $Y=3.085 $X2=6.545 $Y2=5.835
r151 5 94 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.405
+ $Y=3.085 $X2=6.545 $Y2=3.455
r152 4 87 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=5.04
+ $Y=3.085 $X2=5.165 $Y2=5.835
r153 4 84 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=5.04
+ $Y=3.085 $X2=5.165 $Y2=3.795
r154 3 77 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.075
+ $Y=3.085 $X2=4.215 $Y2=5.835
r155 3 74 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.075
+ $Y=3.085 $X2=4.215 $Y2=3.455
r156 2 65 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=2.325 $Y=3.085 $X2=2.465 $Y2=5.835
r157 2 62 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=2.325 $Y=3.085 $X2=2.465 $Y2=3.795
r158 1 53 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=0.575 $Y=3.085 $X2=0.715 $Y2=5.835
r159 1 50 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=0.575 $Y=3.085 $X2=0.715 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%A_75_344# 1 2 11 15 18 22 23 24 25 26 28
+ 31 35 40 41 42 45 47
c86 41 0 5.41559e-20 $X=0.51 $Y=2.765
c87 23 0 1.29912e-19 $X=1.405 $Y=1.765
c88 22 0 1.59851e-19 $X=0.625 $Y=3.1
r89 44 45 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.582 $Y=1.245
+ $X2=1.582 $Y2=1.415
r90 41 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.765
+ $X2=0.51 $Y2=2.93
r91 41 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.765
+ $X2=0.51 $Y2=2.6
r92 40 43 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.765
+ $X2=0.567 $Y2=2.93
r93 40 42 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=2.765
+ $X2=0.567 $Y2=2.6
r94 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=2.765 $X2=0.51 $Y2=2.765
r95 35 37 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.59 $Y=3.455
+ $X2=1.59 $Y2=5.835
r96 33 35 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=1.59 $Y=3.375 $X2=1.59
+ $Y2=3.455
r97 31 44 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.59 $Y=0.825
+ $X2=1.59 $Y2=1.245
r98 28 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.49 $Y=1.68
+ $X2=1.49 $Y2=1.415
r99 25 33 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=1.42 $Y=3.185
+ $X2=1.59 $Y2=3.375
r100 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.42 $Y=3.185
+ $X2=0.71 $Y2=3.185
r101 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.765
+ $X2=1.49 $Y2=1.68
r102 23 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.405 $Y=1.765
+ $X2=0.71 $Y2=1.765
r103 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=3.1
+ $X2=0.71 $Y2=3.185
r104 22 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.625 $Y=3.1
+ $X2=0.625 $Y2=2.93
r105 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.85
+ $X2=0.71 $Y2=1.765
r106 19 42 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.625 $Y=1.85
+ $X2=0.625 $Y2=2.6
r107 18 47 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.45 $Y=1.87
+ $X2=0.45 $Y2=2.6
r108 17 18 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.475 $Y=1.72
+ $X2=0.475 $Y2=1.87
r109 15 48 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.5 $Y=4.585
+ $X2=0.5 $Y2=2.93
r110 11 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.5 $Y=1.075
+ $X2=0.5 $Y2=1.72
r111 2 37 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.365
+ $Y=3.085 $X2=1.59 $Y2=5.835
r112 2 35 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.365
+ $Y=3.085 $X2=1.59 $Y2=3.455
r113 1 31 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.365
+ $Y=0.575 $X2=1.59 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%D 3 7 10 12 16
c43 16 0 1.12321e-19 $X=0.99 $Y=2.22
c44 10 0 1.41836e-19 $X=0.99 $Y=2.22
r45 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=2.22
+ $X2=0.99 $Y2=2.385
r46 16 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=2.22
+ $X2=0.99 $Y2=2.055
r47 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.22 $X2=0.99 $Y2=2.22
r48 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=2.22
+ $X2=0.99 $Y2=2.22
r49 7 18 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.93 $Y=4.585
+ $X2=0.93 $Y2=2.385
r50 3 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.93 $Y=1.075
+ $X2=0.93 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%CK 3 7 10 13 17 18 20 23 24 25 26 30 31
+ 35 36 38 39 40 41 42 43 46 50 52 54 59 63 66 70
c213 63 0 1.29912e-19 $X=1.83 $Y=1.685
c214 59 0 1.41836e-19 $X=1.35 $Y=2.765
c215 39 0 6.79641e-20 $X=3.185 $Y=2.59
c216 30 0 1.98654e-19 $X=1.83 $Y=1.85
c217 26 0 1.86602e-19 $X=1.745 $Y=2.59
r218 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=2.765 $X2=4.575 $Y2=2.765
r219 70 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=2.765
+ $X2=3.58 $Y2=2.93
r220 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=2.765 $X2=3.58 $Y2=2.765
r221 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=2.765
+ $X2=1.35 $Y2=2.93
r222 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=2.765 $X2=1.35 $Y2=2.765
r223 54 74 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.59
+ $X2=4.575 $Y2=2.765
r224 52 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.575 $Y=2.59
+ $X2=4.575 $Y2=2.59
r225 50 69 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.58 $Y=2.59
+ $X2=3.58 $Y2=2.765
r226 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.59
+ $X2=3.58 $Y2=2.59
r227 46 58 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.35 $Y=2.59
+ $X2=1.35 $Y2=2.765
r228 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.35 $Y=2.59
+ $X2=1.35 $Y2=2.59
r229 43 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.725 $Y=2.59
+ $X2=3.58 $Y2=2.59
r230 42 52 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.43 $Y=2.59
+ $X2=4.575 $Y2=2.59
r231 42 43 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=4.43 $Y=2.59
+ $X2=3.725 $Y2=2.59
r232 41 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.495 $Y=2.59
+ $X2=1.35 $Y2=2.59
r233 40 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.435 $Y=2.59
+ $X2=3.58 $Y2=2.59
r234 40 41 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=3.435 $Y=2.59
+ $X2=1.495 $Y2=2.59
r235 38 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.59
+ $X2=3.58 $Y2=2.59
r236 38 39 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.495 $Y=2.59
+ $X2=3.185 $Y2=2.59
r237 36 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.85
+ $X2=3.1 $Y2=1.685
r238 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.85 $X2=3.1 $Y2=1.85
r239 33 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.505
+ $X2=3.185 $Y2=2.59
r240 33 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.1 $Y=2.505
+ $X2=3.1 $Y2=1.85
r241 31 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.85
+ $X2=1.83 $Y2=1.685
r242 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.85 $X2=1.83 $Y2=1.85
r243 28 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.83 $Y=2.505
+ $X2=1.83 $Y2=1.85
r244 27 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.59
+ $X2=1.35 $Y2=2.59
r245 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=2.59
+ $X2=1.83 $Y2=2.505
r246 26 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.745 $Y=2.59
+ $X2=1.435 $Y2=2.59
r247 24 25 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=4.457 $Y=1.685
+ $X2=4.457 $Y2=1.835
r248 23 75 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=4.485 $Y=2.6
+ $X2=4.532 $Y2=2.765
r249 23 25 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.485 $Y=2.6
+ $X2=4.485 $Y2=1.835
r250 18 75 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=4.43 $Y=2.93
+ $X2=4.532 $Y2=2.765
r251 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=4.43 $Y=2.93
+ $X2=4.43 $Y2=4.585
r252 17 24 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.43 $Y=1.075
+ $X2=4.43 $Y2=1.685
r253 13 72 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.64 $Y=4.585
+ $X2=3.64 $Y2=2.93
r254 10 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.04 $Y=1.075
+ $X2=3.04 $Y2=1.685
r255 7 63 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.89 $Y=1.075
+ $X2=1.89 $Y2=1.685
r256 3 61 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.29 $Y=4.585
+ $X2=1.29 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%A_32_115# 1 2 9 13 17 21 23 24 25 26 28
+ 29 31 35 41 46 48 49 55 56
c115 41 0 1.5821e-19 $X=2.42 $Y=2.765
c116 26 0 6.79641e-20 $X=2.605 $Y=2.765
c117 24 0 1.86602e-19 $X=2.325 $Y=2.765
c118 21 0 6.36774e-20 $X=2.68 $Y=4.585
c119 13 0 6.36774e-20 $X=2.25 $Y=4.585
r120 56 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.85 $X2=2.42 $Y2=1.85
r121 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.33 $Y=1.85
+ $X2=2.33 $Y2=1.85
r122 49 51 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.43 $Y=1.85
+ $X2=0.285 $Y2=1.85
r123 48 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.185 $Y=1.85
+ $X2=2.33 $Y2=1.85
r124 48 49 1.68986 $w=1.7e-07 $l=1.755e-06 $layer=MET1_cond $X=2.185 $Y=1.85
+ $X2=0.43 $Y2=1.85
r125 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=2.765 $X2=2.42 $Y2=2.765
r126 39 56 2.3025 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.42 $Y=1.935
+ $X2=2.33 $Y2=1.81
r127 39 41 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.42 $Y=1.935
+ $X2=2.42 $Y2=2.765
r128 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.285 $Y=3.455
+ $X2=0.285 $Y2=5.835
r129 33 46 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.285 $Y=3.345
+ $X2=0.285 $Y2=3.242
r130 33 35 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.285 $Y=3.345
+ $X2=0.285 $Y2=3.455
r131 29 62 4.81931 $w=2.73e-07 $l=1.15e-07 $layer=LI1_cond $X=0.285 $Y=1.797
+ $X2=0.17 $Y2=1.797
r132 29 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.285 $Y=1.85
+ $X2=0.285 $Y2=1.85
r133 29 31 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.285 $Y=1.66
+ $X2=0.285 $Y2=0.825
r134 28 46 6.22173 $w=2.03e-07 $l=1.15e-07 $layer=LI1_cond $X=0.17 $Y=3.242
+ $X2=0.285 $Y2=3.242
r135 27 62 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.17 $Y=1.935
+ $X2=0.17 $Y2=1.797
r136 27 28 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=0.17 $Y=1.935
+ $X2=0.17 $Y2=3.14
r137 26 42 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=2.765
+ $X2=2.42 $Y2=2.765
r138 25 60 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.605 $Y=1.85
+ $X2=2.42 $Y2=1.85
r139 24 42 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=2.765
+ $X2=2.42 $Y2=2.765
r140 23 60 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=2.325 $Y=1.85
+ $X2=2.42 $Y2=1.85
r141 19 26 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.68 $Y=2.9
+ $X2=2.605 $Y2=2.765
r142 19 21 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=2.68 $Y=2.9
+ $X2=2.68 $Y2=4.585
r143 15 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.68 $Y=1.715
+ $X2=2.605 $Y2=1.85
r144 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.68 $Y=1.715
+ $X2=2.68 $Y2=1.075
r145 11 24 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=2.9
+ $X2=2.325 $Y2=2.765
r146 11 13 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=2.25 $Y=2.9
+ $X2=2.25 $Y2=4.585
r147 7 23 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.25 $Y=1.715
+ $X2=2.325 $Y2=1.85
r148 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.25 $Y=1.715 $X2=2.25
+ $Y2=1.075
r149 2 37 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.16
+ $Y=3.085 $X2=0.285 $Y2=5.835
r150 2 35 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.16
+ $Y=3.085 $X2=0.285 $Y2=3.455
r151 1 31 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.575 $X2=0.285 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%A_243_89# 1 2 7 9 11 12 13 16 18 22 24 27
+ 30 33 35 36 37 40 44 47 50 55 56 59 63 66
c174 33 0 1.98654e-19 $X=1.41 $Y=1.76
c175 16 0 1.12321e-19 $X=1.89 $Y=4.585
r176 61 63 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=3.185
+ $X2=4.915 $Y2=3.185
r177 57 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.645 $Y=2.19
+ $X2=4.915 $Y2=2.19
r178 55 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=3.1
+ $X2=4.915 $Y2=3.185
r179 54 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.275
+ $X2=4.915 $Y2=2.19
r180 54 55 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.915 $Y=2.275
+ $X2=4.915 $Y2=3.1
r181 50 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.645 $Y=3.455
+ $X2=4.645 $Y2=5.835
r182 48 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=3.27
+ $X2=4.645 $Y2=3.185
r183 48 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.645 $Y=3.27
+ $X2=4.645 $Y2=3.455
r184 47 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=2.105
+ $X2=4.645 $Y2=2.19
r185 46 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.935
+ $X2=4.645 $Y2=1.85
r186 46 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.645 $Y=1.935
+ $X2=4.645 $Y2=2.105
r187 42 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=1.85
r188 42 44 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=0.825
r189 40 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.85
+ $X2=3.58 $Y2=2.015
r190 40 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.85
+ $X2=3.58 $Y2=1.685
r191 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.85 $X2=3.58 $Y2=1.85
r192 37 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=1.85
+ $X2=4.645 $Y2=1.85
r193 37 39 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.56 $Y=1.85
+ $X2=3.58 $Y2=1.85
r194 31 33 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.29 $Y=1.76
+ $X2=1.41 $Y2=1.76
r195 30 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.64 $Y=1.075
+ $X2=3.64 $Y2=1.685
r196 27 67 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.52 $Y=2.225
+ $X2=3.52 $Y2=2.015
r197 25 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.115 $Y=2.3
+ $X2=3.04 $Y2=2.3
r198 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.445 $Y=2.3
+ $X2=3.52 $Y2=2.225
r199 24 25 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.445 $Y=2.3
+ $X2=3.115 $Y2=2.3
r200 20 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.04 $Y=2.375
+ $X2=3.04 $Y2=2.3
r201 20 22 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=3.04 $Y=2.375
+ $X2=3.04 $Y2=4.585
r202 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=2.3
+ $X2=1.89 $Y2=2.3
r203 18 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.965 $Y=2.3
+ $X2=3.04 $Y2=2.3
r204 18 19 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.965 $Y=2.3
+ $X2=1.965 $Y2=2.3
r205 14 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=2.375
+ $X2=1.89 $Y2=2.3
r206 14 16 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=1.89 $Y=2.375
+ $X2=1.89 $Y2=4.585
r207 12 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=2.3
+ $X2=1.89 $Y2=2.3
r208 12 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.815 $Y=2.3
+ $X2=1.485 $Y2=2.3
r209 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=2.225
+ $X2=1.485 $Y2=2.3
r210 10 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.835
+ $X2=1.41 $Y2=1.76
r211 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.41 $Y=1.835
+ $X2=1.41 $Y2=2.225
r212 7 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.685
+ $X2=1.29 $Y2=1.76
r213 7 9 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.29 $Y=1.685
+ $X2=1.29 $Y2=1.075
r214 2 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.505
+ $Y=3.085 $X2=4.645 $Y2=5.835
r215 2 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.505
+ $Y=3.085 $X2=4.645 $Y2=3.455
r216 1 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.505
+ $Y=0.575 $X2=4.645 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%A_785_89# 1 2 9 13 21 24 25 26 27 28 31
+ 35 40 41 42 45 48 49 53 58 59
c131 58 0 2.20654e-19 $X=6.215 $Y=2.19
c132 27 0 8.77106e-20 $X=6.305 $Y=2.855
r133 58 60 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.217 $Y=2.19
+ $X2=6.217 $Y2=2.355
r134 58 59 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.217 $Y=2.19
+ $X2=6.217 $Y2=2.025
r135 53 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=2.19
+ $X2=4.06 $Y2=2.355
r136 53 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=2.19
+ $X2=4.06 $Y2=2.025
r137 49 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=2.19 $X2=6.215 $Y2=2.19
r138 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=2.19
+ $X2=6.215 $Y2=2.19
r139 45 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=2.19 $X2=4.06 $Y2=2.19
r140 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.06 $Y=2.19
+ $X2=4.06 $Y2=2.19
r141 42 44 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.205 $Y=2.19
+ $X2=4.06 $Y2=2.19
r142 41 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.07 $Y=2.19
+ $X2=6.215 $Y2=2.19
r143 41 42 1.79578 $w=1.7e-07 $l=1.865e-06 $layer=MET1_cond $X=6.07 $Y=2.19
+ $X2=4.205 $Y2=2.19
r144 39 49 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.68 $Y=2.19
+ $X2=6.215 $Y2=2.19
r145 39 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=2.19
+ $X2=5.595 $Y2=2.19
r146 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.595 $Y=3.455
+ $X2=5.595 $Y2=5.835
r147 33 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=2.275
+ $X2=5.595 $Y2=2.19
r148 33 35 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=5.595 $Y=2.275
+ $X2=5.595 $Y2=3.455
r149 29 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=2.105
+ $X2=5.595 $Y2=2.19
r150 29 31 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=5.595 $Y=2.105
+ $X2=5.595 $Y2=0.825
r151 27 28 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=2.855
+ $X2=6.305 $Y2=3.005
r152 27 60 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.28 $Y=2.855
+ $X2=6.28 $Y2=2.355
r153 26 59 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.28 $Y=1.8
+ $X2=6.28 $Y2=2.025
r154 25 26 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.305 $Y=1.65
+ $X2=6.305 $Y2=1.8
r155 24 28 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=6.33 $Y=4.585
+ $X2=6.33 $Y2=3.005
r156 21 25 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.33 $Y=1.075
+ $X2=6.33 $Y2=1.65
r157 13 55 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=4 $Y=4.585 $X2=4
+ $Y2=2.355
r158 9 54 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4 $Y=1.075 $X2=4
+ $Y2=2.025
r159 2 37 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5.455
+ $Y=3.085 $X2=5.595 $Y2=5.835
r160 2 35 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5.455
+ $Y=3.085 $X2=5.595 $Y2=3.455
r161 1 31 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.455
+ $Y=0.575 $X2=5.595 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%A_623_115# 1 2 7 9 12 14 15 16 17 20 24
+ 30 31 34 37 38 44
c115 34 0 1.57671e-19 $X=2.76 $Y=1.85
c116 31 0 1.5821e-19 $X=2.905 $Y=1.85
r117 42 44 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.175 $Y=1.85
+ $X2=5.38 $Y2=1.85
r118 38 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.85 $X2=5.175 $Y2=1.85
r119 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.85
+ $X2=5.175 $Y2=1.85
r120 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.76 $Y=1.85
+ $X2=2.76 $Y2=1.85
r121 31 33 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.905 $Y=1.85
+ $X2=2.76 $Y2=1.85
r122 30 37 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.85
+ $X2=5.175 $Y2=1.85
r123 30 31 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=5.03 $Y=1.85
+ $X2=2.905 $Y2=1.85
r124 29 34 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.76 $Y=3.1
+ $X2=2.76 $Y2=1.85
r125 28 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.76 $Y=1.515
+ $X2=2.76 $Y2=1.85
r126 24 26 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=3.34 $Y=3.455
+ $X2=3.34 $Y2=5.835
r127 22 24 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=3.34 $Y=3.27
+ $X2=3.34 $Y2=3.455
r128 18 20 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=3.34 $Y=1.345
+ $X2=3.34 $Y2=0.825
r129 17 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.845 $Y=3.185
+ $X2=2.76 $Y2=3.1
r130 16 22 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=3.185
+ $X2=3.34 $Y2=3.27
r131 16 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=3.185
+ $X2=2.845 $Y2=3.185
r132 15 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.845 $Y=1.43
+ $X2=2.76 $Y2=1.515
r133 14 18 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.17 $Y=1.43
+ $X2=3.34 $Y2=1.345
r134 14 15 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.17 $Y=1.43
+ $X2=2.845 $Y2=1.43
r135 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=2.015
+ $X2=5.38 $Y2=1.85
r136 10 12 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=5.38 $Y=2.015
+ $X2=5.38 $Y2=4.585
r137 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.685
+ $X2=5.38 $Y2=1.85
r138 7 9 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.38 $Y=1.685
+ $X2=5.38 $Y2=1.075
r139 2 26 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=3.115
+ $Y=3.085 $X2=3.34 $Y2=5.835
r140 2 24 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=3.115
+ $Y=3.085 $X2=3.34 $Y2=3.455
r141 1 20 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=3.115
+ $Y=0.575 $X2=3.34 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%QN 1 2 9 13 17 19 20 21 22 26 27 31 32
c75 32 0 8.77106e-20 $X=6.12 $Y=2.96
c76 27 0 1.98165e-19 $X=6.7 $Y=2.395
c77 21 0 9.99996e-20 $X=6.615 $Y=2.765
c78 19 0 1.20654e-19 $X=6.615 $Y=1.85
r79 39 41 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.115 $Y=3.455
+ $X2=6.115 $Y2=5.835
r80 31 39 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.115 $Y=2.96
+ $X2=6.115 $Y2=3.455
r81 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.115 $Y=2.96
+ $X2=6.115 $Y2=2.96
r82 28 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.115 $Y=2.85
+ $X2=6.115 $Y2=2.96
r83 27 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.395
+ $X2=6.7 $Y2=2.56
r84 27 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=2.395
+ $X2=6.7 $Y2=2.23
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=2.395 $X2=6.7 $Y2=2.395
r86 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.7 $Y=2.68 $X2=6.7
+ $Y2=2.395
r87 23 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.7 $Y=1.935 $X2=6.7
+ $Y2=2.395
r88 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.2 $Y=2.765
+ $X2=6.115 $Y2=2.85
r89 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=2.765
+ $X2=6.7 $Y2=2.68
r90 21 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=2.765
+ $X2=6.2 $Y2=2.765
r91 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.615 $Y=1.85
+ $X2=6.7 $Y2=1.935
r92 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.615 $Y=1.85
+ $X2=6.2 $Y2=1.85
r93 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=1.765
+ $X2=6.2 $Y2=1.85
r94 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.115 $Y=1.765
+ $X2=6.115 $Y2=0.825
r95 13 36 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=6.76 $Y=4.585
+ $X2=6.76 $Y2=2.56
r96 9 35 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=6.76 $Y=1.075
+ $X2=6.76 $Y2=2.23
r97 2 41 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=5.99
+ $Y=3.085 $X2=6.115 $Y2=5.835
r98 2 39 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=5.99
+ $Y=3.085 $X2=6.115 $Y2=3.455
r99 1 17 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=5.99
+ $Y=0.575 $X2=6.115 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFF_1%Q 1 2 9 12 15 20 23 30
r20 25 30 163.428 $w=1.68e-07 $l=2.505e-06 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=6.975 $Y2=5.835
r21 23 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.975 $Y=3.33
+ $X2=6.975 $Y2=3.33
r22 17 20 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=3.245
+ $X2=7.09 $Y2=3.245
r23 17 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=3.245
+ $X2=6.975 $Y2=3.33
r24 13 15 7.08586 $w=1.78e-07 $l=1.15e-07 $layer=LI1_cond $X=6.975 $Y=1.52
+ $X2=7.09 $Y2=1.52
r25 12 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=3.16
+ $X2=7.09 $Y2=3.245
r26 11 15 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.09 $Y=1.61 $X2=7.09
+ $Y2=1.52
r27 11 12 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=7.09 $Y=1.61
+ $X2=7.09 $Y2=3.16
r28 7 13 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.975 $Y=1.43 $X2=6.975
+ $Y2=1.52
r29 7 9 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.975 $Y=1.43
+ $X2=6.975 $Y2=0.825
r30 2 30 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.835
+ $Y=3.085 $X2=6.975 $Y2=5.835
r31 2 25 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.835
+ $Y=3.085 $X2=6.975 $Y2=3.455
r32 1 9 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.835
+ $Y=0.575 $X2=6.975 $Y2=0.825
.ends

