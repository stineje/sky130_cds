magic
tech sky130A
magscale 1 2
timestamp 1612371718
<< nwell >>
rect -9 529 374 1119
<< nmoslvt >>
rect 80 115 110 225
rect 152 115 182 225
rect 252 115 282 225
<< pmos >>
rect 80 713 110 965
rect 166 713 196 965
rect 252 713 282 965
<< ndiff >>
rect 27 199 80 225
rect 27 131 35 199
rect 69 131 80 199
rect 27 115 80 131
rect 110 115 152 225
rect 182 199 252 225
rect 182 131 193 199
rect 227 131 252 199
rect 182 115 252 131
rect 282 199 335 225
rect 282 131 293 199
rect 327 131 335 199
rect 282 115 335 131
<< pdiff >>
rect 27 949 80 965
rect 27 813 35 949
rect 69 813 80 949
rect 27 713 80 813
rect 110 949 166 965
rect 110 813 121 949
rect 155 813 166 949
rect 110 713 166 813
rect 196 949 252 965
rect 196 813 207 949
rect 241 813 252 949
rect 196 713 252 813
rect 282 949 335 965
rect 282 813 293 949
rect 327 813 335 949
rect 282 713 335 813
<< ndiffc >>
rect 35 131 69 199
rect 193 131 227 199
rect 293 131 327 199
<< pdiffc >>
rect 35 813 69 949
rect 121 813 155 949
rect 207 813 241 949
rect 293 813 327 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 991
rect 80 534 110 713
rect 27 518 110 534
rect 27 484 37 518
rect 71 484 110 518
rect 27 468 110 484
rect 80 225 110 468
rect 166 466 196 713
rect 252 540 282 713
rect 252 510 289 540
rect 152 450 217 466
rect 152 416 173 450
rect 207 416 217 450
rect 152 400 217 416
rect 152 225 182 400
rect 259 368 289 510
rect 259 352 313 368
rect 259 332 269 352
rect 252 318 269 332
rect 303 318 313 352
rect 252 302 313 318
rect 252 225 282 302
rect 80 89 110 115
rect 152 89 182 115
rect 252 89 282 115
<< polycont >>
rect 37 484 71 518
rect 173 416 207 450
rect 269 318 303 352
<< locali >>
rect 0 1089 374 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 374 1089
rect 35 949 69 1049
rect 121 949 155 965
rect 35 797 69 813
rect 105 813 121 831
rect 105 797 155 813
rect 207 949 241 1049
rect 207 797 241 813
rect 293 949 327 965
rect 37 518 71 597
rect 37 468 71 484
rect 105 352 139 797
rect 173 450 207 523
rect 293 483 327 813
rect 173 400 207 416
rect 35 318 269 352
rect 303 318 319 352
rect 35 199 69 318
rect 35 115 69 131
rect 193 199 227 215
rect 193 61 227 131
rect 293 199 327 227
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 37 597 71 631
rect 173 523 207 557
rect 293 449 327 483
rect 293 227 327 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 374 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 374 1089
rect 0 1049 374 1055
rect 25 631 83 637
rect 25 597 37 631
rect 71 597 105 631
rect 25 591 83 597
rect 161 557 219 563
rect 140 523 173 557
rect 207 523 219 557
rect 161 517 219 523
rect 281 483 339 489
rect 281 449 293 483
rect 327 449 339 483
rect 281 443 339 449
rect 293 267 327 443
rect 281 261 339 267
rect 281 227 293 261
rect 327 227 339 261
rect 281 221 339 227
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 311 392 311 392 1 Y
port 1 n
rlabel viali 55 614 55 614 1 A
port 2 n
rlabel viali 191 540 191 540 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
