* File: sky130_osu_sc_12T_ls__nand2_l.pxi.spice
* Created: Fri Nov 12 15:38:47 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__NAND2_L%GND N_GND_M1000_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_10_p GND N_GND_c_3_p PM_SKY130_OSU_SC_12T_LS__NAND2_L%GND
x_PM_SKY130_OSU_SC_12T_LS__NAND2_L%VDD N_VDD_M1001_s N_VDD_M1003_d N_VDD_M1001_b
+ N_VDD_c_26_p N_VDD_c_27_p N_VDD_c_36_p VDD N_VDD_c_28_p
+ PM_SKY130_OSU_SC_12T_LS__NAND2_L%VDD
x_PM_SKY130_OSU_SC_12T_LS__NAND2_L%A N_A_M1002_g N_A_M1001_g N_A_c_49_n
+ N_A_c_50_n A PM_SKY130_OSU_SC_12T_LS__NAND2_L%A
x_PM_SKY130_OSU_SC_12T_LS__NAND2_L%B N_B_M1000_g N_B_M1003_g N_B_c_82_n
+ N_B_c_83_n N_B_c_84_n B PM_SKY130_OSU_SC_12T_LS__NAND2_L%B
x_PM_SKY130_OSU_SC_12T_LS__NAND2_L%Y N_Y_M1002_s N_Y_M1001_d N_Y_c_114_n
+ N_Y_c_117_n N_Y_c_118_n N_Y_c_119_n Y N_Y_c_121_n
+ PM_SKY130_OSU_SC_12T_LS__NAND2_L%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.119782f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.755
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.755
cc_3 N_GND_c_3_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.755
cc_4 N_GND_M1002_b N_A_M1001_g 0.00327281f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.445
cc_5 N_GND_M1002_b N_A_c_49_n 0.0487757f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.575
cc_6 N_GND_M1002_b N_A_c_50_n 0.00717647f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.575
cc_7 N_GND_M1002_b A 0.00300043f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.85
cc_8 N_GND_M1002_b N_B_M1000_g 0.0661988f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.755
cc_9 N_GND_c_2_p N_B_M1000_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.755
cc_10 N_GND_c_10_p N_B_M1000_g 0.00502587f $X=1.05 $Y=0.74 $X2=0.835 $Y2=0.755
cc_11 N_GND_c_3_p N_B_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.755
cc_12 N_GND_M1002_b N_B_M1003_g 0.0497877f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.445
cc_13 N_GND_M1002_b N_B_c_82_n 0.0369336f $X=-0.045 $Y=0 $X2=0.915 $Y2=1.825
cc_14 N_GND_M1002_b N_B_c_83_n 0.0293783f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.85
cc_15 N_GND_M1002_b N_B_c_84_n 0.0123076f $X=-0.045 $Y=0 $X2=1.06 $Y2=1.825
cc_16 N_GND_M1002_b B 0.00489846f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.85
cc_17 N_GND_M1002_b N_Y_c_114_n 0.0259786f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.74
cc_18 N_GND_c_2_p N_Y_c_114_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26 $Y2=0.74
cc_19 N_GND_c_3_p N_Y_c_114_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26 $Y2=0.74
cc_20 N_GND_M1002_b N_Y_c_117_n 0.00852443f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.48
cc_21 N_GND_M1002_b N_Y_c_118_n 0.0101912f $X=-0.045 $Y=0 $X2=0.605 $Y2=1.37
cc_22 N_GND_M1002_b N_Y_c_119_n 0.0242516f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.37
cc_23 N_GND_M1002_b Y 0.0166407f $X=-0.045 $Y=0 $X2=0.68 $Y2=2.24
cc_24 N_GND_M1002_b N_Y_c_121_n 0.00524085f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.48
cc_25 N_VDD_M1001_b N_A_M1001_g 0.0263245f $X=-0.045 $Y=2.795 $X2=0.475
+ $Y2=3.445
cc_26 N_VDD_c_26_p N_A_M1001_g 0.00713292f $X=0.26 $Y=3.615 $X2=0.475 $Y2=3.445
cc_27 N_VDD_c_27_p N_A_M1001_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.445
cc_28 N_VDD_c_28_p N_A_M1001_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.445
cc_29 N_VDD_c_26_p N_A_c_49_n 0.00164789f $X=0.26 $Y=3.615 $X2=0.32 $Y2=2.575
cc_30 N_VDD_M1001_b N_A_c_50_n 0.0032924f $X=-0.045 $Y=2.795 $X2=0.32 $Y2=2.575
cc_31 N_VDD_c_26_p N_A_c_50_n 0.00297982f $X=0.26 $Y=3.615 $X2=0.32 $Y2=2.575
cc_32 N_VDD_M1001_b A 0.0117399f $X=-0.045 $Y=2.795 $X2=0.32 $Y2=2.85
cc_33 N_VDD_c_26_p A 0.00538653f $X=0.26 $Y=3.615 $X2=0.32 $Y2=2.85
cc_34 N_VDD_M1001_b N_B_M1003_g 0.0263245f $X=-0.045 $Y=2.795 $X2=0.905
+ $Y2=3.445
cc_35 N_VDD_c_27_p N_B_M1003_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.445
cc_36 N_VDD_c_36_p N_B_M1003_g 0.00713292f $X=1.12 $Y=3.615 $X2=0.905 $Y2=3.445
cc_37 N_VDD_c_28_p N_B_M1003_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.905 $Y2=3.445
cc_38 N_VDD_M1001_b N_B_c_83_n 0.00329491f $X=-0.045 $Y=2.795 $X2=1.06 $Y2=2.85
cc_39 N_VDD_c_36_p N_B_c_83_n 0.00299223f $X=1.12 $Y=3.615 $X2=1.06 $Y2=2.85
cc_40 N_VDD_M1001_b B 0.0117399f $X=-0.045 $Y=2.795 $X2=1.06 $Y2=2.85
cc_41 N_VDD_c_36_p B 0.00538653f $X=1.12 $Y=3.615 $X2=1.06 $Y2=2.85
cc_42 N_VDD_M1001_b N_Y_c_117_n 0.00553429f $X=-0.045 $Y=2.795 $X2=0.69 $Y2=2.48
cc_43 N_VDD_c_27_p N_Y_c_117_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69 $Y2=2.48
cc_44 N_VDD_c_28_p N_Y_c_117_n 0.00475776f $X=1.02 $Y=4.25 $X2=0.69 $Y2=2.48
cc_45 N_A_M1002_g N_B_M1000_g 0.0967758f $X=0.475 $Y=0.755 $X2=0.835 $Y2=0.755
cc_46 N_A_M1002_g N_B_M1003_g 0.0670829f $X=0.475 $Y=0.755 $X2=0.905 $Y2=3.445
cc_47 N_A_M1002_g N_B_c_83_n 0.00248145f $X=0.475 $Y=0.755 $X2=1.06 $Y2=2.85
cc_48 N_A_M1002_g N_B_c_84_n 0.00282768f $X=0.475 $Y=0.755 $X2=1.06 $Y2=1.825
cc_49 A B 0.0182713f $X=0.32 $Y=2.85 $X2=1.06 $Y2=2.85
cc_50 N_A_M1002_g N_Y_c_114_n 0.0190376f $X=0.475 $Y=0.755 $X2=0.26 $Y2=0.74
cc_51 N_A_M1002_g N_Y_c_117_n 0.00813643f $X=0.475 $Y=0.755 $X2=0.69 $Y2=2.48
cc_52 N_A_c_50_n N_Y_c_117_n 0.0288062f $X=0.32 $Y=2.575 $X2=0.69 $Y2=2.48
cc_53 A N_Y_c_117_n 0.00300775f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_54 N_A_M1002_g N_Y_c_118_n 0.0136921f $X=0.475 $Y=0.755 $X2=0.605 $Y2=1.37
cc_55 N_A_M1002_g N_Y_c_119_n 0.00393078f $X=0.475 $Y=0.755 $X2=0.405 $Y2=1.37
cc_56 N_A_M1002_g Y 0.0125133f $X=0.475 $Y=0.755 $X2=0.68 $Y2=2.24
cc_57 N_A_M1002_g N_Y_c_121_n 0.00216533f $X=0.475 $Y=0.755 $X2=0.69 $Y2=2.48
cc_58 N_A_c_49_n N_Y_c_121_n 0.00274987f $X=0.32 $Y=2.575 $X2=0.69 $Y2=2.48
cc_59 N_A_c_50_n N_Y_c_121_n 0.00474021f $X=0.32 $Y=2.575 $X2=0.69 $Y2=2.48
cc_60 A N_Y_c_121_n 0.00280435f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_61 N_B_M1003_g N_Y_c_117_n 0.00772009f $X=0.905 $Y=3.445 $X2=0.69 $Y2=2.48
cc_62 N_B_c_83_n N_Y_c_117_n 0.0295869f $X=1.06 $Y=2.85 $X2=0.69 $Y2=2.48
cc_63 N_B_c_84_n N_Y_c_117_n 5.24123e-19 $X=1.06 $Y=1.825 $X2=0.69 $Y2=2.48
cc_64 B N_Y_c_117_n 0.00301465f $X=1.06 $Y=2.85 $X2=0.69 $Y2=2.48
cc_65 N_B_M1000_g N_Y_c_118_n 0.00853825f $X=0.835 $Y=0.755 $X2=0.605 $Y2=1.37
cc_66 N_B_M1000_g Y 0.00770103f $X=0.835 $Y=0.755 $X2=0.68 $Y2=2.24
cc_67 N_B_M1003_g Y 0.00539744f $X=0.905 $Y=3.445 $X2=0.68 $Y2=2.24
cc_68 N_B_c_82_n Y 0.00401356f $X=0.915 $Y=1.825 $X2=0.68 $Y2=2.24
cc_69 N_B_c_83_n Y 0.0183986f $X=1.06 $Y=2.85 $X2=0.68 $Y2=2.24
cc_70 N_B_c_84_n Y 0.0141623f $X=1.06 $Y=1.825 $X2=0.68 $Y2=2.24
cc_71 N_B_M1003_g N_Y_c_121_n 0.00341272f $X=0.905 $Y=3.445 $X2=0.69 $Y2=2.48
cc_72 N_B_c_82_n N_Y_c_121_n 0.00144278f $X=0.915 $Y=1.825 $X2=0.69 $Y2=2.48
cc_73 N_B_c_83_n N_Y_c_121_n 0.00640429f $X=1.06 $Y=2.85 $X2=0.69 $Y2=2.48
cc_74 N_B_c_84_n N_Y_c_121_n 0.00194461f $X=1.06 $Y=1.825 $X2=0.69 $Y2=2.48
cc_75 B N_Y_c_121_n 0.00280435f $X=1.06 $Y=2.85 $X2=0.69 $Y2=2.48
