* File: sky130_osu_sc_12T_ms__dff_l.pxi.spice
* Created: Fri Nov 12 15:22:30 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%GND N_GND_M1004_d N_GND_M1011_d N_GND_M1023_d
+ N_GND_M1007_s N_GND_M1008_d N_GND_M1004_b N_GND_c_2_p N_GND_c_3_p N_GND_c_16_p
+ N_GND_c_59_p N_GND_c_35_p N_GND_c_39_p N_GND_c_40_p N_GND_c_41_p N_GND_c_116_p
+ N_GND_c_117_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_MS__DFF_L%GND
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%VDD N_VDD_M1019_d N_VDD_M1002_d N_VDD_M1014_d
+ N_VDD_M1021_s N_VDD_M1006_d N_VDD_M1019_b N_VDD_c_182_p N_VDD_c_183_p
+ N_VDD_c_192_p N_VDD_c_218_p N_VDD_c_203_p N_VDD_c_207_p N_VDD_c_208_p
+ N_VDD_c_209_p N_VDD_c_249_p N_VDD_c_250_p N_VDD_c_273_p VDD N_VDD_c_184_p
+ PM_SKY130_OSU_SC_12T_MS__DFF_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%A_75_248# N_A_75_248#_M1022_d
+ N_A_75_248#_M1013_d N_A_75_248#_M1004_g N_A_75_248#_M1019_g
+ N_A_75_248#_c_289_n N_A_75_248#_c_290_n N_A_75_248#_c_291_n
+ N_A_75_248#_c_307_n N_A_75_248#_c_292_n N_A_75_248#_c_294_n
+ N_A_75_248#_c_308_n N_A_75_248#_c_310_n N_A_75_248#_c_296_n
+ N_A_75_248#_c_312_n N_A_75_248#_c_297_n N_A_75_248#_c_298_n
+ N_A_75_248#_c_299_n PM_SKY130_OSU_SC_12T_MS__DFF_L%A_75_248#
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%D N_D_M1003_g N_D_M1018_g N_D_c_377_n
+ N_D_c_378_n D PM_SKY130_OSU_SC_12T_MS__DFF_L%D
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%CK N_CK_M1013_g N_CK_M1016_g N_CK_M1010_g
+ N_CK_M1017_g N_CK_M1024_g N_CK_c_415_n N_CK_M1015_g N_CK_c_416_n N_CK_c_417_n
+ N_CK_c_418_n N_CK_c_419_n N_CK_c_422_n N_CK_c_423_n N_CK_c_426_n N_CK_c_427_n
+ N_CK_c_432_n N_CK_c_433_n N_CK_c_434_n N_CK_c_435_n N_CK_c_436_n N_CK_c_437_n
+ N_CK_c_438_n N_CK_c_439_n N_CK_c_440_n N_CK_c_441_n N_CK_c_442_n N_CK_c_443_n
+ N_CK_c_444_n CK PM_SKY130_OSU_SC_12T_MS__DFF_L%CK
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%A_32_115# N_A_32_115#_M1004_s
+ N_A_32_115#_M1019_s N_A_32_115#_M1011_g N_A_32_115#_M1002_g
+ N_A_32_115#_c_649_n N_A_32_115#_c_651_n N_A_32_115#_c_652_n
+ N_A_32_115#_c_653_n N_A_32_115#_M1012_g N_A_32_115#_M1005_g
+ N_A_32_115#_c_658_n N_A_32_115#_c_659_n N_A_32_115#_c_680_n
+ N_A_32_115#_c_662_n N_A_32_115#_c_663_n N_A_32_115#_c_685_n
+ N_A_32_115#_c_664_n N_A_32_115#_c_666_n N_A_32_115#_c_668_n
+ N_A_32_115#_c_669_n PM_SKY130_OSU_SC_12T_MS__DFF_L%A_32_115#
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%A_243_89# N_A_243_89#_M1024_d
+ N_A_243_89#_M1015_d N_A_243_89#_c_759_n N_A_243_89#_M1022_g
+ N_A_243_89#_c_762_n N_A_243_89#_c_763_n N_A_243_89#_c_764_n
+ N_A_243_89#_M1009_g N_A_243_89#_c_766_n N_A_243_89#_M1000_g
+ N_A_243_89#_c_768_n N_A_243_89#_M1001_g N_A_243_89#_c_772_n
+ N_A_243_89#_c_773_n N_A_243_89#_c_774_n N_A_243_89#_c_775_n
+ N_A_243_89#_c_776_n N_A_243_89#_c_777_n N_A_243_89#_c_792_n
+ N_A_243_89#_c_781_n N_A_243_89#_c_782_n N_A_243_89#_c_797_n
+ N_A_243_89#_c_783_n N_A_243_89#_c_784_n N_A_243_89#_c_785_n
+ PM_SKY130_OSU_SC_12T_MS__DFF_L%A_243_89#
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%A_785_89# N_A_785_89#_M1007_d
+ N_A_785_89#_M1021_d N_A_785_89#_M1023_g N_A_785_89#_M1014_g
+ N_A_785_89#_c_955_n N_A_785_89#_M1008_g N_A_785_89#_M1006_g
+ N_A_785_89#_c_960_n N_A_785_89#_c_962_n N_A_785_89#_c_986_n
+ N_A_785_89#_c_963_n N_A_785_89#_c_964_n N_A_785_89#_c_965_n
+ N_A_785_89#_c_968_n N_A_785_89#_c_969_n N_A_785_89#_c_970_n
+ N_A_785_89#_c_971_n N_A_785_89#_c_972_n N_A_785_89#_c_973_n
+ N_A_785_89#_c_974_n N_A_785_89#_c_975_n N_A_785_89#_c_976_n
+ PM_SKY130_OSU_SC_12T_MS__DFF_L%A_785_89#
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%A_623_115# N_A_623_115#_M1010_d
+ N_A_623_115#_M1000_d N_A_623_115#_c_1116_n N_A_623_115#_M1007_g
+ N_A_623_115#_M1021_g N_A_623_115#_c_1121_n N_A_623_115#_c_1123_n
+ N_A_623_115#_c_1153_n N_A_623_115#_c_1183_n N_A_623_115#_c_1142_n
+ N_A_623_115#_c_1124_n N_A_623_115#_c_1125_n N_A_623_115#_c_1127_n
+ N_A_623_115#_c_1130_n N_A_623_115#_c_1131_n N_A_623_115#_c_1132_n
+ N_A_623_115#_c_1134_n N_A_623_115#_c_1135_n
+ PM_SKY130_OSU_SC_12T_MS__DFF_L%A_623_115#
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%ON N_ON_M1008_s N_ON_M1006_s N_ON_M1025_g
+ N_ON_M1020_g N_ON_c_1240_n N_ON_c_1241_n N_ON_c_1244_n N_ON_c_1245_n
+ N_ON_c_1246_n N_ON_c_1248_n N_ON_c_1249_n N_ON_c_1250_n N_ON_c_1251_n
+ N_ON_c_1252_n ON PM_SKY130_OSU_SC_12T_MS__DFF_L%ON
x_PM_SKY130_OSU_SC_12T_MS__DFF_L%Q N_Q_M1025_d N_Q_M1020_d N_Q_c_1317_n
+ N_Q_c_1323_n N_Q_c_1319_n N_Q_c_1320_n N_Q_c_1327_n N_Q_c_1328_n N_Q_c_1321_n
+ Q PM_SKY130_OSU_SC_12T_MS__DFF_L%Q
cc_1 N_GND_M1004_b N_A_75_248#_M1004_g 0.0223692f $X=-0.045 $Y=0 $X2=0.5
+ $Y2=0.835
cc_2 N_GND_c_2_p N_A_75_248#_M1004_g 0.00606474f $X=0.63 $Y=0.152 $X2=0.5
+ $Y2=0.835
cc_3 N_GND_c_3_p N_A_75_248#_M1004_g 0.00308284f $X=0.715 $Y=0.755 $X2=0.5
+ $Y2=0.835
cc_4 N_GND_c_4_p N_A_75_248#_M1004_g 0.00468827f $X=6.46 $Y=0.19 $X2=0.5
+ $Y2=0.835
cc_5 N_GND_M1004_b N_A_75_248#_c_289_n 0.0143449f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=1.39
cc_6 N_GND_M1004_b N_A_75_248#_c_290_n 0.0223136f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.285
cc_7 N_GND_M1004_b N_A_75_248#_c_291_n 0.0431517f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.12
cc_8 N_GND_M1004_b N_A_75_248#_c_292_n 0.0183015f $X=-0.045 $Y=0 $X2=1.405
+ $Y2=1.285
cc_9 N_GND_c_3_p N_A_75_248#_c_292_n 0.00456782f $X=0.715 $Y=0.755 $X2=1.405
+ $Y2=1.285
cc_10 N_GND_M1004_b N_A_75_248#_c_294_n 0.00315644f $X=-0.045 $Y=0 $X2=0.71
+ $Y2=1.285
cc_11 N_GND_c_3_p N_A_75_248#_c_294_n 0.00460441f $X=0.715 $Y=0.755 $X2=0.71
+ $Y2=1.285
cc_12 N_GND_M1004_b N_A_75_248#_c_296_n 0.00198494f $X=-0.045 $Y=0 $X2=1.49
+ $Y2=1.2
cc_13 N_GND_M1004_b N_A_75_248#_c_297_n 0.00325766f $X=-0.045 $Y=0 $X2=0.51
+ $Y2=2.285
cc_14 N_GND_M1004_b N_A_75_248#_c_298_n 0.0127034f $X=-0.045 $Y=0 $X2=0.567
+ $Y2=2.12
cc_15 N_GND_M1004_b N_A_75_248#_c_299_n 0.00311983f $X=-0.045 $Y=0 $X2=1.49
+ $Y2=0.755
cc_16 N_GND_c_16_p N_A_75_248#_c_299_n 0.0145844f $X=2.38 $Y=0.152 $X2=1.49
+ $Y2=0.755
cc_17 N_GND_c_4_p N_A_75_248#_c_299_n 0.0098977f $X=6.46 $Y=0.19 $X2=1.49
+ $Y2=0.755
cc_18 N_GND_M1004_b N_D_M1003_g 0.0334344f $X=-0.045 $Y=0 $X2=0.93 $Y2=0.835
cc_19 N_GND_c_3_p N_D_M1003_g 0.00308284f $X=0.715 $Y=0.755 $X2=0.93 $Y2=0.835
cc_20 N_GND_c_16_p N_D_M1003_g 0.00606474f $X=2.38 $Y=0.152 $X2=0.93 $Y2=0.835
cc_21 N_GND_c_4_p N_D_M1003_g 0.00468827f $X=6.46 $Y=0.19 $X2=0.93 $Y2=0.835
cc_22 N_GND_M1004_b N_D_M1018_g 0.0299924f $X=-0.045 $Y=0 $X2=0.93 $Y2=3.235
cc_23 N_GND_M1004_b N_D_c_377_n 0.0272793f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.74
cc_24 N_GND_M1004_b N_D_c_378_n 0.00311208f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.74
cc_25 N_GND_M1004_b D 0.00874398f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.74
cc_26 N_GND_M1004_b N_CK_c_415_n 0.0307453f $X=-0.045 $Y=0 $X2=4.43 $Y2=2.45
cc_27 N_GND_M1004_b N_CK_c_416_n 0.0445582f $X=-0.045 $Y=0 $X2=4.485 $Y2=2.12
cc_28 N_GND_M1004_b N_CK_c_417_n 0.0244054f $X=-0.045 $Y=0 $X2=1.35 $Y2=2.285
cc_29 N_GND_M1004_b N_CK_c_418_n 0.0254608f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.37
cc_30 N_GND_M1004_b N_CK_c_419_n 0.0173906f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.205
cc_31 N_GND_c_16_p N_CK_c_419_n 0.00606474f $X=2.38 $Y=0.152 $X2=1.83 $Y2=1.205
cc_32 N_GND_c_4_p N_CK_c_419_n 0.00468827f $X=6.46 $Y=0.19 $X2=1.83 $Y2=1.205
cc_33 N_GND_M1004_b N_CK_c_422_n 0.0268189f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.37
cc_34 N_GND_M1004_b N_CK_c_423_n 0.0174883f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.205
cc_35 N_GND_c_35_p N_CK_c_423_n 0.00606474f $X=4.13 $Y=0.152 $X2=3.1 $Y2=1.205
cc_36 N_GND_c_4_p N_CK_c_423_n 0.00468827f $X=6.46 $Y=0.19 $X2=3.1 $Y2=1.205
cc_37 N_GND_M1004_b N_CK_c_426_n 0.0218864f $X=-0.045 $Y=0 $X2=3.58 $Y2=2.285
cc_38 N_GND_M1004_b N_CK_c_427_n 0.0183851f $X=-0.045 $Y=0 $X2=4.457 $Y2=1.205
cc_39 N_GND_c_39_p N_CK_c_427_n 0.00308284f $X=4.215 $Y=0.755 $X2=4.457
+ $Y2=1.205
cc_40 N_GND_c_40_p N_CK_c_427_n 0.00606474f $X=5.08 $Y=0.152 $X2=4.457 $Y2=1.205
cc_41 N_GND_c_41_p N_CK_c_427_n 0.00365683f $X=5.165 $Y=0.755 $X2=4.457
+ $Y2=1.205
cc_42 N_GND_c_4_p N_CK_c_427_n 0.00468827f $X=6.46 $Y=0.19 $X2=4.457 $Y2=1.205
cc_43 N_GND_M1004_b N_CK_c_432_n 0.0141068f $X=-0.045 $Y=0 $X2=4.457 $Y2=1.355
cc_44 N_GND_M1004_b N_CK_c_433_n 0.00600607f $X=-0.045 $Y=0 $X2=1.745 $Y2=2.11
cc_45 N_GND_M1004_b N_CK_c_434_n 0.0107953f $X=-0.045 $Y=0 $X2=1.83 $Y2=1.37
cc_46 N_GND_M1004_b N_CK_c_435_n 0.00936067f $X=-0.045 $Y=0 $X2=3.1 $Y2=1.37
cc_47 N_GND_M1004_b N_CK_c_436_n 0.00482391f $X=-0.045 $Y=0 $X2=3.495 $Y2=2.11
cc_48 N_GND_M1004_b N_CK_c_437_n 5.00459e-19 $X=-0.045 $Y=0 $X2=3.185 $Y2=2.11
cc_49 N_GND_M1004_b N_CK_c_438_n 7.11312e-19 $X=-0.045 $Y=0 $X2=4.575 $Y2=2.11
cc_50 N_GND_M1004_b N_CK_c_439_n 0.00235115f $X=-0.045 $Y=0 $X2=1.35 $Y2=2.11
cc_51 N_GND_M1004_b N_CK_c_440_n 0.00120157f $X=-0.045 $Y=0 $X2=3.58 $Y2=2.11
cc_52 N_GND_M1004_b N_CK_c_441_n 0.0338553f $X=-0.045 $Y=0 $X2=3.435 $Y2=2.11
cc_53 N_GND_M1004_b N_CK_c_442_n 0.00614962f $X=-0.045 $Y=0 $X2=1.495 $Y2=2.11
cc_54 N_GND_M1004_b N_CK_c_443_n 0.013468f $X=-0.045 $Y=0 $X2=4.43 $Y2=2.11
cc_55 N_GND_M1004_b N_CK_c_444_n 0.00256396f $X=-0.045 $Y=0 $X2=3.725 $Y2=2.11
cc_56 N_GND_M1004_b CK 0.00144547f $X=-0.045 $Y=0 $X2=4.575 $Y2=2.11
cc_57 N_GND_M1004_b N_A_32_115#_M1011_g 0.0171926f $X=-0.045 $Y=0 $X2=2.25
+ $Y2=0.835
cc_58 N_GND_c_16_p N_A_32_115#_M1011_g 0.00606474f $X=2.38 $Y=0.152 $X2=2.25
+ $Y2=0.835
cc_59 N_GND_c_59_p N_A_32_115#_M1011_g 0.00308284f $X=2.465 $Y=0.74 $X2=2.25
+ $Y2=0.835
cc_60 N_GND_c_4_p N_A_32_115#_M1011_g 0.00468827f $X=6.46 $Y=0.19 $X2=2.25
+ $Y2=0.835
cc_61 N_GND_M1004_b N_A_32_115#_c_649_n 0.0241855f $X=-0.045 $Y=0 $X2=2.605
+ $Y2=1.37
cc_62 N_GND_c_59_p N_A_32_115#_c_649_n 9.93645e-19 $X=2.465 $Y=0.74 $X2=2.605
+ $Y2=1.37
cc_63 N_GND_M1004_b N_A_32_115#_c_651_n 0.0105855f $X=-0.045 $Y=0 $X2=2.325
+ $Y2=1.37
cc_64 N_GND_M1004_b N_A_32_115#_c_652_n 0.0232417f $X=-0.045 $Y=0 $X2=2.605
+ $Y2=2.285
cc_65 N_GND_M1004_b N_A_32_115#_c_653_n 0.0105265f $X=-0.045 $Y=0 $X2=2.325
+ $Y2=2.285
cc_66 N_GND_M1004_b N_A_32_115#_M1012_g 0.0171936f $X=-0.045 $Y=0 $X2=2.68
+ $Y2=0.835
cc_67 N_GND_c_59_p N_A_32_115#_M1012_g 0.00308284f $X=2.465 $Y=0.74 $X2=2.68
+ $Y2=0.835
cc_68 N_GND_c_35_p N_A_32_115#_M1012_g 0.00606474f $X=4.13 $Y=0.152 $X2=2.68
+ $Y2=0.835
cc_69 N_GND_c_4_p N_A_32_115#_M1012_g 0.00468827f $X=6.46 $Y=0.19 $X2=2.68
+ $Y2=0.835
cc_70 N_GND_M1004_b N_A_32_115#_c_658_n 0.0456538f $X=-0.045 $Y=0 $X2=0.17
+ $Y2=2.695
cc_71 N_GND_M1004_b N_A_32_115#_c_659_n 0.00613129f $X=-0.045 $Y=0 $X2=0.285
+ $Y2=0.755
cc_72 N_GND_c_2_p N_A_32_115#_c_659_n 0.00729833f $X=0.63 $Y=0.152 $X2=0.285
+ $Y2=0.755
cc_73 N_GND_c_4_p N_A_32_115#_c_659_n 0.00474439f $X=6.46 $Y=0.19 $X2=0.285
+ $Y2=0.755
cc_74 N_GND_M1004_b N_A_32_115#_c_662_n 0.00871176f $X=-0.045 $Y=0 $X2=2.42
+ $Y2=2.285
cc_75 N_GND_M1004_b N_A_32_115#_c_663_n 0.0203007f $X=-0.045 $Y=0 $X2=0.285
+ $Y2=1.37
cc_76 N_GND_M1004_b N_A_32_115#_c_664_n 0.00381957f $X=-0.045 $Y=0 $X2=2.42
+ $Y2=1.37
cc_77 N_GND_c_59_p N_A_32_115#_c_664_n 0.00673193f $X=2.465 $Y=0.74 $X2=2.42
+ $Y2=1.37
cc_78 N_GND_M1004_b N_A_32_115#_c_666_n 0.0225319f $X=-0.045 $Y=0 $X2=2.185
+ $Y2=1.37
cc_79 N_GND_c_3_p N_A_32_115#_c_666_n 0.00118122f $X=0.715 $Y=0.755 $X2=2.185
+ $Y2=1.37
cc_80 N_GND_M1004_b N_A_32_115#_c_668_n 0.00468924f $X=-0.045 $Y=0 $X2=0.43
+ $Y2=1.37
cc_81 N_GND_c_59_p N_A_32_115#_c_669_n 7.02397e-19 $X=2.465 $Y=0.74 $X2=2.33
+ $Y2=1.37
cc_82 N_GND_M1004_b N_A_243_89#_c_759_n 0.0173059f $X=-0.045 $Y=0 $X2=1.29
+ $Y2=1.205
cc_83 N_GND_c_16_p N_A_243_89#_c_759_n 0.00606474f $X=2.38 $Y=0.152 $X2=1.29
+ $Y2=1.205
cc_84 N_GND_c_4_p N_A_243_89#_c_759_n 0.00468827f $X=6.46 $Y=0.19 $X2=1.29
+ $Y2=1.205
cc_85 N_GND_M1004_b N_A_243_89#_c_762_n 0.0202867f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.745
cc_86 N_GND_M1004_b N_A_243_89#_c_763_n 0.0207095f $X=-0.045 $Y=0 $X2=1.815
+ $Y2=1.82
cc_87 N_GND_M1004_b N_A_243_89#_c_764_n 0.00755029f $X=-0.045 $Y=0 $X2=1.485
+ $Y2=1.82
cc_88 N_GND_M1004_b N_A_243_89#_M1009_g 0.032457f $X=-0.045 $Y=0 $X2=1.89
+ $Y2=3.235
cc_89 N_GND_M1004_b N_A_243_89#_c_766_n 0.0559794f $X=-0.045 $Y=0 $X2=2.965
+ $Y2=1.82
cc_90 N_GND_M1004_b N_A_243_89#_M1000_g 0.0313037f $X=-0.045 $Y=0 $X2=3.04
+ $Y2=3.235
cc_91 N_GND_M1004_b N_A_243_89#_c_768_n 0.0211051f $X=-0.045 $Y=0 $X2=3.445
+ $Y2=1.825
cc_92 N_GND_M1004_b N_A_243_89#_M1001_g 0.035333f $X=-0.045 $Y=0 $X2=3.64
+ $Y2=0.835
cc_93 N_GND_c_35_p N_A_243_89#_M1001_g 0.00606474f $X=4.13 $Y=0.152 $X2=3.64
+ $Y2=0.835
cc_94 N_GND_c_4_p N_A_243_89#_M1001_g 0.00468827f $X=6.46 $Y=0.19 $X2=3.64
+ $Y2=0.835
cc_95 N_GND_M1004_b N_A_243_89#_c_772_n 0.0141736f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.28
cc_96 N_GND_M1004_b N_A_243_89#_c_773_n 0.00426512f $X=-0.045 $Y=0 $X2=1.89
+ $Y2=1.82
cc_97 N_GND_M1004_b N_A_243_89#_c_774_n 0.00467948f $X=-0.045 $Y=0 $X2=3.04
+ $Y2=1.825
cc_98 N_GND_M1004_b N_A_243_89#_c_775_n 0.0262245f $X=-0.045 $Y=0 $X2=3.58
+ $Y2=1.74
cc_99 N_GND_M1004_b N_A_243_89#_c_776_n 0.00205129f $X=-0.045 $Y=0 $X2=3.58
+ $Y2=1.74
cc_100 N_GND_M1004_b N_A_243_89#_c_777_n 0.0151485f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=0.755
cc_101 N_GND_c_40_p N_A_243_89#_c_777_n 0.00749582f $X=5.08 $Y=0.152 $X2=4.645
+ $Y2=0.755
cc_102 N_GND_c_41_p N_A_243_89#_c_777_n 0.0153786f $X=5.165 $Y=0.755 $X2=4.645
+ $Y2=0.755
cc_103 N_GND_c_4_p N_A_243_89#_c_777_n 0.00476261f $X=6.46 $Y=0.19 $X2=4.645
+ $Y2=0.755
cc_104 N_GND_M1004_b N_A_243_89#_c_781_n 0.0123446f $X=-0.045 $Y=0 $X2=4.915
+ $Y2=2.62
cc_105 N_GND_M1004_b N_A_243_89#_c_782_n 0.011016f $X=-0.045 $Y=0 $X2=4.915
+ $Y2=1.725
cc_106 N_GND_M1004_b N_A_243_89#_c_783_n 0.00174422f $X=-0.045 $Y=0 $X2=3.725
+ $Y2=1.725
cc_107 N_GND_M1004_b N_A_243_89#_c_784_n 0.00217465f $X=-0.045 $Y=0 $X2=4.645
+ $Y2=1.74
cc_108 N_GND_M1004_b N_A_243_89#_c_785_n 0.00682657f $X=-0.045 $Y=0 $X2=4.5
+ $Y2=1.74
cc_109 N_GND_M1004_b N_A_785_89#_M1023_g 0.0337299f $X=-0.045 $Y=0 $X2=4
+ $Y2=0.835
cc_110 N_GND_c_35_p N_A_785_89#_M1023_g 0.00606474f $X=4.13 $Y=0.152 $X2=4
+ $Y2=0.835
cc_111 N_GND_c_39_p N_A_785_89#_M1023_g 0.00308284f $X=4.215 $Y=0.755 $X2=4
+ $Y2=0.835
cc_112 N_GND_c_4_p N_A_785_89#_M1023_g 0.00468827f $X=6.46 $Y=0.19 $X2=4
+ $Y2=0.835
cc_113 N_GND_M1004_b N_A_785_89#_M1014_g 0.0286123f $X=-0.045 $Y=0 $X2=4
+ $Y2=3.235
cc_114 N_GND_M1004_b N_A_785_89#_c_955_n 0.0524798f $X=-0.045 $Y=0 $X2=6.28
+ $Y2=1.905
cc_115 N_GND_M1004_b N_A_785_89#_M1008_g 0.0332752f $X=-0.045 $Y=0 $X2=6.33
+ $Y2=0.755
cc_116 N_GND_c_116_p N_A_785_89#_M1008_g 0.00606474f $X=6.46 $Y=0.152 $X2=6.33
+ $Y2=0.755
cc_117 N_GND_c_117_p N_A_785_89#_M1008_g 0.00308284f $X=6.545 $Y=0.74 $X2=6.33
+ $Y2=0.755
cc_118 N_GND_c_4_p N_A_785_89#_M1008_g 0.00468827f $X=6.46 $Y=0.19 $X2=6.33
+ $Y2=0.755
cc_119 N_GND_M1004_b N_A_785_89#_c_960_n 0.0262718f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=1.74
cc_120 N_GND_c_39_p N_A_785_89#_c_960_n 0.00144867f $X=4.215 $Y=0.755 $X2=4.06
+ $Y2=1.74
cc_121 N_GND_M1004_b N_A_785_89#_c_962_n 0.0304692f $X=-0.045 $Y=0 $X2=6.305
+ $Y2=2.475
cc_122 N_GND_M1004_b N_A_785_89#_c_963_n 8.68018e-19 $X=-0.045 $Y=0 $X2=4.062
+ $Y2=1.812
cc_123 N_GND_M1004_b N_A_785_89#_c_964_n 0.00374026f $X=-0.045 $Y=0 $X2=4.06
+ $Y2=2.48
cc_124 N_GND_M1004_b N_A_785_89#_c_965_n 0.0143842f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=0.755
cc_125 N_GND_c_116_p N_A_785_89#_c_965_n 0.0074445f $X=6.46 $Y=0.152 $X2=5.595
+ $Y2=0.755
cc_126 N_GND_c_4_p N_A_785_89#_c_965_n 0.00476261f $X=6.46 $Y=0.19 $X2=5.595
+ $Y2=0.755
cc_127 N_GND_M1004_b N_A_785_89#_c_968_n 0.013534f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=2.955
cc_128 N_GND_M1004_b N_A_785_89#_c_969_n 0.0122098f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=1.74
cc_129 N_GND_M1004_b N_A_785_89#_c_970_n 0.00242672f $X=-0.045 $Y=0 $X2=5.595
+ $Y2=1.74
cc_130 N_GND_M1004_b N_A_785_89#_c_971_n 0.00262889f $X=-0.045 $Y=0 $X2=4.935
+ $Y2=2.48
cc_131 N_GND_M1004_b N_A_785_89#_c_972_n 0.00120404f $X=-0.045 $Y=0 $X2=4.205
+ $Y2=2.48
cc_132 N_GND_M1004_b N_A_785_89#_c_973_n 0.0053881f $X=-0.045 $Y=0 $X2=5.007
+ $Y2=2.395
cc_133 N_GND_M1004_b N_A_785_89#_c_974_n 0.0342266f $X=-0.045 $Y=0 $X2=6.08
+ $Y2=1.74
cc_134 N_GND_M1004_b N_A_785_89#_c_975_n 3.47949e-19 $X=-0.045 $Y=0 $X2=5.08
+ $Y2=1.74
cc_135 N_GND_M1004_b N_A_785_89#_c_976_n 0.00114171f $X=-0.045 $Y=0 $X2=6.215
+ $Y2=1.74
cc_136 N_GND_M1004_b N_A_623_115#_c_1116_n 0.0221119f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=1.205
cc_137 N_GND_c_41_p N_A_623_115#_c_1116_n 0.00502587f $X=5.165 $Y=0.755 $X2=5.38
+ $Y2=1.205
cc_138 N_GND_c_116_p N_A_623_115#_c_1116_n 0.00606474f $X=6.46 $Y=0.152 $X2=5.38
+ $Y2=1.205
cc_139 N_GND_c_4_p N_A_623_115#_c_1116_n 0.00468827f $X=6.46 $Y=0.19 $X2=5.38
+ $Y2=1.205
cc_140 N_GND_M1004_b N_A_623_115#_M1021_g 0.0594603f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=3.235
cc_141 N_GND_M1004_b N_A_623_115#_c_1121_n 0.0482869f $X=-0.045 $Y=0 $X2=5.38
+ $Y2=1.37
cc_142 N_GND_c_41_p N_A_623_115#_c_1121_n 0.00386381f $X=5.165 $Y=0.755 $X2=5.38
+ $Y2=1.37
cc_143 N_GND_M1004_b N_A_623_115#_c_1123_n 0.0110483f $X=-0.045 $Y=0 $X2=2.76
+ $Y2=1.37
cc_144 N_GND_M1004_b N_A_623_115#_c_1124_n 0.00919317f $X=-0.045 $Y=0 $X2=3.44
+ $Y2=1.34
cc_145 N_GND_M1004_b N_A_623_115#_c_1125_n 0.00162209f $X=-0.045 $Y=0 $X2=5.175
+ $Y2=1.37
cc_146 N_GND_c_41_p N_A_623_115#_c_1125_n 0.00509685f $X=5.165 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_147 N_GND_M1004_b N_A_623_115#_c_1127_n 0.00312748f $X=-0.045 $Y=0 $X2=3.34
+ $Y2=0.755
cc_148 N_GND_c_35_p N_A_623_115#_c_1127_n 0.0152394f $X=4.13 $Y=0.152 $X2=3.34
+ $Y2=0.755
cc_149 N_GND_c_4_p N_A_623_115#_c_1127_n 0.00994746f $X=6.46 $Y=0.19 $X2=3.34
+ $Y2=0.755
cc_150 N_GND_M1004_b N_A_623_115#_c_1130_n 0.00411356f $X=-0.045 $Y=0 $X2=3.295
+ $Y2=1.37
cc_151 N_GND_M1004_b N_A_623_115#_c_1131_n 0.00645173f $X=-0.045 $Y=0 $X2=2.905
+ $Y2=1.37
cc_152 N_GND_M1004_b N_A_623_115#_c_1132_n 0.0299969f $X=-0.045 $Y=0 $X2=5.03
+ $Y2=1.37
cc_153 N_GND_c_39_p N_A_623_115#_c_1132_n 0.00727398f $X=4.215 $Y=0.755 $X2=5.03
+ $Y2=1.37
cc_154 N_GND_M1004_b N_A_623_115#_c_1134_n 0.00466179f $X=-0.045 $Y=0 $X2=3.585
+ $Y2=1.37
cc_155 N_GND_M1004_b N_A_623_115#_c_1135_n 9.68419e-19 $X=-0.045 $Y=0 $X2=5.175
+ $Y2=1.37
cc_156 N_GND_c_41_p N_A_623_115#_c_1135_n 0.00387325f $X=5.165 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_157 N_GND_M1004_b N_ON_M1025_g 0.0703925f $X=-0.045 $Y=0 $X2=6.76 $Y2=0.755
cc_158 N_GND_c_117_p N_ON_M1025_g 0.00308284f $X=6.545 $Y=0.74 $X2=6.76
+ $Y2=0.755
cc_159 N_GND_c_4_p N_ON_M1025_g 0.00468827f $X=6.46 $Y=0.19 $X2=6.76 $Y2=0.755
cc_160 N_GND_M1004_b N_ON_M1020_g 0.0150123f $X=-0.045 $Y=0 $X2=6.76 $Y2=3.445
cc_161 N_GND_M1004_b N_ON_c_1240_n 0.0285256f $X=-0.045 $Y=0 $X2=6.7 $Y2=2.015
cc_162 N_GND_M1004_b N_ON_c_1241_n 0.00988245f $X=-0.045 $Y=0 $X2=6.115 $Y2=0.74
cc_163 N_GND_c_116_p N_ON_c_1241_n 0.00757793f $X=6.46 $Y=0.152 $X2=6.115
+ $Y2=0.74
cc_164 N_GND_c_4_p N_ON_c_1241_n 0.00476261f $X=6.46 $Y=0.19 $X2=6.115 $Y2=0.74
cc_165 N_GND_M1004_b N_ON_c_1244_n 0.00173247f $X=-0.045 $Y=0 $X2=6.115
+ $Y2=2.195
cc_166 N_GND_M1004_b N_ON_c_1245_n 0.00445021f $X=-0.045 $Y=0 $X2=6.115
+ $Y2=3.615
cc_167 N_GND_M1004_b N_ON_c_1246_n 0.00951514f $X=-0.045 $Y=0 $X2=6.615 $Y2=1.4
cc_168 N_GND_c_117_p N_ON_c_1246_n 0.00738334f $X=6.545 $Y=0.74 $X2=6.615
+ $Y2=1.4
cc_169 N_GND_M1004_b N_ON_c_1248_n 0.0026304f $X=-0.045 $Y=0 $X2=6.2 $Y2=1.4
cc_170 N_GND_M1004_b N_ON_c_1249_n 0.0131198f $X=-0.045 $Y=0 $X2=6.615 $Y2=2.11
cc_171 N_GND_M1004_b N_ON_c_1250_n 0.00154829f $X=-0.045 $Y=0 $X2=6.702
+ $Y2=1.658
cc_172 N_GND_M1004_b N_ON_c_1251_n 5.47532e-19 $X=-0.045 $Y=0 $X2=6.7 $Y2=2.015
cc_173 N_GND_M1004_b N_ON_c_1252_n 5.06249e-19 $X=-0.045 $Y=0 $X2=6.702
+ $Y2=1.745
cc_174 N_GND_M1004_b ON 0.00962953f $X=-0.045 $Y=0 $X2=6.115 $Y2=2.11
cc_175 N_GND_M1004_b N_Q_c_1317_n 0.0118075f $X=-0.045 $Y=0 $X2=6.975 $Y2=0.74
cc_176 N_GND_c_4_p N_Q_c_1317_n 0.00468662f $X=6.46 $Y=0.19 $X2=6.975 $Y2=0.74
cc_177 N_GND_M1004_b N_Q_c_1319_n 0.060171f $X=-0.045 $Y=0 $X2=7.09 $Y2=2.395
cc_178 N_GND_M1004_b N_Q_c_1320_n 0.00345218f $X=-0.045 $Y=0 $X2=7.09 $Y2=2.48
cc_179 N_GND_M1004_b N_Q_c_1321_n 0.0184257f $X=-0.045 $Y=0 $X2=7.09 $Y2=1.07
cc_180 N_GND_M1004_b Q 0.00636397f $X=-0.045 $Y=0 $X2=6.97 $Y2=2.48
cc_181 N_VDD_M1019_b N_A_75_248#_M1019_g 0.0224266f $X=-0.045 $Y=2.425 $X2=0.5
+ $Y2=3.235
cc_182 N_VDD_c_182_p N_A_75_248#_M1019_g 0.00606474f $X=0.63 $Y=4.287 $X2=0.5
+ $Y2=3.235
cc_183 N_VDD_c_183_p N_A_75_248#_M1019_g 0.00337744f $X=0.715 $Y=3.295 $X2=0.5
+ $Y2=3.235
cc_184 N_VDD_c_184_p N_A_75_248#_M1019_g 0.00468827f $X=6.46 $Y=4.25 $X2=0.5
+ $Y2=3.235
cc_185 N_VDD_M1019_b N_A_75_248#_c_290_n 0.00631278f $X=-0.045 $Y=2.425 $X2=0.51
+ $Y2=2.285
cc_186 N_VDD_M1019_b N_A_75_248#_c_307_n 0.00145465f $X=-0.045 $Y=2.425
+ $X2=0.625 $Y2=2.62
cc_187 N_VDD_M1019_d N_A_75_248#_c_308_n 0.00447048f $X=0.575 $Y=2.605 $X2=1.42
+ $Y2=2.705
cc_188 N_VDD_c_183_p N_A_75_248#_c_308_n 0.00499116f $X=0.715 $Y=3.295 $X2=1.42
+ $Y2=2.705
cc_189 N_VDD_M1019_d N_A_75_248#_c_310_n 0.00106276f $X=0.575 $Y=2.605 $X2=0.71
+ $Y2=2.705
cc_190 N_VDD_c_183_p N_A_75_248#_c_310_n 0.00488762f $X=0.715 $Y=3.295 $X2=0.71
+ $Y2=2.705
cc_191 N_VDD_M1019_b N_A_75_248#_c_312_n 0.00313975f $X=-0.045 $Y=2.425 $X2=1.59
+ $Y2=2.955
cc_192 N_VDD_c_192_p N_A_75_248#_c_312_n 0.0149076f $X=2.38 $Y=4.287 $X2=1.59
+ $Y2=2.955
cc_193 N_VDD_c_184_p N_A_75_248#_c_312_n 0.00958198f $X=6.46 $Y=4.25 $X2=1.59
+ $Y2=2.955
cc_194 N_VDD_M1019_b N_A_75_248#_c_297_n 2.30281e-19 $X=-0.045 $Y=2.425 $X2=0.51
+ $Y2=2.285
cc_195 N_VDD_M1019_b N_D_M1018_g 0.0196478f $X=-0.045 $Y=2.425 $X2=0.93
+ $Y2=3.235
cc_196 N_VDD_c_183_p N_D_M1018_g 0.00337744f $X=0.715 $Y=3.295 $X2=0.93
+ $Y2=3.235
cc_197 N_VDD_c_192_p N_D_M1018_g 0.00606474f $X=2.38 $Y=4.287 $X2=0.93 $Y2=3.235
cc_198 N_VDD_c_184_p N_D_M1018_g 0.00468827f $X=6.46 $Y=4.25 $X2=0.93 $Y2=3.235
cc_199 N_VDD_M1019_b N_CK_M1013_g 0.0201249f $X=-0.045 $Y=2.425 $X2=1.29
+ $Y2=3.235
cc_200 N_VDD_c_192_p N_CK_M1013_g 0.00606474f $X=2.38 $Y=4.287 $X2=1.29
+ $Y2=3.235
cc_201 N_VDD_c_184_p N_CK_M1013_g 0.00468827f $X=6.46 $Y=4.25 $X2=1.29 $Y2=3.235
cc_202 N_VDD_M1019_b N_CK_M1017_g 0.0201163f $X=-0.045 $Y=2.425 $X2=3.64
+ $Y2=3.235
cc_203 N_VDD_c_203_p N_CK_M1017_g 0.00606474f $X=4.13 $Y=4.287 $X2=3.64
+ $Y2=3.235
cc_204 N_VDD_c_184_p N_CK_M1017_g 0.00468827f $X=6.46 $Y=4.25 $X2=3.64 $Y2=3.235
cc_205 N_VDD_M1019_b N_CK_c_415_n 0.007968f $X=-0.045 $Y=2.425 $X2=4.43 $Y2=2.45
cc_206 N_VDD_M1019_b N_CK_M1015_g 0.0218804f $X=-0.045 $Y=2.425 $X2=4.43
+ $Y2=3.235
cc_207 N_VDD_c_207_p N_CK_M1015_g 0.0047242f $X=4.215 $Y=3.21 $X2=4.43 $Y2=3.235
cc_208 N_VDD_c_208_p N_CK_M1015_g 0.00606474f $X=5.08 $Y=4.287 $X2=4.43
+ $Y2=3.235
cc_209 N_VDD_c_209_p N_CK_M1015_g 0.00455736f $X=5.165 $Y=3.295 $X2=4.43
+ $Y2=3.235
cc_210 N_VDD_c_184_p N_CK_M1015_g 0.00468827f $X=6.46 $Y=4.25 $X2=4.43 $Y2=3.235
cc_211 N_VDD_M1019_b N_CK_c_417_n 0.00487085f $X=-0.045 $Y=2.425 $X2=1.35
+ $Y2=2.285
cc_212 N_VDD_M1019_b N_CK_c_426_n 0.00486793f $X=-0.045 $Y=2.425 $X2=3.58
+ $Y2=2.285
cc_213 N_VDD_M1019_b N_CK_c_438_n 0.0010436f $X=-0.045 $Y=2.425 $X2=4.575
+ $Y2=2.11
cc_214 N_VDD_M1019_b N_CK_c_439_n 6.42499e-19 $X=-0.045 $Y=2.425 $X2=1.35
+ $Y2=2.11
cc_215 N_VDD_M1019_b N_CK_c_440_n 0.0022456f $X=-0.045 $Y=2.425 $X2=3.58
+ $Y2=2.11
cc_216 N_VDD_M1019_b N_A_32_115#_M1002_g 0.0192219f $X=-0.045 $Y=2.425 $X2=2.25
+ $Y2=3.235
cc_217 N_VDD_c_192_p N_A_32_115#_M1002_g 0.00606474f $X=2.38 $Y=4.287 $X2=2.25
+ $Y2=3.235
cc_218 N_VDD_c_218_p N_A_32_115#_M1002_g 0.00337744f $X=2.465 $Y=3.295 $X2=2.25
+ $Y2=3.235
cc_219 N_VDD_c_184_p N_A_32_115#_M1002_g 0.00468827f $X=6.46 $Y=4.25 $X2=2.25
+ $Y2=3.235
cc_220 N_VDD_c_218_p N_A_32_115#_c_652_n 8.24975e-19 $X=2.465 $Y=3.295 $X2=2.605
+ $Y2=2.285
cc_221 N_VDD_M1019_b N_A_32_115#_M1005_g 0.0181098f $X=-0.045 $Y=2.425 $X2=2.68
+ $Y2=3.235
cc_222 N_VDD_c_218_p N_A_32_115#_M1005_g 0.00337744f $X=2.465 $Y=3.295 $X2=2.68
+ $Y2=3.235
cc_223 N_VDD_c_203_p N_A_32_115#_M1005_g 0.00606474f $X=4.13 $Y=4.287 $X2=2.68
+ $Y2=3.235
cc_224 N_VDD_c_184_p N_A_32_115#_M1005_g 0.00468827f $X=6.46 $Y=4.25 $X2=2.68
+ $Y2=3.235
cc_225 N_VDD_M1019_b N_A_32_115#_c_658_n 0.0120505f $X=-0.045 $Y=2.425 $X2=0.17
+ $Y2=2.695
cc_226 N_VDD_M1019_b N_A_32_115#_c_680_n 0.00156053f $X=-0.045 $Y=2.425
+ $X2=0.285 $Y2=2.955
cc_227 N_VDD_c_182_p N_A_32_115#_c_680_n 0.00736239f $X=0.63 $Y=4.287 $X2=0.285
+ $Y2=2.955
cc_228 N_VDD_c_184_p N_A_32_115#_c_680_n 0.00476261f $X=6.46 $Y=4.25 $X2=0.285
+ $Y2=2.955
cc_229 N_VDD_M1019_b N_A_32_115#_c_662_n 0.00424346f $X=-0.045 $Y=2.425 $X2=2.42
+ $Y2=2.285
cc_230 N_VDD_c_218_p N_A_32_115#_c_662_n 0.004428f $X=2.465 $Y=3.295 $X2=2.42
+ $Y2=2.285
cc_231 N_VDD_M1019_b N_A_32_115#_c_685_n 0.0093744f $X=-0.045 $Y=2.425 $X2=0.285
+ $Y2=2.78
cc_232 N_VDD_M1019_b N_A_243_89#_M1009_g 0.0215131f $X=-0.045 $Y=2.425 $X2=1.89
+ $Y2=3.235
cc_233 N_VDD_c_192_p N_A_243_89#_M1009_g 0.00606474f $X=2.38 $Y=4.287 $X2=1.89
+ $Y2=3.235
cc_234 N_VDD_c_184_p N_A_243_89#_M1009_g 0.00468827f $X=6.46 $Y=4.25 $X2=1.89
+ $Y2=3.235
cc_235 N_VDD_M1019_b N_A_243_89#_M1000_g 0.0214821f $X=-0.045 $Y=2.425 $X2=3.04
+ $Y2=3.235
cc_236 N_VDD_c_203_p N_A_243_89#_M1000_g 0.00606474f $X=4.13 $Y=4.287 $X2=3.04
+ $Y2=3.235
cc_237 N_VDD_c_184_p N_A_243_89#_M1000_g 0.00468827f $X=6.46 $Y=4.25 $X2=3.04
+ $Y2=3.235
cc_238 N_VDD_M1019_b N_A_243_89#_c_792_n 0.00156053f $X=-0.045 $Y=2.425
+ $X2=4.645 $Y2=2.955
cc_239 N_VDD_c_208_p N_A_243_89#_c_792_n 0.00749582f $X=5.08 $Y=4.287 $X2=4.645
+ $Y2=2.955
cc_240 N_VDD_c_209_p N_A_243_89#_c_792_n 0.0341747f $X=5.165 $Y=3.295 $X2=4.645
+ $Y2=2.955
cc_241 N_VDD_c_184_p N_A_243_89#_c_792_n 0.00476261f $X=6.46 $Y=4.25 $X2=4.645
+ $Y2=2.955
cc_242 N_VDD_M1019_b N_A_243_89#_c_781_n 0.00543969f $X=-0.045 $Y=2.425
+ $X2=4.915 $Y2=2.62
cc_243 N_VDD_M1019_b N_A_243_89#_c_797_n 0.0119291f $X=-0.045 $Y=2.425 $X2=4.915
+ $Y2=2.705
cc_244 N_VDD_M1019_b N_A_785_89#_M1014_g 0.0178558f $X=-0.045 $Y=2.425 $X2=4
+ $Y2=3.235
cc_245 N_VDD_c_203_p N_A_785_89#_M1014_g 0.00606474f $X=4.13 $Y=4.287 $X2=4
+ $Y2=3.235
cc_246 N_VDD_c_207_p N_A_785_89#_M1014_g 0.0047242f $X=4.215 $Y=3.21 $X2=4
+ $Y2=3.235
cc_247 N_VDD_c_184_p N_A_785_89#_M1014_g 0.00468827f $X=6.46 $Y=4.25 $X2=4
+ $Y2=3.235
cc_248 N_VDD_M1019_b N_A_785_89#_M1006_g 0.0369702f $X=-0.045 $Y=2.425 $X2=6.33
+ $Y2=3.445
cc_249 N_VDD_c_249_p N_A_785_89#_M1006_g 0.00606474f $X=6.46 $Y=4.287 $X2=6.33
+ $Y2=3.445
cc_250 N_VDD_c_250_p N_A_785_89#_M1006_g 0.00354579f $X=6.545 $Y=3.615 $X2=6.33
+ $Y2=3.445
cc_251 N_VDD_c_184_p N_A_785_89#_M1006_g 0.00468827f $X=6.46 $Y=4.25 $X2=6.33
+ $Y2=3.445
cc_252 N_VDD_M1019_b N_A_785_89#_c_962_n 0.00284353f $X=-0.045 $Y=2.425
+ $X2=6.305 $Y2=2.475
cc_253 N_VDD_M1019_b N_A_785_89#_c_986_n 0.0134942f $X=-0.045 $Y=2.425 $X2=6.305
+ $Y2=2.625
cc_254 N_VDD_M1019_b N_A_785_89#_c_964_n 0.00241422f $X=-0.045 $Y=2.425 $X2=4.06
+ $Y2=2.48
cc_255 N_VDD_c_207_p N_A_785_89#_c_964_n 0.00121222f $X=4.215 $Y=3.21 $X2=4.06
+ $Y2=2.48
cc_256 N_VDD_M1019_b N_A_785_89#_c_968_n 0.00574079f $X=-0.045 $Y=2.425
+ $X2=5.595 $Y2=2.955
cc_257 N_VDD_c_249_p N_A_785_89#_c_968_n 0.0074445f $X=6.46 $Y=4.287 $X2=5.595
+ $Y2=2.955
cc_258 N_VDD_c_184_p N_A_785_89#_c_968_n 0.00476261f $X=6.46 $Y=4.25 $X2=5.595
+ $Y2=2.955
cc_259 N_VDD_M1019_b N_A_785_89#_c_971_n 0.011211f $X=-0.045 $Y=2.425 $X2=4.935
+ $Y2=2.48
cc_260 N_VDD_c_207_p N_A_785_89#_c_971_n 0.00492996f $X=4.215 $Y=3.21 $X2=4.935
+ $Y2=2.48
cc_261 N_VDD_M1019_b N_A_785_89#_c_972_n 0.00594013f $X=-0.045 $Y=2.425
+ $X2=4.205 $Y2=2.48
cc_262 N_VDD_c_207_p N_A_785_89#_c_972_n 0.00366258f $X=4.215 $Y=3.21 $X2=4.205
+ $Y2=2.48
cc_263 N_VDD_M1019_b N_A_623_115#_M1021_g 0.0260072f $X=-0.045 $Y=2.425 $X2=5.38
+ $Y2=3.235
cc_264 N_VDD_c_209_p N_A_623_115#_M1021_g 0.00636672f $X=5.165 $Y=3.295 $X2=5.38
+ $Y2=3.235
cc_265 N_VDD_c_249_p N_A_623_115#_M1021_g 0.00606474f $X=6.46 $Y=4.287 $X2=5.38
+ $Y2=3.235
cc_266 N_VDD_c_184_p N_A_623_115#_M1021_g 0.00468827f $X=6.46 $Y=4.25 $X2=5.38
+ $Y2=3.235
cc_267 N_VDD_M1019_b N_A_623_115#_c_1123_n 0.00168314f $X=-0.045 $Y=2.425
+ $X2=2.76 $Y2=1.37
cc_268 N_VDD_M1019_b N_A_623_115#_c_1142_n 0.00313975f $X=-0.045 $Y=2.425
+ $X2=3.34 $Y2=3.295
cc_269 N_VDD_c_203_p N_A_623_115#_c_1142_n 0.0151257f $X=4.13 $Y=4.287 $X2=3.34
+ $Y2=3.295
cc_270 N_VDD_c_184_p N_A_623_115#_c_1142_n 0.00958198f $X=6.46 $Y=4.25 $X2=3.34
+ $Y2=3.295
cc_271 N_VDD_M1019_b N_ON_M1020_g 0.0504657f $X=-0.045 $Y=2.425 $X2=6.76
+ $Y2=3.445
cc_272 N_VDD_c_250_p N_ON_M1020_g 0.00354579f $X=6.545 $Y=3.615 $X2=6.76
+ $Y2=3.445
cc_273 N_VDD_c_273_p N_ON_M1020_g 0.00606474f $X=6.46 $Y=4.25 $X2=6.76 $Y2=3.445
cc_274 N_VDD_c_184_p N_ON_M1020_g 0.00468827f $X=6.46 $Y=4.25 $X2=6.76 $Y2=3.445
cc_275 N_VDD_M1019_b N_ON_c_1245_n 0.0158117f $X=-0.045 $Y=2.425 $X2=6.115
+ $Y2=3.615
cc_276 N_VDD_c_249_p N_ON_c_1245_n 0.00757793f $X=6.46 $Y=4.287 $X2=6.115
+ $Y2=3.615
cc_277 N_VDD_c_184_p N_ON_c_1245_n 0.00476261f $X=6.46 $Y=4.25 $X2=6.115
+ $Y2=3.615
cc_278 N_VDD_M1019_b N_Q_c_1323_n 0.00156053f $X=-0.045 $Y=2.425 $X2=6.975
+ $Y2=3.615
cc_279 N_VDD_c_273_p N_Q_c_1323_n 0.00757793f $X=6.46 $Y=4.25 $X2=6.975
+ $Y2=3.615
cc_280 N_VDD_c_184_p N_Q_c_1323_n 0.00476261f $X=6.46 $Y=4.25 $X2=6.975
+ $Y2=3.615
cc_281 N_VDD_M1019_b N_Q_c_1320_n 0.0111162f $X=-0.045 $Y=2.425 $X2=7.09
+ $Y2=2.48
cc_282 N_VDD_M1019_b N_Q_c_1327_n 0.0150519f $X=-0.045 $Y=2.425 $X2=6.972
+ $Y2=2.88
cc_283 N_VDD_M1019_b N_Q_c_1328_n 0.00723753f $X=-0.045 $Y=2.425 $X2=6.972
+ $Y2=3.175
cc_284 N_VDD_M1019_b Q 0.00549803f $X=-0.045 $Y=2.425 $X2=6.97 $Y2=2.48
cc_285 N_A_75_248#_M1004_g N_D_M1003_g 0.0247367f $X=0.5 $Y=0.835 $X2=0.93
+ $Y2=0.835
cc_286 N_A_75_248#_c_291_n N_D_M1003_g 0.022942f $X=0.51 $Y=2.12 $X2=0.93
+ $Y2=0.835
cc_287 N_A_75_248#_c_292_n N_D_M1003_g 0.0146235f $X=1.405 $Y=1.285 $X2=0.93
+ $Y2=0.835
cc_288 N_A_75_248#_c_298_n N_D_M1003_g 0.00557207f $X=0.567 $Y=2.12 $X2=0.93
+ $Y2=0.835
cc_289 N_A_75_248#_M1019_g N_D_M1018_g 0.0342437f $X=0.5 $Y=3.235 $X2=0.93
+ $Y2=3.235
cc_290 N_A_75_248#_c_290_n N_D_M1018_g 0.0194268f $X=0.51 $Y=2.285 $X2=0.93
+ $Y2=3.235
cc_291 N_A_75_248#_c_307_n N_D_M1018_g 0.00557207f $X=0.625 $Y=2.62 $X2=0.93
+ $Y2=3.235
cc_292 N_A_75_248#_c_308_n N_D_M1018_g 0.019095f $X=1.42 $Y=2.705 $X2=0.93
+ $Y2=3.235
cc_293 N_A_75_248#_c_292_n N_D_c_377_n 0.00207628f $X=1.405 $Y=1.285 $X2=0.99
+ $Y2=1.74
cc_294 N_A_75_248#_c_297_n N_D_c_377_n 0.00557207f $X=0.51 $Y=2.285 $X2=0.99
+ $Y2=1.74
cc_295 N_A_75_248#_c_292_n N_D_c_378_n 0.0086486f $X=1.405 $Y=1.285 $X2=0.99
+ $Y2=1.74
cc_296 N_A_75_248#_c_298_n N_D_c_378_n 0.0187793f $X=0.567 $Y=2.12 $X2=0.99
+ $Y2=1.74
cc_297 N_A_75_248#_c_292_n D 0.00200799f $X=1.405 $Y=1.285 $X2=0.99 $Y2=1.74
cc_298 N_A_75_248#_c_298_n D 0.007232f $X=0.567 $Y=2.12 $X2=0.99 $Y2=1.74
cc_299 N_A_75_248#_c_308_n N_CK_M1013_g 0.0153724f $X=1.42 $Y=2.705 $X2=1.29
+ $Y2=3.235
cc_300 N_A_75_248#_c_308_n N_CK_c_417_n 0.00150627f $X=1.42 $Y=2.705 $X2=1.35
+ $Y2=2.285
cc_301 N_A_75_248#_c_292_n N_CK_c_418_n 9.45214e-19 $X=1.405 $Y=1.285 $X2=1.83
+ $Y2=1.37
cc_302 N_A_75_248#_c_299_n N_CK_c_418_n 0.00196448f $X=1.49 $Y=0.755 $X2=1.83
+ $Y2=1.37
cc_303 N_A_75_248#_c_296_n N_CK_c_419_n 0.00540119f $X=1.49 $Y=1.2 $X2=1.83
+ $Y2=1.205
cc_304 N_A_75_248#_c_292_n N_CK_c_433_n 0.0019742f $X=1.405 $Y=1.285 $X2=1.745
+ $Y2=2.11
cc_305 N_A_75_248#_c_308_n N_CK_c_433_n 0.00904674f $X=1.42 $Y=2.705 $X2=1.745
+ $Y2=2.11
cc_306 N_A_75_248#_c_292_n N_CK_c_434_n 0.012316f $X=1.405 $Y=1.285 $X2=1.83
+ $Y2=1.37
cc_307 N_A_75_248#_c_299_n N_CK_c_434_n 6.67366e-19 $X=1.49 $Y=0.755 $X2=1.83
+ $Y2=1.37
cc_308 N_A_75_248#_c_292_n N_CK_c_439_n 0.00224443f $X=1.405 $Y=1.285 $X2=1.35
+ $Y2=2.11
cc_309 N_A_75_248#_c_308_n N_CK_c_439_n 0.0101098f $X=1.42 $Y=2.705 $X2=1.35
+ $Y2=2.11
cc_310 N_A_75_248#_c_298_n N_CK_c_439_n 0.0103407f $X=0.567 $Y=2.12 $X2=1.35
+ $Y2=2.11
cc_311 N_A_75_248#_c_308_n N_CK_c_441_n 0.00613532f $X=1.42 $Y=2.705 $X2=3.435
+ $Y2=2.11
cc_312 N_A_75_248#_c_308_n N_CK_c_442_n 0.00409373f $X=1.42 $Y=2.705 $X2=1.495
+ $Y2=2.11
cc_313 N_A_75_248#_c_298_n N_CK_c_442_n 0.00642105f $X=0.567 $Y=2.12 $X2=1.495
+ $Y2=2.11
cc_314 N_A_75_248#_M1019_g N_A_32_115#_c_658_n 0.00498045f $X=0.5 $Y=3.235
+ $X2=0.17 $Y2=2.695
cc_315 N_A_75_248#_c_291_n N_A_32_115#_c_658_n 0.0218335f $X=0.51 $Y=2.12
+ $X2=0.17 $Y2=2.695
cc_316 N_A_75_248#_c_307_n N_A_32_115#_c_658_n 0.00821014f $X=0.625 $Y=2.62
+ $X2=0.17 $Y2=2.695
cc_317 N_A_75_248#_c_310_n N_A_32_115#_c_658_n 0.00395316f $X=0.71 $Y=2.705
+ $X2=0.17 $Y2=2.695
cc_318 N_A_75_248#_c_297_n N_A_32_115#_c_658_n 0.0245251f $X=0.51 $Y=2.285
+ $X2=0.17 $Y2=2.695
cc_319 N_A_75_248#_c_298_n N_A_32_115#_c_658_n 0.0334082f $X=0.567 $Y=2.12
+ $X2=0.17 $Y2=2.695
cc_320 N_A_75_248#_M1004_g N_A_32_115#_c_659_n 0.00605682f $X=0.5 $Y=0.835
+ $X2=0.285 $Y2=0.755
cc_321 N_A_75_248#_M1004_g N_A_32_115#_c_663_n 0.00165831f $X=0.5 $Y=0.835
+ $X2=0.285 $Y2=1.37
cc_322 N_A_75_248#_c_289_n N_A_32_115#_c_663_n 0.00460749f $X=0.475 $Y=1.39
+ $X2=0.285 $Y2=1.37
cc_323 N_A_75_248#_c_294_n N_A_32_115#_c_663_n 0.0125535f $X=0.71 $Y=1.285
+ $X2=0.285 $Y2=1.37
cc_324 N_A_75_248#_c_298_n N_A_32_115#_c_663_n 0.00592135f $X=0.567 $Y=2.12
+ $X2=0.285 $Y2=1.37
cc_325 N_A_75_248#_c_289_n N_A_32_115#_c_666_n 0.0047054f $X=0.475 $Y=1.39
+ $X2=2.185 $Y2=1.37
cc_326 N_A_75_248#_c_291_n N_A_32_115#_c_666_n 0.0043937f $X=0.51 $Y=2.12
+ $X2=2.185 $Y2=1.37
cc_327 N_A_75_248#_c_292_n N_A_32_115#_c_666_n 0.0597745f $X=1.405 $Y=1.285
+ $X2=2.185 $Y2=1.37
cc_328 N_A_75_248#_c_294_n N_A_32_115#_c_666_n 0.00750079f $X=0.71 $Y=1.285
+ $X2=2.185 $Y2=1.37
cc_329 N_A_75_248#_c_298_n N_A_32_115#_c_666_n 0.0143756f $X=0.567 $Y=2.12
+ $X2=2.185 $Y2=1.37
cc_330 N_A_75_248#_c_299_n N_A_32_115#_c_666_n 0.00707072f $X=1.49 $Y=0.755
+ $X2=2.185 $Y2=1.37
cc_331 N_A_75_248#_c_289_n N_A_32_115#_c_668_n 0.00387046f $X=0.475 $Y=1.39
+ $X2=0.43 $Y2=1.37
cc_332 N_A_75_248#_c_291_n N_A_32_115#_c_668_n 0.00369116f $X=0.51 $Y=2.12
+ $X2=0.43 $Y2=1.37
cc_333 N_A_75_248#_c_294_n N_A_32_115#_c_668_n 8.15236e-19 $X=0.71 $Y=1.285
+ $X2=0.43 $Y2=1.37
cc_334 N_A_75_248#_c_298_n N_A_32_115#_c_668_n 8.59347e-19 $X=0.567 $Y=2.12
+ $X2=0.43 $Y2=1.37
cc_335 N_A_75_248#_c_292_n N_A_243_89#_c_759_n 0.0066768f $X=1.405 $Y=1.285
+ $X2=1.29 $Y2=1.205
cc_336 N_A_75_248#_c_296_n N_A_243_89#_c_759_n 0.00377845f $X=1.49 $Y=1.2
+ $X2=1.29 $Y2=1.205
cc_337 N_A_75_248#_c_292_n N_A_243_89#_c_762_n 0.00326059f $X=1.405 $Y=1.285
+ $X2=1.41 $Y2=1.745
cc_338 N_A_75_248#_c_292_n N_A_243_89#_c_763_n 0.00156949f $X=1.405 $Y=1.285
+ $X2=1.815 $Y2=1.82
cc_339 N_A_75_248#_c_292_n N_A_243_89#_c_772_n 0.00984832f $X=1.405 $Y=1.285
+ $X2=1.41 $Y2=1.28
cc_340 N_A_75_248#_c_308_n A_201_521# 0.00732587f $X=1.42 $Y=2.705 $X2=1.005
+ $Y2=2.605
cc_341 N_D_M1018_g N_CK_c_417_n 0.113471f $X=0.93 $Y=3.235 $X2=1.35 $Y2=2.285
cc_342 N_D_c_377_n N_CK_c_434_n 2.89615e-19 $X=0.99 $Y=1.74 $X2=1.83 $Y2=1.37
cc_343 N_D_c_378_n N_CK_c_434_n 0.00478177f $X=0.99 $Y=1.74 $X2=1.83 $Y2=1.37
cc_344 D N_CK_c_434_n 0.00551577f $X=0.99 $Y=1.74 $X2=1.83 $Y2=1.37
cc_345 N_D_M1018_g N_CK_c_439_n 0.0030898f $X=0.93 $Y=3.235 $X2=1.35 $Y2=2.11
cc_346 N_D_M1018_g N_CK_c_442_n 0.00515433f $X=0.93 $Y=3.235 $X2=1.495 $Y2=2.11
cc_347 D N_CK_c_442_n 0.00375733f $X=0.99 $Y=1.74 $X2=1.495 $Y2=2.11
cc_348 N_D_M1003_g N_A_32_115#_c_666_n 0.00223521f $X=0.93 $Y=0.835 $X2=2.185
+ $Y2=1.37
cc_349 N_D_c_377_n N_A_32_115#_c_666_n 7.9412e-19 $X=0.99 $Y=1.74 $X2=2.185
+ $Y2=1.37
cc_350 N_D_c_378_n N_A_32_115#_c_666_n 0.00111625f $X=0.99 $Y=1.74 $X2=2.185
+ $Y2=1.37
cc_351 D N_A_32_115#_c_666_n 0.0353362f $X=0.99 $Y=1.74 $X2=2.185 $Y2=1.37
cc_352 N_D_M1003_g N_A_243_89#_c_759_n 0.0553906f $X=0.93 $Y=0.835 $X2=1.29
+ $Y2=1.205
cc_353 N_D_M1003_g N_A_243_89#_c_762_n 0.00886317f $X=0.93 $Y=0.835 $X2=1.41
+ $Y2=1.745
cc_354 N_D_c_377_n N_A_243_89#_c_762_n 0.0210215f $X=0.99 $Y=1.74 $X2=1.41
+ $Y2=1.745
cc_355 N_D_c_378_n N_A_243_89#_c_762_n 0.00164409f $X=0.99 $Y=1.74 $X2=1.41
+ $Y2=1.745
cc_356 D N_A_243_89#_c_762_n 0.00342011f $X=0.99 $Y=1.74 $X2=1.41 $Y2=1.745
cc_357 D N_A_243_89#_c_764_n 4.62757e-19 $X=0.99 $Y=1.74 $X2=1.485 $Y2=1.82
cc_358 N_CK_c_419_n N_A_32_115#_M1011_g 0.0333294f $X=1.83 $Y=1.205 $X2=2.25
+ $Y2=0.835
cc_359 N_CK_c_434_n N_A_32_115#_M1011_g 0.00109079f $X=1.83 $Y=1.37 $X2=2.25
+ $Y2=0.835
cc_360 N_CK_c_422_n N_A_32_115#_c_649_n 0.0329411f $X=3.1 $Y=1.37 $X2=2.605
+ $Y2=1.37
cc_361 N_CK_c_435_n N_A_32_115#_c_649_n 2.90013e-19 $X=3.1 $Y=1.37 $X2=2.605
+ $Y2=1.37
cc_362 N_CK_c_418_n N_A_32_115#_c_651_n 0.0333294f $X=1.83 $Y=1.37 $X2=2.325
+ $Y2=1.37
cc_363 N_CK_c_441_n N_A_32_115#_c_652_n 0.00772879f $X=3.435 $Y=2.11 $X2=2.605
+ $Y2=2.285
cc_364 N_CK_c_441_n N_A_32_115#_c_653_n 0.00679967f $X=3.435 $Y=2.11 $X2=2.325
+ $Y2=2.285
cc_365 N_CK_c_423_n N_A_32_115#_M1012_g 0.0329411f $X=3.1 $Y=1.205 $X2=2.68
+ $Y2=0.835
cc_366 N_CK_c_435_n N_A_32_115#_M1012_g 2.72781e-19 $X=3.1 $Y=1.37 $X2=2.68
+ $Y2=0.835
cc_367 N_CK_c_418_n N_A_32_115#_c_662_n 7.30049e-19 $X=1.83 $Y=1.37 $X2=2.42
+ $Y2=2.285
cc_368 N_CK_c_433_n N_A_32_115#_c_662_n 0.00401809f $X=1.745 $Y=2.11 $X2=2.42
+ $Y2=2.285
cc_369 N_CK_c_434_n N_A_32_115#_c_662_n 0.0203851f $X=1.83 $Y=1.37 $X2=2.42
+ $Y2=2.285
cc_370 N_CK_c_441_n N_A_32_115#_c_662_n 0.0206884f $X=3.435 $Y=2.11 $X2=2.42
+ $Y2=2.285
cc_371 N_CK_c_418_n N_A_32_115#_c_664_n 7.18106e-19 $X=1.83 $Y=1.37 $X2=2.42
+ $Y2=1.37
cc_372 N_CK_c_434_n N_A_32_115#_c_664_n 0.00742068f $X=1.83 $Y=1.37 $X2=2.42
+ $Y2=1.37
cc_373 N_CK_c_435_n N_A_32_115#_c_664_n 0.00183328f $X=3.1 $Y=1.37 $X2=2.42
+ $Y2=1.37
cc_374 N_CK_c_441_n N_A_32_115#_c_664_n 0.00102309f $X=3.435 $Y=2.11 $X2=2.42
+ $Y2=1.37
cc_375 N_CK_c_418_n N_A_32_115#_c_666_n 0.00576782f $X=1.83 $Y=1.37 $X2=2.185
+ $Y2=1.37
cc_376 N_CK_c_433_n N_A_32_115#_c_666_n 0.00443421f $X=1.745 $Y=2.11 $X2=2.185
+ $Y2=1.37
cc_377 N_CK_c_434_n N_A_32_115#_c_666_n 0.0204779f $X=1.83 $Y=1.37 $X2=2.185
+ $Y2=1.37
cc_378 N_CK_c_439_n N_A_32_115#_c_666_n 7.12046e-19 $X=1.35 $Y=2.11 $X2=2.185
+ $Y2=1.37
cc_379 N_CK_c_442_n N_A_32_115#_c_666_n 0.0126164f $X=1.495 $Y=2.11 $X2=2.185
+ $Y2=1.37
cc_380 N_CK_c_418_n N_A_32_115#_c_669_n 3.3031e-19 $X=1.83 $Y=1.37 $X2=2.33
+ $Y2=1.37
cc_381 N_CK_c_434_n N_A_32_115#_c_669_n 0.00143592f $X=1.83 $Y=1.37 $X2=2.33
+ $Y2=1.37
cc_382 N_CK_c_441_n N_A_32_115#_c_669_n 0.0129652f $X=3.435 $Y=2.11 $X2=2.33
+ $Y2=1.37
cc_383 N_CK_c_419_n N_A_243_89#_c_759_n 0.0152095f $X=1.83 $Y=1.205 $X2=1.29
+ $Y2=1.205
cc_384 N_CK_c_434_n N_A_243_89#_c_762_n 0.00613747f $X=1.83 $Y=1.37 $X2=1.41
+ $Y2=1.745
cc_385 N_CK_c_418_n N_A_243_89#_c_763_n 0.0183603f $X=1.83 $Y=1.37 $X2=1.815
+ $Y2=1.82
cc_386 N_CK_c_434_n N_A_243_89#_c_763_n 0.00630484f $X=1.83 $Y=1.37 $X2=1.815
+ $Y2=1.82
cc_387 N_CK_c_441_n N_A_243_89#_c_763_n 0.00558832f $X=3.435 $Y=2.11 $X2=1.815
+ $Y2=1.82
cc_388 N_CK_c_417_n N_A_243_89#_c_764_n 0.00904036f $X=1.35 $Y=2.285 $X2=1.485
+ $Y2=1.82
cc_389 N_CK_c_433_n N_A_243_89#_c_764_n 0.00810782f $X=1.745 $Y=2.11 $X2=1.485
+ $Y2=1.82
cc_390 N_CK_c_439_n N_A_243_89#_c_764_n 0.00109468f $X=1.35 $Y=2.11 $X2=1.485
+ $Y2=1.82
cc_391 N_CK_c_442_n N_A_243_89#_c_764_n 0.00131242f $X=1.495 $Y=2.11 $X2=1.485
+ $Y2=1.82
cc_392 N_CK_M1013_g N_A_243_89#_M1009_g 0.0315947f $X=1.29 $Y=3.235 $X2=1.89
+ $Y2=3.235
cc_393 N_CK_c_417_n N_A_243_89#_M1009_g 0.0128384f $X=1.35 $Y=2.285 $X2=1.89
+ $Y2=3.235
cc_394 N_CK_c_433_n N_A_243_89#_M1009_g 0.0081071f $X=1.745 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_395 N_CK_c_434_n N_A_243_89#_M1009_g 0.00478024f $X=1.83 $Y=1.37 $X2=1.89
+ $Y2=3.235
cc_396 N_CK_c_439_n N_A_243_89#_M1009_g 0.00184124f $X=1.35 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_397 N_CK_c_441_n N_A_243_89#_M1009_g 0.00938974f $X=3.435 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_398 N_CK_c_442_n N_A_243_89#_M1009_g 4.2e-19 $X=1.495 $Y=2.11 $X2=1.89
+ $Y2=3.235
cc_399 N_CK_c_441_n N_A_243_89#_c_766_n 0.00607908f $X=3.435 $Y=2.11 $X2=2.965
+ $Y2=1.82
cc_400 N_CK_M1017_g N_A_243_89#_M1000_g 0.0316011f $X=3.64 $Y=3.235 $X2=3.04
+ $Y2=3.235
cc_401 N_CK_c_426_n N_A_243_89#_M1000_g 0.0118393f $X=3.58 $Y=2.285 $X2=3.04
+ $Y2=3.235
cc_402 N_CK_c_435_n N_A_243_89#_M1000_g 0.00368284f $X=3.1 $Y=1.37 $X2=3.04
+ $Y2=3.235
cc_403 N_CK_c_437_n N_A_243_89#_M1000_g 0.00654233f $X=3.185 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_404 N_CK_c_440_n N_A_243_89#_M1000_g 0.00128351f $X=3.58 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_405 N_CK_c_441_n N_A_243_89#_M1000_g 0.00497421f $X=3.435 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_406 N_CK_c_444_n N_A_243_89#_M1000_g 4.2e-19 $X=3.725 $Y=2.11 $X2=3.04
+ $Y2=3.235
cc_407 N_CK_c_435_n N_A_243_89#_c_768_n 0.00679428f $X=3.1 $Y=1.37 $X2=3.445
+ $Y2=1.825
cc_408 N_CK_c_436_n N_A_243_89#_c_768_n 0.00791072f $X=3.495 $Y=2.11 $X2=3.445
+ $Y2=1.825
cc_409 N_CK_c_441_n N_A_243_89#_c_768_n 0.00549267f $X=3.435 $Y=2.11 $X2=3.445
+ $Y2=1.825
cc_410 N_CK_c_444_n N_A_243_89#_c_768_n 0.00125393f $X=3.725 $Y=2.11 $X2=3.445
+ $Y2=1.825
cc_411 N_CK_c_422_n N_A_243_89#_M1001_g 0.0129208f $X=3.1 $Y=1.37 $X2=3.64
+ $Y2=0.835
cc_412 N_CK_c_423_n N_A_243_89#_M1001_g 0.0151224f $X=3.1 $Y=1.205 $X2=3.64
+ $Y2=0.835
cc_413 N_CK_c_435_n N_A_243_89#_M1001_g 0.00166016f $X=3.1 $Y=1.37 $X2=3.64
+ $Y2=0.835
cc_414 N_CK_c_418_n N_A_243_89#_c_772_n 0.0216263f $X=1.83 $Y=1.37 $X2=1.41
+ $Y2=1.28
cc_415 N_CK_c_439_n N_A_243_89#_c_772_n 2.45465e-19 $X=1.35 $Y=2.11 $X2=1.41
+ $Y2=1.28
cc_416 N_CK_c_434_n N_A_243_89#_c_773_n 0.00568091f $X=1.83 $Y=1.37 $X2=1.89
+ $Y2=1.82
cc_417 N_CK_c_422_n N_A_243_89#_c_774_n 0.0183777f $X=3.1 $Y=1.37 $X2=3.04
+ $Y2=1.825
cc_418 N_CK_c_435_n N_A_243_89#_c_774_n 0.00451735f $X=3.1 $Y=1.37 $X2=3.04
+ $Y2=1.825
cc_419 N_CK_c_426_n N_A_243_89#_c_775_n 0.017377f $X=3.58 $Y=2.285 $X2=3.58
+ $Y2=1.74
cc_420 N_CK_c_435_n N_A_243_89#_c_775_n 0.00308518f $X=3.1 $Y=1.37 $X2=3.58
+ $Y2=1.74
cc_421 N_CK_c_440_n N_A_243_89#_c_775_n 0.00108353f $X=3.58 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_422 N_CK_c_426_n N_A_243_89#_c_776_n 7.72371e-19 $X=3.58 $Y=2.285 $X2=3.58
+ $Y2=1.74
cc_423 N_CK_c_435_n N_A_243_89#_c_776_n 0.00780691f $X=3.1 $Y=1.37 $X2=3.58
+ $Y2=1.74
cc_424 N_CK_c_436_n N_A_243_89#_c_776_n 0.00456947f $X=3.495 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_425 N_CK_c_440_n N_A_243_89#_c_776_n 0.00979766f $X=3.58 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_426 N_CK_c_443_n N_A_243_89#_c_776_n 5.17303e-19 $X=4.43 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_427 N_CK_c_444_n N_A_243_89#_c_776_n 0.00182452f $X=3.725 $Y=2.11 $X2=3.58
+ $Y2=1.74
cc_428 N_CK_c_427_n N_A_243_89#_c_777_n 0.00700796f $X=4.457 $Y=1.205 $X2=4.645
+ $Y2=0.755
cc_429 N_CK_c_432_n N_A_243_89#_c_777_n 0.0118432f $X=4.457 $Y=1.355 $X2=4.645
+ $Y2=0.755
cc_430 N_CK_c_415_n N_A_243_89#_c_781_n 0.00318866f $X=4.43 $Y=2.45 $X2=4.915
+ $Y2=2.62
cc_431 N_CK_M1015_g N_A_243_89#_c_781_n 0.00395773f $X=4.43 $Y=3.235 $X2=4.915
+ $Y2=2.62
cc_432 N_CK_c_416_n N_A_243_89#_c_781_n 0.00643904f $X=4.485 $Y=2.12 $X2=4.915
+ $Y2=2.62
cc_433 N_CK_c_438_n N_A_243_89#_c_781_n 0.0277441f $X=4.575 $Y=2.11 $X2=4.915
+ $Y2=2.62
cc_434 CK N_A_243_89#_c_781_n 0.00256489f $X=4.575 $Y=2.11 $X2=4.915 $Y2=2.62
cc_435 N_CK_c_415_n N_A_243_89#_c_782_n 0.0016621f $X=4.43 $Y=2.45 $X2=4.915
+ $Y2=1.725
cc_436 N_CK_c_416_n N_A_243_89#_c_782_n 0.00536103f $X=4.485 $Y=2.12 $X2=4.915
+ $Y2=1.725
cc_437 N_CK_c_438_n N_A_243_89#_c_782_n 0.00607622f $X=4.575 $Y=2.11 $X2=4.915
+ $Y2=1.725
cc_438 CK N_A_243_89#_c_782_n 7.74944e-19 $X=4.575 $Y=2.11 $X2=4.915 $Y2=1.725
cc_439 N_CK_c_415_n N_A_243_89#_c_797_n 0.00233394f $X=4.43 $Y=2.45 $X2=4.915
+ $Y2=2.705
cc_440 N_CK_c_438_n N_A_243_89#_c_797_n 0.00601935f $X=4.575 $Y=2.11 $X2=4.915
+ $Y2=2.705
cc_441 N_CK_c_435_n N_A_243_89#_c_783_n 0.00361908f $X=3.1 $Y=1.37 $X2=3.725
+ $Y2=1.725
cc_442 N_CK_c_436_n N_A_243_89#_c_783_n 2.38605e-19 $X=3.495 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_443 N_CK_c_440_n N_A_243_89#_c_783_n 4.76324e-19 $X=3.58 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_444 N_CK_c_441_n N_A_243_89#_c_783_n 0.00163817f $X=3.435 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_445 N_CK_c_444_n N_A_243_89#_c_783_n 0.0296305f $X=3.725 $Y=2.11 $X2=3.725
+ $Y2=1.725
cc_446 N_CK_c_415_n N_A_243_89#_c_784_n 2.36275e-19 $X=4.43 $Y=2.45 $X2=4.645
+ $Y2=1.74
cc_447 N_CK_c_416_n N_A_243_89#_c_784_n 0.00216028f $X=4.485 $Y=2.12 $X2=4.645
+ $Y2=1.74
cc_448 N_CK_c_438_n N_A_243_89#_c_784_n 0.00129914f $X=4.575 $Y=2.11 $X2=4.645
+ $Y2=1.74
cc_449 CK N_A_243_89#_c_784_n 0.0226506f $X=4.575 $Y=2.11 $X2=4.645 $Y2=1.74
cc_450 N_CK_c_416_n N_A_243_89#_c_785_n 0.00278025f $X=4.485 $Y=2.12 $X2=4.5
+ $Y2=1.74
cc_451 N_CK_c_432_n N_A_243_89#_c_785_n 2.64649e-19 $X=4.457 $Y=1.355 $X2=4.5
+ $Y2=1.74
cc_452 N_CK_c_443_n N_A_243_89#_c_785_n 0.0538111f $X=4.43 $Y=2.11 $X2=4.5
+ $Y2=1.74
cc_453 CK N_A_243_89#_c_785_n 0.00582134f $X=4.575 $Y=2.11 $X2=4.5 $Y2=1.74
cc_454 N_CK_c_416_n N_A_785_89#_M1023_g 0.00866378f $X=4.485 $Y=2.12 $X2=4
+ $Y2=0.835
cc_455 N_CK_c_427_n N_A_785_89#_M1023_g 0.0236863f $X=4.457 $Y=1.205 $X2=4
+ $Y2=0.835
cc_456 N_CK_c_415_n N_A_785_89#_M1014_g 0.0389285f $X=4.43 $Y=2.45 $X2=4
+ $Y2=3.235
cc_457 N_CK_c_416_n N_A_785_89#_M1014_g 0.0139901f $X=4.485 $Y=2.12 $X2=4
+ $Y2=3.235
cc_458 N_CK_c_426_n N_A_785_89#_M1014_g 0.11248f $X=3.58 $Y=2.285 $X2=4
+ $Y2=3.235
cc_459 N_CK_c_438_n N_A_785_89#_M1014_g 5.87562e-19 $X=4.575 $Y=2.11 $X2=4
+ $Y2=3.235
cc_460 N_CK_c_440_n N_A_785_89#_M1014_g 0.0022769f $X=3.58 $Y=2.11 $X2=4
+ $Y2=3.235
cc_461 N_CK_c_443_n N_A_785_89#_M1014_g 0.00290457f $X=4.43 $Y=2.11 $X2=4
+ $Y2=3.235
cc_462 N_CK_c_444_n N_A_785_89#_M1014_g 0.00113587f $X=3.725 $Y=2.11 $X2=4
+ $Y2=3.235
cc_463 N_CK_c_416_n N_A_785_89#_c_960_n 0.0205813f $X=4.485 $Y=2.12 $X2=4.06
+ $Y2=1.74
cc_464 N_CK_c_443_n N_A_785_89#_c_960_n 7.38456e-19 $X=4.43 $Y=2.11 $X2=4.06
+ $Y2=1.74
cc_465 N_CK_c_416_n N_A_785_89#_c_963_n 8.19109e-19 $X=4.485 $Y=2.12 $X2=4.062
+ $Y2=1.812
cc_466 N_CK_c_415_n N_A_785_89#_c_964_n 0.00276728f $X=4.43 $Y=2.45 $X2=4.06
+ $Y2=2.48
cc_467 N_CK_c_416_n N_A_785_89#_c_964_n 0.00446139f $X=4.485 $Y=2.12 $X2=4.06
+ $Y2=2.48
cc_468 N_CK_c_426_n N_A_785_89#_c_964_n 0.00225599f $X=3.58 $Y=2.285 $X2=4.06
+ $Y2=2.48
cc_469 N_CK_c_438_n N_A_785_89#_c_964_n 0.0149594f $X=4.575 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_470 N_CK_c_440_n N_A_785_89#_c_964_n 0.0150983f $X=3.58 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_471 N_CK_c_443_n N_A_785_89#_c_964_n 0.0141643f $X=4.43 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_472 N_CK_c_444_n N_A_785_89#_c_964_n 0.00206546f $X=3.725 $Y=2.11 $X2=4.06
+ $Y2=2.48
cc_473 CK N_A_785_89#_c_964_n 0.00191287f $X=4.575 $Y=2.11 $X2=4.06 $Y2=2.48
cc_474 N_CK_c_415_n N_A_785_89#_c_971_n 0.00433056f $X=4.43 $Y=2.45 $X2=4.935
+ $Y2=2.48
cc_475 N_CK_M1015_g N_A_785_89#_c_971_n 0.00888384f $X=4.43 $Y=3.235 $X2=4.935
+ $Y2=2.48
cc_476 N_CK_c_438_n N_A_785_89#_c_971_n 0.00642492f $X=4.575 $Y=2.11 $X2=4.935
+ $Y2=2.48
cc_477 N_CK_c_443_n N_A_785_89#_c_971_n 0.0190758f $X=4.43 $Y=2.11 $X2=4.935
+ $Y2=2.48
cc_478 CK N_A_785_89#_c_971_n 0.025144f $X=4.575 $Y=2.11 $X2=4.935 $Y2=2.48
cc_479 N_CK_c_415_n N_A_785_89#_c_972_n 4.83733e-19 $X=4.43 $Y=2.45 $X2=4.205
+ $Y2=2.48
cc_480 N_CK_M1015_g N_A_785_89#_c_972_n 4.63789e-19 $X=4.43 $Y=3.235 $X2=4.205
+ $Y2=2.48
cc_481 N_CK_c_426_n N_A_785_89#_c_972_n 0.00405956f $X=3.58 $Y=2.285 $X2=4.205
+ $Y2=2.48
cc_482 N_CK_c_438_n N_A_785_89#_c_972_n 7.97287e-19 $X=4.575 $Y=2.11 $X2=4.205
+ $Y2=2.48
cc_483 N_CK_c_440_n N_A_785_89#_c_972_n 0.0025579f $X=3.58 $Y=2.11 $X2=4.205
+ $Y2=2.48
cc_484 N_CK_c_443_n N_A_785_89#_c_972_n 0.0252575f $X=4.43 $Y=2.11 $X2=4.205
+ $Y2=2.48
cc_485 N_CK_c_438_n N_A_785_89#_c_973_n 0.00120049f $X=4.575 $Y=2.11 $X2=5.007
+ $Y2=2.395
cc_486 CK N_A_785_89#_c_973_n 0.0189169f $X=4.575 $Y=2.11 $X2=5.007 $Y2=2.395
cc_487 N_CK_c_415_n N_A_623_115#_M1021_g 0.00468822f $X=4.43 $Y=2.45 $X2=5.38
+ $Y2=3.235
cc_488 N_CK_c_432_n N_A_623_115#_c_1121_n 0.00712865f $X=4.457 $Y=1.355 $X2=5.38
+ $Y2=1.37
cc_489 N_CK_c_422_n N_A_623_115#_c_1123_n 0.00171905f $X=3.1 $Y=1.37 $X2=2.76
+ $Y2=1.37
cc_490 N_CK_c_435_n N_A_623_115#_c_1123_n 0.0516647f $X=3.1 $Y=1.37 $X2=2.76
+ $Y2=1.37
cc_491 N_CK_c_437_n N_A_623_115#_c_1123_n 0.0116326f $X=3.185 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_492 N_CK_c_440_n N_A_623_115#_c_1123_n 0.00613815f $X=3.58 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_493 N_CK_c_441_n N_A_623_115#_c_1123_n 0.020361f $X=3.435 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_494 N_CK_c_444_n N_A_623_115#_c_1123_n 6.61118e-19 $X=3.725 $Y=2.11 $X2=2.76
+ $Y2=1.37
cc_495 N_CK_c_426_n N_A_623_115#_c_1153_n 0.00150627f $X=3.58 $Y=2.285 $X2=3.17
+ $Y2=2.705
cc_496 N_CK_c_436_n N_A_623_115#_c_1153_n 0.00843004f $X=3.495 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_497 N_CK_c_437_n N_A_623_115#_c_1153_n 0.00323798f $X=3.185 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_498 N_CK_c_440_n N_A_623_115#_c_1153_n 0.00103871f $X=3.58 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_499 N_CK_c_441_n N_A_623_115#_c_1153_n 0.012754f $X=3.435 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_500 N_CK_c_444_n N_A_623_115#_c_1153_n 0.00146098f $X=3.725 $Y=2.11 $X2=3.17
+ $Y2=2.705
cc_501 N_CK_c_422_n N_A_623_115#_c_1124_n 0.0015339f $X=3.1 $Y=1.37 $X2=3.44
+ $Y2=1.34
cc_502 N_CK_c_423_n N_A_623_115#_c_1124_n 0.00346504f $X=3.1 $Y=1.205 $X2=3.44
+ $Y2=1.34
cc_503 N_CK_c_435_n N_A_623_115#_c_1124_n 0.0166762f $X=3.1 $Y=1.37 $X2=3.44
+ $Y2=1.34
cc_504 N_CK_c_436_n N_A_623_115#_c_1124_n 0.00112312f $X=3.495 $Y=2.11 $X2=3.44
+ $Y2=1.34
cc_505 N_CK_c_441_n N_A_623_115#_c_1124_n 9.66728e-19 $X=3.435 $Y=2.11 $X2=3.44
+ $Y2=1.34
cc_506 N_CK_c_422_n N_A_623_115#_c_1127_n 0.00224296f $X=3.1 $Y=1.37 $X2=3.34
+ $Y2=0.755
cc_507 N_CK_c_435_n N_A_623_115#_c_1127_n 9.81838e-19 $X=3.1 $Y=1.37 $X2=3.34
+ $Y2=0.755
cc_508 N_CK_c_422_n N_A_623_115#_c_1130_n 0.00610106f $X=3.1 $Y=1.37 $X2=3.295
+ $Y2=1.37
cc_509 N_CK_c_435_n N_A_623_115#_c_1130_n 0.0178696f $X=3.1 $Y=1.37 $X2=3.295
+ $Y2=1.37
cc_510 N_CK_c_436_n N_A_623_115#_c_1130_n 0.00291459f $X=3.495 $Y=2.11 $X2=3.295
+ $Y2=1.37
cc_511 N_CK_c_422_n N_A_623_115#_c_1131_n 6.81488e-19 $X=3.1 $Y=1.37 $X2=2.905
+ $Y2=1.37
cc_512 N_CK_c_435_n N_A_623_115#_c_1131_n 0.00134743f $X=3.1 $Y=1.37 $X2=2.905
+ $Y2=1.37
cc_513 N_CK_c_441_n N_A_623_115#_c_1131_n 0.0128239f $X=3.435 $Y=2.11 $X2=2.905
+ $Y2=1.37
cc_514 N_CK_c_416_n N_A_623_115#_c_1132_n 0.00321559f $X=4.485 $Y=2.12 $X2=5.03
+ $Y2=1.37
cc_515 N_CK_c_432_n N_A_623_115#_c_1132_n 0.0102303f $X=4.457 $Y=1.355 $X2=5.03
+ $Y2=1.37
cc_516 N_CK_c_422_n N_A_623_115#_c_1134_n 7.09529e-19 $X=3.1 $Y=1.37 $X2=3.585
+ $Y2=1.37
cc_517 N_CK_c_435_n N_A_623_115#_c_1134_n 0.00114929f $X=3.1 $Y=1.37 $X2=3.585
+ $Y2=1.37
cc_518 N_A_32_115#_c_666_n N_A_243_89#_c_762_n 0.00252532f $X=2.185 $Y=1.37
+ $X2=1.41 $Y2=1.745
cc_519 N_A_32_115#_c_666_n N_A_243_89#_c_763_n 0.004711f $X=2.185 $Y=1.37
+ $X2=1.815 $Y2=1.82
cc_520 N_A_32_115#_c_653_n N_A_243_89#_M1009_g 0.113994f $X=2.325 $Y=2.285
+ $X2=1.89 $Y2=3.235
cc_521 N_A_32_115#_c_662_n N_A_243_89#_M1009_g 0.00486364f $X=2.42 $Y=2.285
+ $X2=1.89 $Y2=3.235
cc_522 N_A_32_115#_c_651_n N_A_243_89#_c_766_n 0.0342351f $X=2.325 $Y=1.37
+ $X2=2.965 $Y2=1.82
cc_523 N_A_32_115#_c_653_n N_A_243_89#_c_766_n 0.0307748f $X=2.325 $Y=2.285
+ $X2=2.965 $Y2=1.82
cc_524 N_A_32_115#_c_662_n N_A_243_89#_c_766_n 0.0113171f $X=2.42 $Y=2.285
+ $X2=2.965 $Y2=1.82
cc_525 N_A_32_115#_c_664_n N_A_243_89#_c_766_n 8.69982e-19 $X=2.42 $Y=1.37
+ $X2=2.965 $Y2=1.82
cc_526 N_A_32_115#_c_666_n N_A_243_89#_c_766_n 0.00486036f $X=2.185 $Y=1.37
+ $X2=2.965 $Y2=1.82
cc_527 N_A_32_115#_c_669_n N_A_243_89#_c_766_n 4.12801e-19 $X=2.33 $Y=1.37
+ $X2=2.965 $Y2=1.82
cc_528 N_A_32_115#_c_652_n N_A_243_89#_M1000_g 0.110621f $X=2.605 $Y=2.285
+ $X2=3.04 $Y2=3.235
cc_529 N_A_32_115#_M1002_g N_A_623_115#_c_1123_n 9.36754e-19 $X=2.25 $Y=3.235
+ $X2=2.76 $Y2=1.37
cc_530 N_A_32_115#_c_649_n N_A_623_115#_c_1123_n 0.0070068f $X=2.605 $Y=1.37
+ $X2=2.76 $Y2=1.37
cc_531 N_A_32_115#_c_652_n N_A_623_115#_c_1123_n 0.00738718f $X=2.605 $Y=2.285
+ $X2=2.76 $Y2=1.37
cc_532 N_A_32_115#_M1005_g N_A_623_115#_c_1123_n 0.00479454f $X=2.68 $Y=3.235
+ $X2=2.76 $Y2=1.37
cc_533 N_A_32_115#_c_662_n N_A_623_115#_c_1123_n 0.0702347f $X=2.42 $Y=2.285
+ $X2=2.76 $Y2=1.37
cc_534 N_A_32_115#_c_664_n N_A_623_115#_c_1123_n 0.0104545f $X=2.42 $Y=1.37
+ $X2=2.76 $Y2=1.37
cc_535 N_A_32_115#_c_669_n N_A_623_115#_c_1123_n 3.63286e-19 $X=2.33 $Y=1.37
+ $X2=2.76 $Y2=1.37
cc_536 N_A_32_115#_M1002_g N_A_623_115#_c_1183_n 9.13132e-19 $X=2.25 $Y=3.235
+ $X2=2.845 $Y2=2.705
cc_537 N_A_32_115#_M1005_g N_A_623_115#_c_1183_n 0.0096885f $X=2.68 $Y=3.235
+ $X2=2.845 $Y2=2.705
cc_538 N_A_32_115#_c_649_n N_A_623_115#_c_1131_n 0.00776295f $X=2.605 $Y=1.37
+ $X2=2.905 $Y2=1.37
cc_539 N_A_32_115#_c_664_n N_A_623_115#_c_1131_n 0.00134369f $X=2.42 $Y=1.37
+ $X2=2.905 $Y2=1.37
cc_540 N_A_32_115#_c_669_n N_A_623_115#_c_1131_n 0.0241863f $X=2.33 $Y=1.37
+ $X2=2.905 $Y2=1.37
cc_541 N_A_243_89#_M1001_g N_A_785_89#_M1023_g 0.04635f $X=3.64 $Y=0.835 $X2=4
+ $Y2=0.835
cc_542 N_A_243_89#_c_775_n N_A_785_89#_c_960_n 0.04635f $X=3.58 $Y=1.74 $X2=4.06
+ $Y2=1.74
cc_543 N_A_243_89#_c_776_n N_A_785_89#_c_960_n 8.11121e-19 $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_544 N_A_243_89#_c_782_n N_A_785_89#_c_960_n 6.38549e-19 $X=4.915 $Y=1.725
+ $X2=4.06 $Y2=1.74
cc_545 N_A_243_89#_c_783_n N_A_785_89#_c_960_n 9.00828e-19 $X=3.725 $Y=1.725
+ $X2=4.06 $Y2=1.74
cc_546 N_A_243_89#_c_784_n N_A_785_89#_c_960_n 4.49351e-19 $X=4.645 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_547 N_A_243_89#_c_785_n N_A_785_89#_c_960_n 0.00295157f $X=4.5 $Y=1.74
+ $X2=4.06 $Y2=1.74
cc_548 N_A_243_89#_c_775_n N_A_785_89#_c_963_n 7.47762e-19 $X=3.58 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_549 N_A_243_89#_c_776_n N_A_785_89#_c_963_n 0.0079274f $X=3.58 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_550 N_A_243_89#_c_777_n N_A_785_89#_c_963_n 0.00183874f $X=4.645 $Y=0.755
+ $X2=4.062 $Y2=1.812
cc_551 N_A_243_89#_c_782_n N_A_785_89#_c_963_n 0.00400058f $X=4.915 $Y=1.725
+ $X2=4.062 $Y2=1.812
cc_552 N_A_243_89#_c_783_n N_A_785_89#_c_963_n 0.00135239f $X=3.725 $Y=1.725
+ $X2=4.062 $Y2=1.812
cc_553 N_A_243_89#_c_784_n N_A_785_89#_c_963_n 0.00102352f $X=4.645 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_554 N_A_243_89#_c_785_n N_A_785_89#_c_963_n 0.0115044f $X=4.5 $Y=1.74
+ $X2=4.062 $Y2=1.812
cc_555 N_A_243_89#_c_775_n N_A_785_89#_c_964_n 5.35826e-19 $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_556 N_A_243_89#_c_776_n N_A_785_89#_c_964_n 6.26362e-19 $X=3.58 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_557 N_A_243_89#_c_782_n N_A_785_89#_c_964_n 2.40837e-19 $X=4.915 $Y=1.725
+ $X2=4.06 $Y2=2.48
cc_558 N_A_243_89#_c_783_n N_A_785_89#_c_964_n 0.00136024f $X=3.725 $Y=1.725
+ $X2=4.06 $Y2=2.48
cc_559 N_A_243_89#_c_784_n N_A_785_89#_c_964_n 0.0012974f $X=4.645 $Y=1.74
+ $X2=4.06 $Y2=2.48
cc_560 N_A_243_89#_c_782_n N_A_785_89#_c_965_n 0.00107657f $X=4.915 $Y=1.725
+ $X2=5.595 $Y2=0.755
cc_561 N_A_243_89#_c_781_n N_A_785_89#_c_968_n 0.0168304f $X=4.915 $Y=2.62
+ $X2=5.595 $Y2=2.955
cc_562 N_A_243_89#_c_782_n N_A_785_89#_c_970_n 0.0038359f $X=4.915 $Y=1.725
+ $X2=5.595 $Y2=1.74
cc_563 N_A_243_89#_c_781_n N_A_785_89#_c_971_n 0.0136501f $X=4.915 $Y=2.62
+ $X2=4.935 $Y2=2.48
cc_564 N_A_243_89#_c_782_n N_A_785_89#_c_971_n 0.0020334f $X=4.915 $Y=1.725
+ $X2=4.935 $Y2=2.48
cc_565 N_A_243_89#_c_797_n N_A_785_89#_c_971_n 0.0134665f $X=4.915 $Y=2.705
+ $X2=4.935 $Y2=2.48
cc_566 N_A_243_89#_c_784_n N_A_785_89#_c_971_n 0.00360662f $X=4.645 $Y=1.74
+ $X2=4.935 $Y2=2.48
cc_567 N_A_243_89#_c_781_n N_A_785_89#_c_973_n 0.0185071f $X=4.915 $Y=2.62
+ $X2=5.007 $Y2=2.395
cc_568 N_A_243_89#_c_782_n N_A_785_89#_c_975_n 0.00779877f $X=4.915 $Y=1.725
+ $X2=5.08 $Y2=1.74
cc_569 N_A_243_89#_c_784_n N_A_785_89#_c_975_n 0.0198607f $X=4.645 $Y=1.74
+ $X2=5.08 $Y2=1.74
cc_570 N_A_243_89#_c_777_n N_A_623_115#_c_1116_n 0.00662411f $X=4.645 $Y=0.755
+ $X2=5.38 $Y2=1.205
cc_571 N_A_243_89#_c_777_n N_A_623_115#_M1021_g 0.00201047f $X=4.645 $Y=0.755
+ $X2=5.38 $Y2=3.235
cc_572 N_A_243_89#_c_792_n N_A_623_115#_M1021_g 0.00781432f $X=4.645 $Y=2.955
+ $X2=5.38 $Y2=3.235
cc_573 N_A_243_89#_c_781_n N_A_623_115#_M1021_g 0.0110692f $X=4.915 $Y=2.62
+ $X2=5.38 $Y2=3.235
cc_574 N_A_243_89#_c_782_n N_A_623_115#_M1021_g 0.00299487f $X=4.915 $Y=1.725
+ $X2=5.38 $Y2=3.235
cc_575 N_A_243_89#_c_797_n N_A_623_115#_M1021_g 0.00340068f $X=4.915 $Y=2.705
+ $X2=5.38 $Y2=3.235
cc_576 N_A_243_89#_c_777_n N_A_623_115#_c_1121_n 0.00361086f $X=4.645 $Y=0.755
+ $X2=5.38 $Y2=1.37
cc_577 N_A_243_89#_c_766_n N_A_623_115#_c_1123_n 0.0122297f $X=2.965 $Y=1.82
+ $X2=2.76 $Y2=1.37
cc_578 N_A_243_89#_c_774_n N_A_623_115#_c_1123_n 0.0112175f $X=3.04 $Y=1.825
+ $X2=2.76 $Y2=1.37
cc_579 N_A_243_89#_M1000_g N_A_623_115#_c_1153_n 0.0162544f $X=3.04 $Y=3.235
+ $X2=3.17 $Y2=2.705
cc_580 N_A_243_89#_c_768_n N_A_623_115#_c_1124_n 0.0013046f $X=3.445 $Y=1.825
+ $X2=3.44 $Y2=1.34
cc_581 N_A_243_89#_M1001_g N_A_623_115#_c_1124_n 0.011734f $X=3.64 $Y=0.835
+ $X2=3.44 $Y2=1.34
cc_582 N_A_243_89#_c_775_n N_A_623_115#_c_1124_n 0.00190498f $X=3.58 $Y=1.74
+ $X2=3.44 $Y2=1.34
cc_583 N_A_243_89#_c_776_n N_A_623_115#_c_1124_n 0.00649516f $X=3.58 $Y=1.74
+ $X2=3.44 $Y2=1.34
cc_584 N_A_243_89#_c_783_n N_A_623_115#_c_1124_n 3.68943e-19 $X=3.725 $Y=1.725
+ $X2=3.44 $Y2=1.34
cc_585 N_A_243_89#_c_777_n N_A_623_115#_c_1125_n 0.00736723f $X=4.645 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_586 N_A_243_89#_c_766_n N_A_623_115#_c_1130_n 0.00156696f $X=2.965 $Y=1.82
+ $X2=3.295 $Y2=1.37
cc_587 N_A_243_89#_c_768_n N_A_623_115#_c_1130_n 0.00252279f $X=3.445 $Y=1.825
+ $X2=3.295 $Y2=1.37
cc_588 N_A_243_89#_c_774_n N_A_623_115#_c_1130_n 5.21392e-19 $X=3.04 $Y=1.825
+ $X2=3.295 $Y2=1.37
cc_589 N_A_243_89#_c_766_n N_A_623_115#_c_1131_n 0.00120486f $X=2.965 $Y=1.82
+ $X2=2.905 $Y2=1.37
cc_590 N_A_243_89#_M1001_g N_A_623_115#_c_1132_n 0.0076805f $X=3.64 $Y=0.835
+ $X2=5.03 $Y2=1.37
cc_591 N_A_243_89#_c_777_n N_A_623_115#_c_1132_n 0.0227582f $X=4.645 $Y=0.755
+ $X2=5.03 $Y2=1.37
cc_592 N_A_243_89#_c_782_n N_A_623_115#_c_1132_n 0.00916047f $X=4.915 $Y=1.725
+ $X2=5.03 $Y2=1.37
cc_593 N_A_243_89#_c_784_n N_A_623_115#_c_1132_n 0.0251703f $X=4.645 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_594 N_A_243_89#_c_785_n N_A_623_115#_c_1132_n 0.0641247f $X=4.5 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_595 N_A_243_89#_M1001_g N_A_623_115#_c_1134_n 0.00331631f $X=3.64 $Y=0.835
+ $X2=3.585 $Y2=1.37
cc_596 N_A_243_89#_c_775_n N_A_623_115#_c_1134_n 6.43748e-19 $X=3.58 $Y=1.74
+ $X2=3.585 $Y2=1.37
cc_597 N_A_243_89#_c_776_n N_A_623_115#_c_1134_n 0.00311003f $X=3.58 $Y=1.74
+ $X2=3.585 $Y2=1.37
cc_598 N_A_243_89#_c_783_n N_A_623_115#_c_1134_n 0.0279665f $X=3.725 $Y=1.725
+ $X2=3.585 $Y2=1.37
cc_599 N_A_243_89#_c_777_n N_A_623_115#_c_1135_n 0.00257549f $X=4.645 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_600 N_A_785_89#_c_965_n N_A_623_115#_c_1116_n 0.0220174f $X=5.595 $Y=0.755
+ $X2=5.38 $Y2=1.205
cc_601 N_A_785_89#_c_955_n N_A_623_115#_M1021_g 0.00462538f $X=6.28 $Y=1.905
+ $X2=5.38 $Y2=3.235
cc_602 N_A_785_89#_c_968_n N_A_623_115#_M1021_g 0.023277f $X=5.595 $Y=2.955
+ $X2=5.38 $Y2=3.235
cc_603 N_A_785_89#_c_970_n N_A_623_115#_M1021_g 0.00244533f $X=5.595 $Y=1.74
+ $X2=5.38 $Y2=3.235
cc_604 N_A_785_89#_c_973_n N_A_623_115#_M1021_g 0.0141612f $X=5.007 $Y=2.395
+ $X2=5.38 $Y2=3.235
cc_605 N_A_785_89#_c_974_n N_A_623_115#_M1021_g 0.0162569f $X=6.08 $Y=1.74
+ $X2=5.38 $Y2=3.235
cc_606 N_A_785_89#_c_975_n N_A_623_115#_c_1121_n 0.00415861f $X=5.08 $Y=1.74
+ $X2=5.38 $Y2=1.37
cc_607 N_A_785_89#_c_965_n N_A_623_115#_c_1125_n 0.0115453f $X=5.595 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_608 N_A_785_89#_c_974_n N_A_623_115#_c_1125_n 7.4919e-19 $X=6.08 $Y=1.74
+ $X2=5.175 $Y2=1.37
cc_609 N_A_785_89#_c_975_n N_A_623_115#_c_1125_n 0.00428868f $X=5.08 $Y=1.74
+ $X2=5.175 $Y2=1.37
cc_610 N_A_785_89#_M1023_g N_A_623_115#_c_1132_n 0.0105151f $X=4 $Y=0.835
+ $X2=5.03 $Y2=1.37
cc_611 N_A_785_89#_c_960_n N_A_623_115#_c_1132_n 7.90759e-19 $X=4.06 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_612 N_A_785_89#_c_963_n N_A_623_115#_c_1132_n 0.00516488f $X=4.062 $Y=1.812
+ $X2=5.03 $Y2=1.37
cc_613 N_A_785_89#_c_975_n N_A_623_115#_c_1132_n 0.00830534f $X=5.08 $Y=1.74
+ $X2=5.03 $Y2=1.37
cc_614 N_A_785_89#_c_965_n N_A_623_115#_c_1135_n 0.00389142f $X=5.595 $Y=0.755
+ $X2=5.175 $Y2=1.37
cc_615 N_A_785_89#_c_975_n N_A_623_115#_c_1135_n 0.0270542f $X=5.08 $Y=1.74
+ $X2=5.175 $Y2=1.37
cc_616 N_A_785_89#_c_955_n N_ON_M1025_g 0.0154305f $X=6.28 $Y=1.905 $X2=6.76
+ $Y2=0.755
cc_617 N_A_785_89#_M1008_g N_ON_M1025_g 0.0253877f $X=6.33 $Y=0.755 $X2=6.76
+ $Y2=0.755
cc_618 N_A_785_89#_c_969_n N_ON_M1025_g 6.55283e-19 $X=6.215 $Y=1.74 $X2=6.76
+ $Y2=0.755
cc_619 N_A_785_89#_c_962_n N_ON_M1020_g 0.0102677f $X=6.305 $Y=2.475 $X2=6.76
+ $Y2=3.445
cc_620 N_A_785_89#_c_986_n N_ON_M1020_g 0.0457815f $X=6.305 $Y=2.625 $X2=6.76
+ $Y2=3.445
cc_621 N_A_785_89#_c_955_n N_ON_c_1240_n 0.0212297f $X=6.28 $Y=1.905 $X2=6.7
+ $Y2=2.015
cc_622 N_A_785_89#_c_955_n N_ON_c_1241_n 0.00188672f $X=6.28 $Y=1.905 $X2=6.115
+ $Y2=0.74
cc_623 N_A_785_89#_M1008_g N_ON_c_1241_n 0.0129631f $X=6.33 $Y=0.755 $X2=6.115
+ $Y2=0.74
cc_624 N_A_785_89#_c_965_n N_ON_c_1241_n 0.0324824f $X=5.595 $Y=0.755 $X2=6.115
+ $Y2=0.74
cc_625 N_A_785_89#_c_955_n N_ON_c_1244_n 0.00289364f $X=6.28 $Y=1.905 $X2=6.115
+ $Y2=2.195
cc_626 N_A_785_89#_c_968_n N_ON_c_1244_n 0.00525727f $X=5.595 $Y=2.955 $X2=6.115
+ $Y2=2.195
cc_627 N_A_785_89#_c_969_n N_ON_c_1244_n 0.0101349f $X=6.215 $Y=1.74 $X2=6.115
+ $Y2=2.195
cc_628 N_A_785_89#_c_976_n N_ON_c_1244_n 3.37612e-19 $X=6.215 $Y=1.74 $X2=6.115
+ $Y2=2.195
cc_629 N_A_785_89#_M1006_g N_ON_c_1245_n 0.0241057f $X=6.33 $Y=3.445 $X2=6.115
+ $Y2=3.615
cc_630 N_A_785_89#_c_962_n N_ON_c_1245_n 0.0176611f $X=6.305 $Y=2.475 $X2=6.115
+ $Y2=3.615
cc_631 N_A_785_89#_c_968_n N_ON_c_1245_n 0.0727346f $X=5.595 $Y=2.955 $X2=6.115
+ $Y2=3.615
cc_632 N_A_785_89#_c_955_n N_ON_c_1246_n 0.0192889f $X=6.28 $Y=1.905 $X2=6.615
+ $Y2=1.4
cc_633 N_A_785_89#_c_969_n N_ON_c_1246_n 0.0110497f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=1.4
cc_634 N_A_785_89#_c_976_n N_ON_c_1246_n 0.00387586f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=1.4
cc_635 N_A_785_89#_c_955_n N_ON_c_1248_n 0.00308111f $X=6.28 $Y=1.905 $X2=6.2
+ $Y2=1.4
cc_636 N_A_785_89#_c_965_n N_ON_c_1248_n 0.00869401f $X=5.595 $Y=0.755 $X2=6.2
+ $Y2=1.4
cc_637 N_A_785_89#_c_969_n N_ON_c_1248_n 0.0120752f $X=6.215 $Y=1.74 $X2=6.2
+ $Y2=1.4
cc_638 N_A_785_89#_c_974_n N_ON_c_1248_n 0.00132729f $X=6.08 $Y=1.74 $X2=6.2
+ $Y2=1.4
cc_639 N_A_785_89#_c_976_n N_ON_c_1248_n 0.00306734f $X=6.215 $Y=1.74 $X2=6.2
+ $Y2=1.4
cc_640 N_A_785_89#_c_955_n N_ON_c_1249_n 2.65797e-19 $X=6.28 $Y=1.905 $X2=6.615
+ $Y2=2.11
cc_641 N_A_785_89#_c_962_n N_ON_c_1249_n 0.0142383f $X=6.305 $Y=2.475 $X2=6.615
+ $Y2=2.11
cc_642 N_A_785_89#_c_986_n N_ON_c_1249_n 0.00184481f $X=6.305 $Y=2.625 $X2=6.615
+ $Y2=2.11
cc_643 N_A_785_89#_c_969_n N_ON_c_1249_n 0.00957265f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=2.11
cc_644 N_A_785_89#_c_976_n N_ON_c_1249_n 0.00261089f $X=6.215 $Y=1.74 $X2=6.615
+ $Y2=2.11
cc_645 N_A_785_89#_c_955_n N_ON_c_1250_n 0.00380215f $X=6.28 $Y=1.905 $X2=6.702
+ $Y2=1.658
cc_646 N_A_785_89#_c_969_n N_ON_c_1250_n 0.00996181f $X=6.215 $Y=1.74 $X2=6.702
+ $Y2=1.658
cc_647 N_A_785_89#_c_976_n N_ON_c_1250_n 0.00251327f $X=6.215 $Y=1.74 $X2=6.702
+ $Y2=1.658
cc_648 N_A_785_89#_c_955_n N_ON_c_1251_n 0.00152939f $X=6.28 $Y=1.905 $X2=6.7
+ $Y2=2.015
cc_649 N_A_785_89#_c_976_n N_ON_c_1251_n 0.00137139f $X=6.215 $Y=1.74 $X2=6.7
+ $Y2=2.015
cc_650 N_A_785_89#_c_955_n ON 0.00197254f $X=6.28 $Y=1.905 $X2=6.115 $Y2=2.11
cc_651 N_A_785_89#_c_962_n ON 0.00400769f $X=6.305 $Y=2.475 $X2=6.115 $Y2=2.11
cc_652 N_A_785_89#_c_968_n ON 0.00761812f $X=5.595 $Y=2.955 $X2=6.115 $Y2=2.11
cc_653 N_A_785_89#_c_969_n ON 0.00222181f $X=6.215 $Y=1.74 $X2=6.115 $Y2=2.11
cc_654 N_A_785_89#_c_974_n ON 0.0192933f $X=6.08 $Y=1.74 $X2=6.115 $Y2=2.11
cc_655 N_A_785_89#_c_976_n ON 0.0183431f $X=6.215 $Y=1.74 $X2=6.115 $Y2=2.11
cc_656 N_A_785_89#_c_962_n Q 5.37537e-19 $X=6.305 $Y=2.475 $X2=6.97 $Y2=2.48
cc_657 N_A_785_89#_c_986_n Q 6.11581e-19 $X=6.305 $Y=2.625 $X2=6.97 $Y2=2.48
cc_658 N_A_623_115#_c_1153_n A_551_521# 0.00342591f $X=3.17 $Y=2.705 $X2=2.755
+ $Y2=2.605
cc_659 N_A_623_115#_c_1183_n A_551_521# 0.00144354f $X=2.845 $Y=2.705 $X2=2.755
+ $Y2=2.605
cc_660 N_ON_M1025_g N_Q_c_1317_n 0.00192093f $X=6.76 $Y=0.755 $X2=6.975 $Y2=0.74
cc_661 N_ON_M1025_g N_Q_c_1319_n 0.0301628f $X=6.76 $Y=0.755 $X2=7.09 $Y2=2.395
cc_662 N_ON_c_1246_n N_Q_c_1319_n 0.0113726f $X=6.615 $Y=1.4 $X2=7.09 $Y2=2.395
cc_663 N_ON_c_1249_n N_Q_c_1319_n 0.0111434f $X=6.615 $Y=2.11 $X2=7.09 $Y2=2.395
cc_664 N_ON_c_1250_n N_Q_c_1319_n 0.0155777f $X=6.702 $Y=1.658 $X2=7.09
+ $Y2=2.395
cc_665 N_ON_c_1251_n N_Q_c_1319_n 0.0164341f $X=6.7 $Y=2.015 $X2=7.09 $Y2=2.395
cc_666 N_ON_M1020_g N_Q_c_1320_n 0.00583168f $X=6.76 $Y=3.445 $X2=7.09 $Y2=2.48
cc_667 N_ON_M1020_g N_Q_c_1327_n 0.0206543f $X=6.76 $Y=3.445 $X2=6.972 $Y2=2.88
cc_668 N_ON_M1025_g N_Q_c_1321_n 0.00695117f $X=6.76 $Y=0.755 $X2=7.09 $Y2=1.07
cc_669 N_ON_M1020_g Q 0.0140617f $X=6.76 $Y=3.445 $X2=6.97 $Y2=2.48
cc_670 N_ON_c_1245_n Q 0.00550321f $X=6.115 $Y=3.615 $X2=6.97 $Y2=2.48
cc_671 N_ON_c_1249_n Q 0.00287022f $X=6.615 $Y=2.11 $X2=6.97 $Y2=2.48
