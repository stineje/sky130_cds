magic
tech sky130A
magscale 1 2
timestamp 1606864575
<< checkpaint >>
rect -1269 -242 1459 2379
rect -1209 -1243 1345 -242
<< nwell >>
rect -9 529 199 1119
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1049 85 1083
<< locali >>
rect 0 1089 198 1110
rect 0 1049 51 1089
rect 85 1049 198 1089
rect 35 483 69 965
rect 121 589 155 1049
rect 31 449 47 483
rect 81 449 97 483
rect 35 365 69 449
rect 35 331 155 365
rect 35 115 69 331
rect 121 115 155 331
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 47 449 81 483
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1089 198 1110
rect 0 1055 51 1089
rect 85 1055 198 1089
rect 0 1049 198 1055
rect 35 483 108 489
rect 35 449 47 483
rect 81 449 108 483
rect 35 443 108 449
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel viali 64 466 64 466 1 A
port 1 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
