* File: sky130_osu_sc_12T_ls__or2_l.pex.spice
* Created: Fri Nov 12 15:40:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__OR2_L%GND 1 2 21 25 27 35 42 44 47
r36 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r37 33 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r38 33 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.74
r39 27 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r40 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r41 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r42 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r43 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r44 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r45 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r46 2 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.74
r47 1 25 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OR2_L%VDD 1 13 15 24 28 30 33
r21 30 33 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r22 22 28 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r23 22 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=3.615
r24 20 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r25 17 20 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r26 15 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r27 15 20 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r28 13 20 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r29 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r30 1 24 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=3.025 $X2=1.12 $Y2=3.615
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OR2_L%B 3 7 12 15 21
r30 15 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.48
r31 15 18 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.48
+ $X2=0.27 $Y2=2.565
r32 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.565 $X2=0.27 $Y2=2.565
r33 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.565
+ $X2=0.475 $Y2=2.565
r34 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.73
+ $X2=0.475 $Y2=2.565
r35 5 7 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=0.475 $Y=2.73
+ $X2=0.475 $Y2=3.445
r36 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.4
+ $X2=0.475 $Y2=2.565
r37 1 3 843.5 $w=1.5e-07 $l=1.645e-06 $layer=POLY_cond $X=0.475 $Y=2.4 $X2=0.475
+ $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OR2_L%A 3 7 10 14 20
c42 10 0 7.14041e-20 $X=0.95 $Y=2.275
c43 7 0 3.10762e-20 $X=0.905 $Y=3.445
r44 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.48
+ $X2=0.95 $Y2=2.48
r45 14 17 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.95 $Y=2.275
+ $X2=0.95 $Y2=2.48
r46 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.275 $X2=0.95 $Y2=2.275
r47 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.275
+ $X2=0.95 $Y2=2.44
r48 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.275
+ $X2=0.95 $Y2=2.11
r49 7 12 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=0.905 $Y=3.445
+ $X2=0.905 $Y2=2.44
r50 3 11 694.798 $w=1.5e-07 $l=1.355e-06 $layer=POLY_cond $X=0.905 $Y=0.755
+ $X2=0.905 $Y2=2.11
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OR2_L%A_27_605# 1 3 11 15 17 19 20 25 27 28 30
+ 33 37 39
r74 35 39 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.825
+ $X2=0.65 $Y2=1.825
r75 35 37 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.825
+ $X2=1.43 $Y2=1.825
r76 31 39 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.74
+ $X2=0.65 $Y2=1.825
r77 31 33 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=0.69 $Y=1.74 $X2=0.69
+ $Y2=0.74
r78 29 39 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=1.91
+ $X2=0.65 $Y2=1.825
r79 29 30 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.61 $Y=1.91
+ $X2=0.61 $Y2=2.935
r80 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.02
+ $X2=0.61 $Y2=2.935
r81 27 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.02
+ $X2=0.345 $Y2=3.02
r82 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.105
+ $X2=0.345 $Y2=3.02
r83 23 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.26 $Y=3.105
+ $X2=0.26 $Y2=3.615
r84 22 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.825 $X2=1.43 $Y2=1.825
r85 19 20 49.8721 $w=1.85e-07 $l=1.35e-07 $layer=POLY_cond $X=1.352 $Y=2.7
+ $X2=1.352 $Y2=2.835
r86 17 22 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=1.99
+ $X2=1.412 $Y2=1.825
r87 17 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.99
+ $X2=1.37 $Y2=2.7
r88 15 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.335 $Y=3.445
+ $X2=1.335 $Y2=2.835
r89 9 22 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.66
+ $X2=1.412 $Y2=1.825
r90 9 11 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.335 $Y=1.66
+ $X2=1.335 $Y2=0.755
r91 3 25 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.615
r92 1 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__OR2_L%Y 1 3 10 16 24 27 30
c34 30 0 1.0248e-19 $X=1.55 $Y=2.48
r35 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.48
r36 22 24 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.11
r37 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.485
+ $X2=1.55 $Y2=1.37
r38 21 24 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.485
+ $X2=1.55 $Y2=2.11
r39 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.48
r40 16 19 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=3.615
r41 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.37
+ $X2=1.55 $Y2=1.37
r42 10 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.37
r43 3 19 600 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=3.025 $X2=1.55 $Y2=3.615
r44 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

