* File: sky130_osu_sc_15T_ls__tielo.pxi.spice
* Created: Fri Nov 12 15:00:19 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__TIELO%GND N_GND_M1001_s N_GND_M1001_b N_GND_c_2_p
+ N_GND_c_3_p GND PM_SKY130_OSU_SC_15T_LS__TIELO%GND
x_PM_SKY130_OSU_SC_15T_LS__TIELO%VDD N_VDD_M1000_s N_VDD_M1000_b N_VDD_c_12_p
+ N_VDD_c_13_p VDD PM_SKY130_OSU_SC_15T_LS__TIELO%VDD
x_PM_SKY130_OSU_SC_15T_LS__TIELO%A_80_89# N_A_80_89#_M1000_d N_A_80_89#_M1001_g
+ N_A_80_89#_M1000_g N_A_80_89#_c_22_n N_A_80_89#_c_23_n N_A_80_89#_c_24_n
+ PM_SKY130_OSU_SC_15T_LS__TIELO%A_80_89#
x_PM_SKY130_OSU_SC_15T_LS__TIELO%Y N_Y_M1001_d N_Y_c_38_n Y
+ PM_SKY130_OSU_SC_15T_LS__TIELO%Y
cc_1 N_GND_M1001_b N_A_80_89#_M1001_g 0.114871f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=0.945
cc_2 N_GND_c_2_p N_A_80_89#_M1001_g 0.00866533f $X=0.26 $Y=0.865 $X2=0.475
+ $Y2=0.945
cc_3 N_GND_c_3_p N_A_80_89#_M1001_g 0.00468827f $X=0.34 $Y=0.19 $X2=0.475
+ $Y2=0.945
cc_4 N_GND_M1001_b N_A_80_89#_M1000_g 0.00665813f $X=-0.045 $Y=0 $X2=0.475
+ $Y2=3.825
cc_5 N_GND_M1001_b N_A_80_89#_c_22_n 0.0423935f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.4
cc_6 N_GND_M1001_b N_A_80_89#_c_23_n 0.00652005f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=3.205
cc_7 N_GND_M1001_b N_A_80_89#_c_24_n 0.0167595f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.4
cc_8 N_GND_M1001_b N_Y_c_38_n 0.024976f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.865
cc_9 N_GND_c_3_p N_Y_c_38_n 0.00476261f $X=0.34 $Y=0.19 $X2=0.69 $Y2=0.865
cc_10 N_GND_M1001_b Y 0.0182702f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.59
cc_11 N_VDD_M1000_b N_A_80_89#_M1000_g 0.0303814f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_12 N_VDD_c_12_p N_A_80_89#_M1000_g 0.00751602f $X=0.26 $Y=3.205 $X2=0.475
+ $Y2=3.825
cc_13 N_VDD_c_13_p N_A_80_89#_M1000_g 0.00496961f $X=0.34 $Y=5.36 $X2=0.475
+ $Y2=3.825
cc_14 VDD N_A_80_89#_M1000_g 0.00429146f $X=0.34 $Y=5.31 $X2=0.475 $Y2=3.825
cc_15 N_VDD_M1000_b N_A_80_89#_c_23_n 0.0103047f $X=-0.045 $Y=2.645 $X2=0.69
+ $Y2=3.205
cc_16 N_VDD_c_13_p N_A_80_89#_c_23_n 0.00477009f $X=0.34 $Y=5.36 $X2=0.69
+ $Y2=3.205
cc_17 VDD N_A_80_89#_c_23_n 0.00435496f $X=0.34 $Y=5.31 $X2=0.69 $Y2=3.205
cc_18 N_A_80_89#_M1001_g N_Y_c_38_n 0.019532f $X=0.475 $Y=0.945 $X2=0.69
+ $Y2=0.865
cc_19 N_A_80_89#_c_22_n N_Y_c_38_n 0.001024f $X=0.535 $Y=2.4 $X2=0.69 $Y2=0.865
cc_20 N_A_80_89#_c_24_n N_Y_c_38_n 0.00263908f $X=0.69 $Y=2.4 $X2=0.69 $Y2=0.865
cc_21 N_A_80_89#_M1001_g Y 0.0167084f $X=0.475 $Y=0.945 $X2=0.69 $Y2=1.59
cc_22 N_A_80_89#_c_22_n Y 0.00251432f $X=0.535 $Y=2.4 $X2=0.69 $Y2=1.59
cc_23 N_A_80_89#_c_24_n Y 0.00701253f $X=0.69 $Y=2.4 $X2=0.69 $Y2=1.59
