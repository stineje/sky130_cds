* File: sky130_osu_sc_15T_hs__xnor2_l.pxi.spice
* Created: Fri Nov 12 14:34:04 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%GND N_GND_M1003_d N_GND_M1008_d N_GND_M1003_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_9_p N_GND_c_51_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_15T_HS__XNOR2_L%GND
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%VDD N_VDD_M1005_d N_VDD_M1011_d N_VDD_M1005_b
+ N_VDD_c_76_p N_VDD_c_77_p N_VDD_c_73_p N_VDD_c_91_p N_VDD_c_93_p VDD
+ N_VDD_c_74_p PM_SKY130_OSU_SC_15T_HS__XNOR2_L%VDD
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%A N_A_M1003_g N_A_M1005_g N_A_c_116_n
+ N_A_M1001_g N_A_M1009_g N_A_c_123_n N_A_c_124_n N_A_c_125_n N_A_c_126_n
+ N_A_c_127_n N_A_c_128_n N_A_c_131_n N_A_c_132_n N_A_c_133_n N_A_c_134_n A
+ N_A_c_137_n PM_SKY130_OSU_SC_15T_HS__XNOR2_L%A
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1005_s N_A_27_115#_M1002_g N_A_27_115#_M1007_g
+ N_A_27_115#_c_231_n N_A_27_115#_c_232_n N_A_27_115#_c_233_n
+ N_A_27_115#_c_236_n N_A_27_115#_c_237_n N_A_27_115#_c_238_n
+ N_A_27_115#_c_239_n PM_SKY130_OSU_SC_15T_HS__XNOR2_L%A_27_115#
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%A_238_89# N_A_238_89#_M1004_d
+ N_A_238_89#_M1006_d N_A_238_89#_M1010_g N_A_238_89#_M1000_g
+ N_A_238_89#_c_308_n N_A_238_89#_c_309_n N_A_238_89#_c_310_n
+ N_A_238_89#_c_312_n N_A_238_89#_c_313_n
+ PM_SKY130_OSU_SC_15T_HS__XNOR2_L%A_238_89#
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%B N_B_M1008_g N_B_c_382_n N_B_M1011_g
+ N_B_c_369_n N_B_c_370_n N_B_M1004_g N_B_c_374_n N_B_c_389_n N_B_M1006_g
+ N_B_c_375_n N_B_c_377_n N_B_c_378_n B PM_SKY130_OSU_SC_15T_HS__XNOR2_L%B
x_PM_SKY130_OSU_SC_15T_HS__XNOR2_L%Y N_Y_M1010_d N_Y_M1000_d N_Y_c_422_n
+ N_Y_c_423_n N_Y_c_454_n N_Y_c_428_n N_Y_c_438_n Y N_Y_c_427_n N_Y_c_432_n
+ PM_SKY130_OSU_SC_15T_HS__XNOR2_L%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.0237592f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_A_M1003_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_A_M1003_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.895
cc_4 N_GND_c_4_p N_A_M1003_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=0.895
cc_5 N_GND_M1003_b N_A_c_116_n 0.00577419f $X=-0.045 $Y=0 $X2=0.71 $Y2=1.465
cc_6 N_GND_c_3_p N_A_c_116_n 0.0033834f $X=0.69 $Y=0.74 $X2=0.71 $Y2=1.465
cc_7 N_GND_M1003_b N_A_M1001_g 0.0175294f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.895
cc_8 N_GND_c_3_p N_A_M1001_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.895
cc_9 N_GND_c_9_p N_A_M1001_g 0.00606474f $X=2.355 $Y=0.152 $X2=0.905 $Y2=0.895
cc_10 N_GND_c_4_p N_A_M1001_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.905 $Y2=0.895
cc_11 N_GND_M1003_b N_A_M1009_g 0.0214281f $X=-0.045 $Y=0 $X2=1.865 $Y2=3.825
cc_12 N_GND_M1003_b N_A_c_123_n 0.00962022f $X=-0.045 $Y=0 $X2=0.45 $Y2=1.465
cc_13 N_GND_M1003_b N_A_c_124_n 0.0608283f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.6
cc_14 N_GND_M1003_b N_A_c_125_n 0.00432809f $X=-0.045 $Y=0 $X2=0.45 $Y2=2.75
cc_15 N_GND_M1003_b N_A_c_126_n 0.0240171f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.465
cc_16 N_GND_M1003_b N_A_c_127_n 0.052624f $X=-0.045 $Y=0 $X2=1.865 $Y2=2.145
cc_17 N_GND_M1003_d N_A_c_128_n 8.79072e-19 $X=0.55 $Y=0.575 $X2=0.845 $Y2=1.22
cc_18 N_GND_M1003_b N_A_c_128_n 0.00255856f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.22
cc_19 N_GND_c_3_p N_A_c_128_n 6.39251e-19 $X=0.69 $Y=0.74 $X2=0.845 $Y2=1.22
cc_20 N_GND_M1003_b N_A_c_131_n 0.0106735f $X=-0.045 $Y=0 $X2=2.145 $Y2=1.22
cc_21 N_GND_M1003_b N_A_c_132_n 0.00276199f $X=-0.045 $Y=0 $X2=2.225 $Y2=2.13
cc_22 N_GND_M1003_b N_A_c_133_n 0.0134259f $X=-0.045 $Y=0 $X2=2 $Y2=1.22
cc_23 N_GND_M1003_d N_A_c_134_n 0.00408434f $X=0.55 $Y=0.575 $X2=0.99 $Y2=1.22
cc_24 N_GND_M1003_b N_A_c_134_n 0.00274472f $X=-0.045 $Y=0 $X2=0.99 $Y2=1.22
cc_25 N_GND_c_3_p N_A_c_134_n 0.0036198f $X=0.69 $Y=0.74 $X2=0.99 $Y2=1.22
cc_26 N_GND_M1003_b N_A_c_137_n 0.00259705f $X=-0.045 $Y=0 $X2=2.145 $Y2=1.22
cc_27 N_GND_M1003_b N_A_27_115#_M1002_g 0.0184711f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=3.825
cc_28 N_GND_M1003_b N_A_27_115#_M1007_g 0.0222165f $X=-0.045 $Y=0 $X2=1.865
+ $Y2=0.895
cc_29 N_GND_c_9_p N_A_27_115#_M1007_g 0.00606474f $X=2.355 $Y=0.152 $X2=1.865
+ $Y2=0.895
cc_30 N_GND_c_4_p N_A_27_115#_M1007_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.865
+ $Y2=0.895
cc_31 N_GND_M1003_b N_A_27_115#_c_231_n 0.0277923f $X=-0.045 $Y=0 $X2=0.845
+ $Y2=2.13
cc_32 N_GND_M1003_b N_A_27_115#_c_232_n 0.0362346f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.59
cc_33 N_GND_M1003_b N_A_27_115#_c_233_n 0.0407947f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_34 N_GND_c_2_p N_A_27_115#_c_233_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_35 N_GND_c_4_p N_A_27_115#_c_233_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_36 N_GND_M1003_b N_A_27_115#_c_236_n 0.0201658f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.205
cc_37 N_GND_M1003_b N_A_27_115#_c_237_n 0.0354732f $X=-0.045 $Y=0 $X2=1.68
+ $Y2=2.13
cc_38 N_GND_M1003_b N_A_27_115#_c_238_n 0.00497247f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.59
cc_39 N_GND_M1003_b N_A_27_115#_c_239_n 0.00692367f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.13
cc_40 N_GND_M1003_b N_A_238_89#_M1010_g 0.0751109f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=0.895
cc_41 N_GND_c_9_p N_A_238_89#_M1010_g 0.00606474f $X=2.355 $Y=0.152 $X2=1.265
+ $Y2=0.895
cc_42 N_GND_c_4_p N_A_238_89#_M1010_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.265
+ $Y2=0.895
cc_43 N_GND_M1003_b N_A_238_89#_c_308_n 0.021482f $X=-0.045 $Y=0 $X2=1.325
+ $Y2=2.505
cc_44 N_GND_M1003_b N_A_238_89#_c_309_n 0.0330247f $X=-0.045 $Y=0 $X2=2.785
+ $Y2=2.505
cc_45 N_GND_M1003_b N_A_238_89#_c_310_n 0.0660509f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=0.865
cc_46 N_GND_c_4_p N_A_238_89#_c_310_n 0.00476261f $X=2.38 $Y=0.19 $X2=2.87
+ $Y2=0.865
cc_47 N_GND_M1003_b N_A_238_89#_c_312_n 0.00243339f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=3.205
cc_48 N_GND_M1003_b N_A_238_89#_c_313_n 0.00720662f $X=-0.045 $Y=0 $X2=2.87
+ $Y2=2.505
cc_49 N_GND_M1003_b N_B_M1008_g 0.0178481f $X=-0.045 $Y=0 $X2=2.225 $Y2=0.895
cc_50 N_GND_c_9_p N_B_M1008_g 0.00606474f $X=2.355 $Y=0.152 $X2=2.225 $Y2=0.895
cc_51 N_GND_c_51_p N_B_M1008_g 0.00308284f $X=2.44 $Y=0.74 $X2=2.225 $Y2=0.895
cc_52 N_GND_c_4_p N_B_M1008_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.225 $Y2=0.895
cc_53 N_GND_M1003_b N_B_c_369_n 0.00761231f $X=-0.045 $Y=0 $X2=2.58 $Y2=2.675
cc_54 N_GND_M1003_b N_B_c_370_n 0.00457156f $X=-0.045 $Y=0 $X2=2.3 $Y2=2.675
cc_55 N_GND_M1003_b N_B_M1004_g 0.0298422f $X=-0.045 $Y=0 $X2=2.655 $Y2=0.895
cc_56 N_GND_c_51_p N_B_M1004_g 0.00308284f $X=2.44 $Y=0.74 $X2=2.655 $Y2=0.895
cc_57 N_GND_c_4_p N_B_M1004_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.655 $Y2=0.895
cc_58 N_GND_M1003_b N_B_c_374_n 0.0472661f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.6
cc_59 N_GND_M1003_b N_B_c_375_n 0.0457888f $X=-0.045 $Y=0 $X2=2.655 $Y2=1.572
cc_60 N_GND_c_51_p N_B_c_375_n 0.0026533f $X=2.44 $Y=0.74 $X2=2.655 $Y2=1.572
cc_61 N_GND_M1003_b N_B_c_377_n 0.00181559f $X=-0.045 $Y=0 $X2=2.655 $Y2=2.675
cc_62 N_GND_M1003_b N_B_c_378_n 0.00227638f $X=-0.045 $Y=0 $X2=2.53 $Y2=1.59
cc_63 N_GND_c_51_p N_B_c_378_n 0.00210748f $X=2.44 $Y=0.74 $X2=2.53 $Y2=1.59
cc_64 N_GND_M1003_b B 0.00236483f $X=-0.045 $Y=0 $X2=2.53 $Y2=1.59
cc_65 N_GND_c_51_p B 0.00356087f $X=2.44 $Y=0.74 $X2=2.53 $Y2=1.59
cc_66 N_GND_M1003_b N_Y_c_422_n 0.00998803f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.59
cc_67 N_GND_M1003_b N_Y_c_423_n 0.00313365f $X=-0.045 $Y=0 $X2=1.565 $Y2=0.865
cc_68 N_GND_c_9_p N_Y_c_423_n 0.0148236f $X=2.355 $Y=0.152 $X2=1.565 $Y2=0.865
cc_69 N_GND_c_4_p N_Y_c_423_n 0.00954899f $X=2.38 $Y=0.19 $X2=1.565 $Y2=0.865
cc_70 N_GND_M1003_b Y 0.00698114f $X=-0.045 $Y=0 $X2=1.42 $Y2=1.875
cc_71 N_GND_M1003_b N_Y_c_427_n 0.00238374f $X=-0.045 $Y=0 $X2=1.425 $Y2=1.59
cc_72 N_VDD_M1005_b N_A_M1009_g 0.0219053f $X=-0.045 $Y=2.645 $X2=1.865
+ $Y2=3.825
cc_73 N_VDD_c_73_p N_A_M1009_g 0.00496961f $X=2.355 $Y=5.397 $X2=1.865 $Y2=3.825
cc_74 N_VDD_c_74_p N_A_M1009_g 0.00429146f $X=2.38 $Y=5.36 $X2=1.865 $Y2=3.825
cc_75 N_VDD_M1005_b N_A_c_125_n 0.0283712f $X=-0.045 $Y=2.645 $X2=0.45 $Y2=2.75
cc_76 N_VDD_c_76_p N_A_c_125_n 0.00496961f $X=0.605 $Y=5.397 $X2=0.45 $Y2=2.75
cc_77 N_VDD_c_77_p N_A_c_125_n 0.00362996f $X=0.69 $Y=3.205 $X2=0.45 $Y2=2.75
cc_78 N_VDD_c_74_p N_A_c_125_n 0.00429146f $X=2.38 $Y=5.36 $X2=0.45 $Y2=2.75
cc_79 N_VDD_M1005_b N_A_27_115#_M1002_g 0.0201514f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_80 N_VDD_c_77_p N_A_27_115#_M1002_g 0.00362996f $X=0.69 $Y=3.205 $X2=0.905
+ $Y2=3.825
cc_81 N_VDD_c_73_p N_A_27_115#_M1002_g 0.00496961f $X=2.355 $Y=5.397 $X2=0.905
+ $Y2=3.825
cc_82 N_VDD_c_74_p N_A_27_115#_M1002_g 0.00429146f $X=2.38 $Y=5.36 $X2=0.905
+ $Y2=3.825
cc_83 N_VDD_c_77_p N_A_27_115#_c_231_n 0.0017177f $X=0.69 $Y=3.205 $X2=0.845
+ $Y2=2.13
cc_84 N_VDD_M1005_b N_A_27_115#_c_236_n 0.0109193f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.205
cc_85 N_VDD_c_76_p N_A_27_115#_c_236_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=3.205
cc_86 N_VDD_c_74_p N_A_27_115#_c_236_n 0.00435496f $X=2.38 $Y=5.36 $X2=0.26
+ $Y2=3.205
cc_87 N_VDD_M1005_b N_A_238_89#_M1000_g 0.0196878f $X=-0.045 $Y=2.645 $X2=1.265
+ $Y2=3.825
cc_88 N_VDD_c_73_p N_A_238_89#_M1000_g 0.00496961f $X=2.355 $Y=5.397 $X2=1.265
+ $Y2=3.825
cc_89 N_VDD_c_74_p N_A_238_89#_M1000_g 0.00429146f $X=2.38 $Y=5.36 $X2=1.265
+ $Y2=3.825
cc_90 N_VDD_M1005_b N_A_238_89#_c_308_n 0.00559382f $X=-0.045 $Y=2.645 $X2=1.325
+ $Y2=2.505
cc_91 N_VDD_c_91_p N_A_238_89#_c_309_n 0.00811678f $X=2.44 $Y=3.205 $X2=2.785
+ $Y2=2.505
cc_92 N_VDD_M1005_b N_A_238_89#_c_312_n 0.0103574f $X=-0.045 $Y=2.645 $X2=2.87
+ $Y2=3.205
cc_93 N_VDD_c_93_p N_A_238_89#_c_312_n 0.00477009f $X=2.38 $Y=5.36 $X2=2.87
+ $Y2=3.205
cc_94 N_VDD_c_74_p N_A_238_89#_c_312_n 0.00435496f $X=2.38 $Y=5.36 $X2=2.87
+ $Y2=3.205
cc_95 N_VDD_M1005_b N_B_c_382_n 0.01436f $X=-0.045 $Y=2.645 $X2=2.225 $Y2=2.75
cc_96 N_VDD_c_73_p N_B_c_382_n 0.00496961f $X=2.355 $Y=5.397 $X2=2.225 $Y2=2.75
cc_97 N_VDD_c_91_p N_B_c_382_n 0.00362996f $X=2.44 $Y=3.205 $X2=2.225 $Y2=2.75
cc_98 N_VDD_c_74_p N_B_c_382_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.225 $Y2=2.75
cc_99 N_VDD_M1005_b N_B_c_369_n 0.00535962f $X=-0.045 $Y=2.645 $X2=2.58
+ $Y2=2.675
cc_100 N_VDD_c_91_p N_B_c_369_n 0.00221017f $X=2.44 $Y=3.205 $X2=2.58 $Y2=2.675
cc_101 N_VDD_M1005_b N_B_c_370_n 0.00345657f $X=-0.045 $Y=2.645 $X2=2.3
+ $Y2=2.675
cc_102 N_VDD_M1005_b N_B_c_389_n 0.0187201f $X=-0.045 $Y=2.645 $X2=2.655
+ $Y2=2.75
cc_103 N_VDD_c_91_p N_B_c_389_n 0.00362996f $X=2.44 $Y=3.205 $X2=2.655 $Y2=2.75
cc_104 N_VDD_c_93_p N_B_c_389_n 0.00496961f $X=2.38 $Y=5.36 $X2=2.655 $Y2=2.75
cc_105 N_VDD_c_74_p N_B_c_389_n 0.00429146f $X=2.38 $Y=5.36 $X2=2.655 $Y2=2.75
cc_106 N_VDD_M1005_b N_B_c_377_n 0.00423637f $X=-0.045 $Y=2.645 $X2=2.655
+ $Y2=2.675
cc_107 N_VDD_M1005_b N_Y_c_428_n 0.00402069f $X=-0.045 $Y=2.645 $X2=1.565
+ $Y2=3.205
cc_108 N_VDD_c_73_p N_Y_c_428_n 0.00925108f $X=2.355 $Y=5.397 $X2=1.565
+ $Y2=3.205
cc_109 N_VDD_c_74_p N_Y_c_428_n 0.00876183f $X=2.38 $Y=5.36 $X2=1.565 $Y2=3.205
cc_110 N_VDD_M1005_b Y 0.00321849f $X=-0.045 $Y=2.645 $X2=1.42 $Y2=1.875
cc_111 N_VDD_c_77_p N_Y_c_432_n 0.0045586f $X=0.69 $Y=3.205 $X2=1.425 $Y2=3.07
cc_112 N_A_c_124_n N_A_27_115#_M1002_g 0.0111858f $X=0.45 $Y=2.6 $X2=0.905
+ $Y2=3.825
cc_113 N_A_c_125_n N_A_27_115#_M1002_g 0.0252253f $X=0.45 $Y=2.75 $X2=0.905
+ $Y2=3.825
cc_114 N_A_c_131_n N_A_27_115#_M1007_g 0.00311835f $X=2.145 $Y=1.22 $X2=1.865
+ $Y2=0.895
cc_115 N_A_c_133_n N_A_27_115#_M1007_g 0.0134125f $X=2 $Y=1.22 $X2=1.865
+ $Y2=0.895
cc_116 N_A_c_137_n N_A_27_115#_M1007_g 9.56269e-19 $X=2.145 $Y=1.22 $X2=1.865
+ $Y2=0.895
cc_117 N_A_c_124_n N_A_27_115#_c_231_n 0.0212638f $X=0.45 $Y=2.6 $X2=0.845
+ $Y2=2.13
cc_118 N_A_c_126_n N_A_27_115#_c_231_n 0.0184269f $X=0.845 $Y=1.465 $X2=0.845
+ $Y2=2.13
cc_119 N_A_c_128_n N_A_27_115#_c_231_n 6.74966e-19 $X=0.845 $Y=1.22 $X2=0.845
+ $Y2=2.13
cc_120 N_A_c_134_n N_A_27_115#_c_231_n 4.48459e-19 $X=0.99 $Y=1.22 $X2=0.845
+ $Y2=2.13
cc_121 N_A_c_127_n N_A_27_115#_c_232_n 0.00515091f $X=1.865 $Y=2.145 $X2=1.765
+ $Y2=1.59
cc_122 N_A_c_131_n N_A_27_115#_c_232_n 0.00194908f $X=2.145 $Y=1.22 $X2=1.765
+ $Y2=1.59
cc_123 N_A_c_133_n N_A_27_115#_c_232_n 0.00130191f $X=2 $Y=1.22 $X2=1.765
+ $Y2=1.59
cc_124 N_A_M1003_g N_A_27_115#_c_233_n 0.00917829f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=0.865
cc_125 N_A_c_123_n N_A_27_115#_c_233_n 0.022872f $X=0.45 $Y=1.465 $X2=0.26
+ $Y2=0.865
cc_126 N_A_c_128_n N_A_27_115#_c_233_n 0.0197497f $X=0.845 $Y=1.22 $X2=0.26
+ $Y2=0.865
cc_127 N_A_c_134_n N_A_27_115#_c_233_n 0.00710152f $X=0.99 $Y=1.22 $X2=0.26
+ $Y2=0.865
cc_128 N_A_c_124_n N_A_27_115#_c_236_n 0.0221084f $X=0.45 $Y=2.6 $X2=0.26
+ $Y2=3.205
cc_129 N_A_c_125_n N_A_27_115#_c_236_n 0.00766083f $X=0.45 $Y=2.75 $X2=0.26
+ $Y2=3.205
cc_130 N_A_c_116_n N_A_27_115#_c_237_n 8.76512e-19 $X=0.71 $Y=1.465 $X2=1.68
+ $Y2=2.13
cc_131 N_A_c_124_n N_A_27_115#_c_237_n 0.0199699f $X=0.45 $Y=2.6 $X2=1.68
+ $Y2=2.13
cc_132 N_A_c_125_n N_A_27_115#_c_237_n 0.00165231f $X=0.45 $Y=2.75 $X2=1.68
+ $Y2=2.13
cc_133 N_A_c_126_n N_A_27_115#_c_237_n 8.34298e-19 $X=0.845 $Y=1.465 $X2=1.68
+ $Y2=2.13
cc_134 N_A_c_127_n N_A_27_115#_c_237_n 0.00528869f $X=1.865 $Y=2.145 $X2=1.68
+ $Y2=2.13
cc_135 N_A_c_128_n N_A_27_115#_c_237_n 0.00826927f $X=0.845 $Y=1.22 $X2=1.68
+ $Y2=2.13
cc_136 N_A_c_132_n N_A_27_115#_c_237_n 0.0116688f $X=2.225 $Y=2.13 $X2=1.68
+ $Y2=2.13
cc_137 N_A_c_127_n N_A_27_115#_c_238_n 5.00447e-19 $X=1.865 $Y=2.145 $X2=1.765
+ $Y2=1.59
cc_138 N_A_c_131_n N_A_27_115#_c_238_n 0.0360591f $X=2.145 $Y=1.22 $X2=1.765
+ $Y2=1.59
cc_139 N_A_c_133_n N_A_27_115#_c_238_n 0.00737704f $X=2 $Y=1.22 $X2=1.765
+ $Y2=1.59
cc_140 N_A_M1001_g N_A_238_89#_M1010_g 0.0806795f $X=0.905 $Y=0.895 $X2=1.265
+ $Y2=0.895
cc_141 N_A_c_124_n N_A_238_89#_M1010_g 0.00462097f $X=0.45 $Y=2.6 $X2=1.265
+ $Y2=0.895
cc_142 N_A_c_127_n N_A_238_89#_M1010_g 0.00525031f $X=1.865 $Y=2.145 $X2=1.265
+ $Y2=0.895
cc_143 N_A_c_128_n N_A_238_89#_M1010_g 0.00228168f $X=0.845 $Y=1.22 $X2=1.265
+ $Y2=0.895
cc_144 N_A_c_133_n N_A_238_89#_M1010_g 0.0133678f $X=2 $Y=1.22 $X2=1.265
+ $Y2=0.895
cc_145 N_A_c_134_n N_A_238_89#_M1010_g 8.6716e-19 $X=0.99 $Y=1.22 $X2=1.265
+ $Y2=0.895
cc_146 N_A_M1009_g N_A_238_89#_M1000_g 0.0446488f $X=1.865 $Y=3.825 $X2=1.265
+ $Y2=3.825
cc_147 N_A_M1009_g N_A_238_89#_c_308_n 0.0126871f $X=1.865 $Y=3.825 $X2=1.325
+ $Y2=2.505
cc_148 N_A_M1009_g N_A_238_89#_c_309_n 0.018341f $X=1.865 $Y=3.825 $X2=2.785
+ $Y2=2.505
cc_149 N_A_c_127_n N_A_238_89#_c_309_n 0.00796541f $X=1.865 $Y=2.145 $X2=2.785
+ $Y2=2.505
cc_150 N_A_c_132_n N_A_238_89#_c_309_n 0.0206305f $X=2.225 $Y=2.13 $X2=2.785
+ $Y2=2.505
cc_151 N_A_c_131_n N_A_238_89#_c_310_n 0.0141947f $X=2.145 $Y=1.22 $X2=2.87
+ $Y2=0.865
cc_152 N_A_c_132_n N_A_238_89#_c_310_n 0.00742262f $X=2.225 $Y=2.13 $X2=2.87
+ $Y2=0.865
cc_153 N_A_c_137_n N_A_238_89#_c_310_n 0.00547471f $X=2.145 $Y=1.22 $X2=2.87
+ $Y2=0.865
cc_154 N_A_c_131_n N_B_M1008_g 0.00753906f $X=2.145 $Y=1.22 $X2=2.225 $Y2=0.895
cc_155 N_A_c_137_n N_B_M1008_g 0.00991486f $X=2.145 $Y=1.22 $X2=2.225 $Y2=0.895
cc_156 N_A_M1009_g N_B_c_370_n 0.141103f $X=1.865 $Y=3.825 $X2=2.3 $Y2=2.675
cc_157 N_A_c_127_n N_B_c_370_n 0.00779298f $X=1.865 $Y=2.145 $X2=2.3 $Y2=2.675
cc_158 N_A_c_131_n N_B_M1004_g 0.00106222f $X=2.145 $Y=1.22 $X2=2.655 $Y2=0.895
cc_159 N_A_c_137_n N_B_M1004_g 0.00122438f $X=2.145 $Y=1.22 $X2=2.655 $Y2=0.895
cc_160 N_A_M1009_g N_B_c_374_n 0.00402444f $X=1.865 $Y=3.825 $X2=2.655 $Y2=2.6
cc_161 N_A_c_127_n N_B_c_374_n 0.0193201f $X=1.865 $Y=2.145 $X2=2.655 $Y2=2.6
cc_162 N_A_c_131_n N_B_c_374_n 0.00243832f $X=2.145 $Y=1.22 $X2=2.655 $Y2=2.6
cc_163 N_A_c_132_n N_B_c_374_n 0.00131152f $X=2.225 $Y=2.13 $X2=2.655 $Y2=2.6
cc_164 N_A_c_127_n N_B_c_375_n 0.00620704f $X=1.865 $Y=2.145 $X2=2.655 $Y2=1.572
cc_165 N_A_c_131_n N_B_c_375_n 0.00728935f $X=2.145 $Y=1.22 $X2=2.655 $Y2=1.572
cc_166 N_A_c_132_n N_B_c_375_n 0.00132282f $X=2.225 $Y=2.13 $X2=2.655 $Y2=1.572
cc_167 N_A_c_131_n N_B_c_378_n 0.0165474f $X=2.145 $Y=1.22 $X2=2.53 $Y2=1.59
cc_168 N_A_c_127_n B 0.00116112f $X=1.865 $Y=2.145 $X2=2.53 $Y2=1.59
cc_169 N_A_c_131_n B 0.007568f $X=2.145 $Y=1.22 $X2=2.53 $Y2=1.59
cc_170 N_A_c_132_n B 0.00408329f $X=2.225 $Y=2.13 $X2=2.53 $Y2=1.59
cc_171 N_A_c_137_n B 0.00136805f $X=2.145 $Y=1.22 $X2=2.53 $Y2=1.59
cc_172 N_A_c_133_n N_Y_M1010_d 0.00209203f $X=2 $Y=1.22 $X2=1.34 $Y2=0.575
cc_173 N_A_c_131_n N_Y_c_422_n 0.00631055f $X=2.145 $Y=1.22 $X2=1.425 $Y2=1.59
cc_174 N_A_c_133_n N_Y_c_422_n 0.0115606f $X=2 $Y=1.22 $X2=1.425 $Y2=1.59
cc_175 N_A_c_134_n N_Y_c_422_n 7.8621e-19 $X=0.99 $Y=1.22 $X2=1.425 $Y2=1.59
cc_176 N_A_c_137_n N_Y_c_422_n 7.10974e-19 $X=2.145 $Y=1.22 $X2=1.425 $Y2=1.59
cc_177 N_A_c_128_n N_Y_c_438_n 0.0143881f $X=0.845 $Y=1.22 $X2=1.537 $Y2=1.155
cc_178 N_A_c_131_n N_Y_c_438_n 5.37889e-19 $X=2.145 $Y=1.22 $X2=1.537 $Y2=1.155
cc_179 N_A_c_133_n N_Y_c_438_n 0.0271638f $X=2 $Y=1.22 $X2=1.537 $Y2=1.155
cc_180 N_A_c_134_n N_Y_c_438_n 0.00133183f $X=0.99 $Y=1.22 $X2=1.537 $Y2=1.155
cc_181 N_A_c_137_n N_Y_c_438_n 0.00144576f $X=2.145 $Y=1.22 $X2=1.537 $Y2=1.155
cc_182 N_A_c_126_n Y 2.24638e-19 $X=0.845 $Y=1.465 $X2=1.42 $Y2=1.875
cc_183 N_A_c_127_n Y 0.00743805f $X=1.865 $Y=2.145 $X2=1.42 $Y2=1.875
cc_184 N_A_c_128_n Y 0.00146257f $X=0.845 $Y=1.22 $X2=1.42 $Y2=1.875
cc_185 N_A_c_132_n Y 6.70937e-19 $X=2.225 $Y=2.13 $X2=1.42 $Y2=1.875
cc_186 N_A_c_126_n N_Y_c_427_n 0.0011785f $X=0.845 $Y=1.465 $X2=1.425 $Y2=1.59
cc_187 N_A_c_128_n N_Y_c_427_n 0.00531647f $X=0.845 $Y=1.22 $X2=1.425 $Y2=1.59
cc_188 N_A_c_133_n N_Y_c_427_n 0.0259642f $X=2 $Y=1.22 $X2=1.425 $Y2=1.59
cc_189 N_A_c_133_n A_196_115# 0.0077095f $X=2 $Y=1.22 $X2=0.98 $Y2=0.575
cc_190 N_A_c_134_n A_196_115# 7.14422e-19 $X=0.99 $Y=1.22 $X2=0.98 $Y2=0.575
cc_191 N_A_c_131_n A_388_115# 0.00143201f $X=2.145 $Y=1.22 $X2=1.94 $Y2=0.575
cc_192 N_A_c_133_n A_388_115# 0.00228573f $X=2 $Y=1.22 $X2=1.94 $Y2=0.575
cc_193 N_A_c_137_n A_388_115# 0.00626365f $X=2.145 $Y=1.22 $X2=1.94 $Y2=0.575
cc_194 N_A_27_115#_M1007_g N_A_238_89#_M1010_g 0.0208808f $X=1.865 $Y=0.895
+ $X2=1.265 $Y2=0.895
cc_195 N_A_27_115#_c_231_n N_A_238_89#_M1010_g 0.0904081f $X=0.845 $Y=2.13
+ $X2=1.265 $Y2=0.895
cc_196 N_A_27_115#_c_232_n N_A_238_89#_M1010_g 0.0141925f $X=1.765 $Y=1.59
+ $X2=1.265 $Y2=0.895
cc_197 N_A_27_115#_c_237_n N_A_238_89#_M1010_g 0.0146245f $X=1.68 $Y=2.13
+ $X2=1.265 $Y2=0.895
cc_198 N_A_27_115#_c_238_n N_A_238_89#_M1010_g 0.00755502f $X=1.765 $Y=1.59
+ $X2=1.265 $Y2=0.895
cc_199 N_A_27_115#_M1002_g N_A_238_89#_c_308_n 0.0904081f $X=0.905 $Y=3.825
+ $X2=1.325 $Y2=2.505
cc_200 N_A_27_115#_c_237_n N_A_238_89#_c_308_n 0.00220335f $X=1.68 $Y=2.13
+ $X2=1.325 $Y2=2.505
cc_201 N_A_27_115#_M1002_g N_A_238_89#_c_309_n 0.00444529f $X=0.905 $Y=3.825
+ $X2=2.785 $Y2=2.505
cc_202 N_A_27_115#_c_232_n N_A_238_89#_c_309_n 6.30959e-19 $X=1.765 $Y=1.59
+ $X2=2.785 $Y2=2.505
cc_203 N_A_27_115#_c_237_n N_A_238_89#_c_309_n 0.0436145f $X=1.68 $Y=2.13
+ $X2=2.785 $Y2=2.505
cc_204 N_A_27_115#_M1007_g N_B_M1008_g 0.0335733f $X=1.865 $Y=0.895 $X2=2.225
+ $Y2=0.895
cc_205 N_A_27_115#_c_232_n N_B_c_375_n 0.0379418f $X=1.765 $Y=1.59 $X2=2.655
+ $Y2=1.572
cc_206 N_A_27_115#_M1007_g N_Y_c_422_n 0.00208671f $X=1.865 $Y=0.895 $X2=1.425
+ $Y2=1.59
cc_207 N_A_27_115#_c_232_n N_Y_c_422_n 0.00161977f $X=1.765 $Y=1.59 $X2=1.425
+ $Y2=1.59
cc_208 N_A_27_115#_c_237_n N_Y_c_422_n 0.00556015f $X=1.68 $Y=2.13 $X2=1.425
+ $Y2=1.59
cc_209 N_A_27_115#_c_238_n N_Y_c_422_n 0.0159901f $X=1.765 $Y=1.59 $X2=1.425
+ $Y2=1.59
cc_210 N_A_27_115#_M1002_g N_Y_c_454_n 7.92921e-19 $X=0.905 $Y=3.825 $X2=1.565
+ $Y2=3.185
cc_211 N_A_27_115#_M1007_g N_Y_c_438_n 0.00368227f $X=1.865 $Y=0.895 $X2=1.537
+ $Y2=1.155
cc_212 N_A_27_115#_c_232_n N_Y_c_438_n 0.00192667f $X=1.765 $Y=1.59 $X2=1.537
+ $Y2=1.155
cc_213 N_A_27_115#_c_238_n N_Y_c_438_n 0.00214495f $X=1.765 $Y=1.59 $X2=1.537
+ $Y2=1.155
cc_214 N_A_27_115#_M1002_g Y 0.00191867f $X=0.905 $Y=3.825 $X2=1.42 $Y2=1.875
cc_215 N_A_27_115#_c_231_n Y 9.27207e-19 $X=0.845 $Y=2.13 $X2=1.42 $Y2=1.875
cc_216 N_A_27_115#_c_232_n Y 7.0267e-19 $X=1.765 $Y=1.59 $X2=1.42 $Y2=1.875
cc_217 N_A_27_115#_c_237_n Y 0.0160336f $X=1.68 $Y=2.13 $X2=1.42 $Y2=1.875
cc_218 N_A_27_115#_c_238_n Y 0.015499f $X=1.765 $Y=1.59 $X2=1.42 $Y2=1.875
cc_219 N_A_27_115#_c_232_n N_Y_c_427_n 0.00394131f $X=1.765 $Y=1.59 $X2=1.425
+ $Y2=1.59
cc_220 N_A_27_115#_c_237_n N_Y_c_427_n 0.00440188f $X=1.68 $Y=2.13 $X2=1.425
+ $Y2=1.59
cc_221 N_A_27_115#_c_238_n N_Y_c_427_n 0.00746221f $X=1.765 $Y=1.59 $X2=1.425
+ $Y2=1.59
cc_222 N_A_27_115#_M1002_g N_Y_c_432_n 0.00108503f $X=0.905 $Y=3.825 $X2=1.425
+ $Y2=3.07
cc_223 N_A_238_89#_c_309_n N_B_c_370_n 0.0133212f $X=2.785 $Y=2.505 $X2=2.3
+ $Y2=2.675
cc_224 N_A_238_89#_c_310_n N_B_M1004_g 0.0401968f $X=2.87 $Y=0.865 $X2=2.655
+ $Y2=0.895
cc_225 N_A_238_89#_c_309_n N_B_c_374_n 0.020054f $X=2.785 $Y=2.505 $X2=2.655
+ $Y2=2.6
cc_226 N_A_238_89#_c_312_n N_B_c_374_n 0.0149444f $X=2.87 $Y=3.205 $X2=2.655
+ $Y2=2.6
cc_227 N_A_238_89#_c_309_n N_B_c_375_n 0.00180943f $X=2.785 $Y=2.505 $X2=2.655
+ $Y2=1.572
cc_228 N_A_238_89#_c_309_n N_B_c_378_n 0.00433845f $X=2.785 $Y=2.505 $X2=2.53
+ $Y2=1.59
cc_229 N_A_238_89#_c_310_n N_B_c_378_n 0.0214571f $X=2.87 $Y=0.865 $X2=2.53
+ $Y2=1.59
cc_230 N_A_238_89#_c_310_n B 0.00642833f $X=2.87 $Y=0.865 $X2=2.53 $Y2=1.59
cc_231 N_A_238_89#_M1000_g N_Y_c_454_n 0.0034761f $X=1.265 $Y=3.825 $X2=1.565
+ $Y2=3.185
cc_232 N_A_238_89#_c_308_n N_Y_c_454_n 0.00170549f $X=1.325 $Y=2.505 $X2=1.565
+ $Y2=3.185
cc_233 N_A_238_89#_c_309_n N_Y_c_454_n 0.015078f $X=2.785 $Y=2.505 $X2=1.565
+ $Y2=3.185
cc_234 N_A_238_89#_M1010_g N_Y_c_438_n 0.00718079f $X=1.265 $Y=0.895 $X2=1.537
+ $Y2=1.155
cc_235 N_A_238_89#_M1010_g Y 0.00982251f $X=1.265 $Y=0.895 $X2=1.42 $Y2=1.875
cc_236 N_A_238_89#_M1000_g Y 0.00464698f $X=1.265 $Y=3.825 $X2=1.42 $Y2=1.875
cc_237 N_A_238_89#_c_308_n Y 0.00651733f $X=1.325 $Y=2.505 $X2=1.42 $Y2=1.875
cc_238 N_A_238_89#_c_309_n Y 0.0165306f $X=2.785 $Y=2.505 $X2=1.42 $Y2=1.875
cc_239 N_A_238_89#_M1010_g N_Y_c_427_n 0.00425916f $X=1.265 $Y=0.895 $X2=1.425
+ $Y2=1.59
cc_240 N_A_238_89#_M1000_g N_Y_c_432_n 0.00624758f $X=1.265 $Y=3.825 $X2=1.425
+ $Y2=3.07
cc_241 N_A_238_89#_c_309_n N_Y_c_432_n 0.00233457f $X=2.785 $Y=2.505 $X2=1.425
+ $Y2=3.07
