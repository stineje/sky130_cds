* File: sky130_osu_sc_12T_hs__dffsr_1.pex.spice
* Created: Fri Nov 12 15:09:47 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%GND 1 2 3 4 5 6 7 8 9 127 131 133 140
+ 142 152 154 158 160 170 172 182 184 191 193 203 205 212 238 240
c265 191 0 1.63226e-19 $X=7.47 $Y=0.755
c266 182 0 3.34232e-19 $X=6.52 $Y=0.755
c267 158 0 3.07651e-19 $X=3.02 $Y=0.755
c268 152 0 2.98797e-19 $X=2.5 $Y=0.755
c269 127 0 2.70767e-19 $X=-0.05 $Y=0
r270 238 240 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.855 $Y2=0.152
r271 214 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=0.152
+ $X2=9.71 $Y2=0.152
r272 210 234 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.152
r273 210 212 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.71 $Y=0.305
+ $X2=9.71 $Y2=0.755
r274 206 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.152
+ $X2=8.75 $Y2=0.152
r275 205 234 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=0.152
+ $X2=9.71 $Y2=0.152
r276 201 233 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.152
r277 201 203 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.75 $Y=0.305
+ $X2=8.75 $Y2=0.74
r278 194 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.152
+ $X2=7.47 $Y2=0.152
r279 193 233 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.152
+ $X2=8.75 $Y2=0.152
r280 189 232 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.152
r281 189 191 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.47 $Y=0.305
+ $X2=7.47 $Y2=0.755
r282 184 232 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=0.152
+ $X2=7.47 $Y2=0.152
r283 180 182 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.52 $Y=0.305
+ $X2=6.52 $Y2=0.755
r284 173 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.152
+ $X2=4.77 $Y2=0.152
r285 168 228 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.152
r286 168 170 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.77 $Y=0.305
+ $X2=4.77 $Y2=0.74
r287 160 228 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.152
+ $X2=4.77 $Y2=0.152
r288 156 158 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.02 $Y=0.305
+ $X2=3.02 $Y2=0.755
r289 155 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.152
+ $X2=2.5 $Y2=0.152
r290 154 155 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=2.935 $Y=0.152
+ $X2=2.585 $Y2=0.152
r291 150 224 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.152
r292 150 152 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.5 $Y=0.305
+ $X2=2.5 $Y2=0.755
r293 143 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0.152
+ $X2=1.22 $Y2=0.152
r294 142 224 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.152
+ $X2=2.5 $Y2=0.152
r295 138 223 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.152
r296 138 140 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.22 $Y=0.305
+ $X2=1.22 $Y2=0.74
r297 133 223 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.152
+ $X2=1.22 $Y2=0.152
r298 129 131 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r299 127 240 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=0.19
+ $X2=9.855 $Y2=0.19
r300 127 238 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r301 127 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.52 $Y2=0.305
r302 127 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.435 $Y2=0.152
r303 127 185 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.152
+ $X2=6.605 $Y2=0.152
r304 127 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.02 $Y2=0.305
r305 127 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=2.935 $Y2=0.152
r306 127 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.152
+ $X2=3.105 $Y2=0.152
r307 127 129 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r308 127 134 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r309 127 214 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.855 $Y=0.152
+ $X2=9.795 $Y2=0.152
r310 127 205 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=9.625 $Y2=0.152
r311 127 206 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.835 $Y2=0.152
r312 127 193 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.665 $Y2=0.152
r313 127 194 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=7.815 $Y=0.152
+ $X2=7.555 $Y2=0.152
r314 127 184 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.385 $Y2=0.152
r315 127 185 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.605 $Y2=0.152
r316 127 172 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.435 $Y2=0.152
r317 127 173 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.855 $Y2=0.152
r318 127 160 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=4.685 $Y2=0.152
r319 127 161 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.105 $Y2=0.152
r320 127 142 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.415 $Y2=0.152
r321 127 143 14.7362 $w=3.03e-07 $l=3.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.305 $Y2=0.152
r322 127 133 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.135 $Y2=0.152
r323 127 134 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r324 9 212 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.57
+ $Y=0.575 $X2=9.71 $Y2=0.755
r325 8 203 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.61
+ $Y=0.575 $X2=8.75 $Y2=0.74
r326 7 191 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.755
r327 6 182 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.755
r328 5 170 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.575 $X2=4.77 $Y2=0.74
r329 4 158 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.575 $X2=3.02 $Y2=0.755
r330 3 152 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.575 $X2=2.5 $Y2=0.755
r331 2 140 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.575 $X2=1.22 $Y2=0.74
r332 1 131 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%VDD 1 2 3 4 5 6 7 89 93 95 103 105 111
+ 113 121 123 131 133 139 141 149 155 170 174
c165 149 0 1.98165e-19 $X=9.71 $Y=2.955
r166 170 174 4.43367 $w=3.05e-07 $l=9.52e-06 $layer=MET1_cond $X=0.335 $Y=4.287
+ $X2=9.855 $Y2=4.287
r167 158 170 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.335 $Y=4.25
+ $X2=0.335 $Y2=4.25
r168 155 174 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=9.855 $Y=4.25
+ $X2=9.855 $Y2=4.25
r169 153 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=4.287
+ $X2=9.71 $Y2=4.287
r170 153 155 2.4 $w=3.05e-07 $l=6e-08 $layer=LI1_cond $X=9.795 $Y=4.287
+ $X2=9.855 $Y2=4.287
r171 149 152 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.71 $Y=2.955
+ $X2=9.71 $Y2=3.635
r172 147 168 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.71 $Y=4.135
+ $X2=9.71 $Y2=4.287
r173 147 152 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.71 $Y=4.135
+ $X2=9.71 $Y2=3.635
r174 144 146 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=8.495 $Y=4.287
+ $X2=9.175 $Y2=4.287
r175 142 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=4.287
+ $X2=7.9 $Y2=4.287
r176 142 144 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=7.985 $Y=4.287
+ $X2=8.495 $Y2=4.287
r177 141 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.625 $Y=4.287
+ $X2=9.71 $Y2=4.287
r178 141 146 17.0033 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=9.625 $Y=4.287
+ $X2=9.175 $Y2=4.287
r179 137 167 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=4.287
r180 137 139 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=4.135
+ $X2=7.9 $Y2=3.7
r181 134 165 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=4.287
+ $X2=6.52 $Y2=4.287
r182 134 136 20.0261 $w=3.03e-07 $l=5.3e-07 $layer=LI1_cond $X=6.605 $Y=4.287
+ $X2=7.135 $Y2=4.287
r183 133 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=4.287
+ $X2=7.9 $Y2=4.287
r184 133 136 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=4.287
+ $X2=7.135 $Y2=4.287
r185 129 165 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.52 $Y=4.135
+ $X2=6.52 $Y2=4.287
r186 129 131 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.52 $Y=4.135
+ $X2=6.52 $Y2=3.21
r187 126 128 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=4.287
+ $X2=5.775 $Y2=4.287
r188 124 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=4.287
+ $X2=4.77 $Y2=4.287
r189 124 126 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=4.855 $Y=4.287
+ $X2=5.095 $Y2=4.287
r190 123 165 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=4.287
+ $X2=6.52 $Y2=4.287
r191 123 128 24.9381 $w=3.03e-07 $l=6.6e-07 $layer=LI1_cond $X=6.435 $Y=4.287
+ $X2=5.775 $Y2=4.287
r192 119 163 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.77 $Y=4.135
+ $X2=4.77 $Y2=4.287
r193 119 121 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.77 $Y=4.135
+ $X2=4.77 $Y2=3.295
r194 116 118 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=4.287
+ $X2=4.415 $Y2=4.287
r195 114 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=4.287
+ $X2=3.02 $Y2=4.287
r196 114 116 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=3.105 $Y=4.287
+ $X2=3.735 $Y2=4.287
r197 113 163 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=4.287
+ $X2=4.77 $Y2=4.287
r198 113 118 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=4.685 $Y=4.287
+ $X2=4.415 $Y2=4.287
r199 109 162 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.02 $Y=4.135
+ $X2=3.02 $Y2=4.287
r200 109 111 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.02 $Y=4.135
+ $X2=3.02 $Y2=3.295
r201 106 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=4.287
+ $X2=2.07 $Y2=4.287
r202 106 108 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.155 $Y=4.287
+ $X2=2.375 $Y2=4.287
r203 105 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=4.287
+ $X2=3.02 $Y2=4.287
r204 105 108 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=2.935 $Y=4.287
+ $X2=2.375 $Y2=4.287
r205 101 160 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.07 $Y=4.135
+ $X2=2.07 $Y2=4.287
r206 101 103 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=4.135
+ $X2=2.07 $Y2=3.7
r207 98 100 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=4.287
+ $X2=1.695 $Y2=4.287
r208 96 158 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r209 96 98 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.015 $Y2=4.287
r210 95 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=4.287
+ $X2=2.07 $Y2=4.287
r211 95 100 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.985 $Y=4.287
+ $X2=1.695 $Y2=4.287
r212 91 158 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r213 91 93 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r214 89 155 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=9.65 $Y=4.135 $X2=9.855 $Y2=4.22
r215 89 146 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=4.135 $X2=9.175 $Y2=4.22
r216 89 144 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=4.135 $X2=8.495 $Y2=4.22
r217 89 167 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=4.135 $X2=7.815 $Y2=4.22
r218 89 136 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=4.135 $X2=7.135 $Y2=4.22
r219 89 165 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=4.135 $X2=6.455 $Y2=4.22
r220 89 128 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=4.135 $X2=5.775 $Y2=4.22
r221 89 126 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=4.135 $X2=5.095 $Y2=4.22
r222 89 118 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=4.135 $X2=4.415 $Y2=4.22
r223 89 116 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=4.135 $X2=3.735 $Y2=4.22
r224 89 162 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=4.135 $X2=3.055 $Y2=4.22
r225 89 108 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=4.135 $X2=2.375 $Y2=4.22
r226 89 100 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=4.135 $X2=1.695 $Y2=4.22
r227 89 98 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=4.135 $X2=1.015 $Y2=4.22
r228 89 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=4.135 $X2=0.335 $Y2=4.22
r229 7 152 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=9.57
+ $Y=2.605 $X2=9.71 $Y2=3.635
r230 7 149 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=9.57
+ $Y=2.605 $X2=9.71 $Y2=2.955
r231 6 139 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.605 $X2=7.9 $Y2=3.7
r232 5 131 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=3.21
r233 4 121 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=4.63
+ $Y=2.605 $X2=4.77 $Y2=3.295
r234 3 111 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.605 $X2=3.02 $Y2=3.295
r235 2 103 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.605 $X2=2.07 $Y2=3.7
r236 1 93 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%RN 3 5 7 13 15 21
c42 21 0 7.48684e-20 $X=0.325 $Y=2.85
c43 3 0 1.41286e-20 $X=0.475 $Y=0.85
r44 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=2.85
+ $X2=0.325 $Y2=2.85
r45 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.53 $Y2=1.825
r46 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r47 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=1.99
+ $X2=0.32 $Y2=1.825
r48 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=1.99 $X2=0.32
+ $Y2=2.85
r49 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.825 $X2=0.53 $Y2=1.825
r50 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.53 $Y2=1.825
r51 5 7 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=3.235
r52 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.53 $Y2=1.825
r53 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.475 $Y2=0.85
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_110_115# 1 3 10 13 15 17 18 20 23 26
+ 29 33 36 39 43 47 54 55 57 64 67 71 72 73 77 80 81
c230 77 0 1.63455e-19 $X=0.87 $Y=1.37
c231 71 0 1.41286e-20 $X=0.87 $Y=1.255
c232 67 0 3.77772e-20 $X=8.86 $Y=1.27
c233 64 0 7.48684e-20 $X=0.87 $Y=2.26
c234 57 0 1.98452e-19 $X=1.23 $Y=1.27
c235 39 0 1.09867e-19 $X=8.545 $Y=2.27
c236 26 0 8.31638e-20 $X=8.8 $Y=2.125
r237 80 81 0.0806629 $w=2.95e-07 $l=1.15e-07 $layer=MET1_cond $X=8.862 $Y=1.37
+ $X2=8.862 $Y2=1.255
r238 74 81 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=8.86 $Y=1.085
+ $X2=8.86 $Y2=1.255
r239 72 74 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=8.775 $Y=1
+ $X2=8.86 $Y2=1.085
r240 72 73 7.52974 $w=1.7e-07 $l=7.82e-06 $layer=MET1_cond $X=8.775 $Y=1
+ $X2=0.955 $Y2=1
r241 71 77 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.87 $Y=1.255
+ $X2=0.87 $Y2=1.37
r242 70 73 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.87 $Y=1.085
+ $X2=0.955 $Y2=1
r243 70 71 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=0.87 $Y=1.085
+ $X2=0.87 $Y2=1.255
r244 69 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.86 $Y=1.37
+ $X2=8.86 $Y2=1.37
r245 67 69 4.51852 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=8.86 $Y=1.27 $X2=8.86
+ $Y2=1.37
r246 62 64 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.26
+ $X2=0.87 $Y2=2.26
r247 59 61 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.27
+ $X2=0.87 $Y2=1.27
r248 55 61 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.27
+ $X2=0.87 $Y2=1.27
r249 55 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.955 $Y=1.27
+ $X2=1.23 $Y2=1.27
r250 54 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.87 $Y=1.37
+ $X2=0.87 $Y2=1.37
r251 52 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=2.26
r252 52 54 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=1.37
r253 51 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.355
+ $X2=0.87 $Y2=1.27
r254 51 54 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.87 $Y=1.355
+ $X2=0.87 $Y2=1.37
r255 47 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r256 45 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.26
r257 45 47 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.955
r258 41 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.185
+ $X2=0.69 $Y2=1.27
r259 41 43 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.69 $Y=1.185
+ $X2=0.69 $Y2=0.755
r260 39 40 60.25 $w=2.04e-07 $l=2.55e-07 $layer=POLY_cond $X=8.545 $Y=2.27
+ $X2=8.8 $Y2=2.27
r261 38 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.86
+ $Y=1.27 $X2=8.86 $Y2=1.27
r262 36 38 12.05 $w=2.4e-07 $l=6e-08 $layer=POLY_cond $X=8.8 $Y=1.27 $X2=8.86
+ $Y2=1.27
r263 32 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.27 $X2=1.23 $Y2=1.27
r264 32 33 10.7111 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=1.23 $Y=1.27 $X2=1.29
+ $Y2=1.27
r265 27 29 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.29 $Y=2.395
+ $X2=1.425 $Y2=2.395
r266 26 40 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.8 $Y=2.125
+ $X2=8.8 $Y2=2.27
r267 25 36 13.7767 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=1.435
+ $X2=8.8 $Y2=1.27
r268 25 26 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.8 $Y=1.435
+ $X2=8.8 $Y2=2.125
r269 21 39 10.0333 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.545 $Y=2.415
+ $X2=8.545 $Y2=2.27
r270 21 23 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.545 $Y=2.415
+ $X2=8.545 $Y2=3.235
r271 18 36 53.2208 $w=2.4e-07 $l=3.37565e-07 $layer=POLY_cond $X=8.535 $Y=1.105
+ $X2=8.8 $Y2=1.27
r272 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.535 $Y=1.105
+ $X2=8.535 $Y2=0.785
r273 15 33 25.8852 $w=2.7e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.435 $Y=1.105
+ $X2=1.29 $Y2=1.27
r274 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.435 $Y=1.105
+ $X2=1.435 $Y2=0.785
r275 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=2.47
+ $X2=1.425 $Y2=2.395
r276 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.425 $Y=2.47
+ $X2=1.425 $Y2=3.235
r277 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=2.32
+ $X2=1.29 $Y2=2.395
r278 9 33 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.435
+ $X2=1.29 $Y2=1.27
r279 9 10 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=1.29 $Y=1.435
+ $X2=1.29 $Y2=2.32
r280 3 49 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r281 3 47 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r282 1 43 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%SN 1 2 5 9 13 17 22 25 29 32 34 37 39
+ 45 47 48 49 56
c193 48 0 1.36413e-19 $X=7.79 $Y=2.85
c194 29 0 1.5152e-19 $X=1.71 $Y=2.62
c195 2 0 1.95862e-19 $X=1.89 $Y=1.785
c196 1 0 1.98452e-19 $X=1.89 $Y=1.405
r197 54 56 0.00223214 $w=2.8e-07 $l=5e-09 $layer=MET1_cond $X=7.935 $Y=2.802
+ $X2=7.94 $Y2=2.802
r198 49 51 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=2.195 $Y=2.85
+ $X2=2.055 $Y2=2.85
r199 48 54 0.0838839 $w=2.8e-07 $l=1.67287e-07 $layer=MET1_cond $X=7.79 $Y=2.85
+ $X2=7.935 $Y2=2.802
r200 48 49 5.38733 $w=1.7e-07 $l=5.595e-06 $layer=MET1_cond $X=7.79 $Y=2.85
+ $X2=2.195 $Y2=2.85
r201 42 45 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=1.815
+ $X2=8.02 $Y2=1.815
r202 41 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.055 $Y=2.85
+ $X2=2.055 $Y2=2.85
r203 39 41 17.9872 $w=2.34e-07 $l=3.45e-07 $layer=LI1_cond $X=1.71 $Y=2.777
+ $X2=2.055 $Y2=2.777
r204 34 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.935 $Y=2.845
+ $X2=7.935 $Y2=2.845
r205 32 47 5.51377 $w=1.73e-07 $l=8.7e-08 $layer=LI1_cond $X=7.937 $Y=2.482
+ $X2=7.937 $Y2=2.395
r206 32 34 23.0057 $w=1.73e-07 $l=3.63e-07 $layer=LI1_cond $X=7.937 $Y=2.482
+ $X2=7.937 $Y2=2.845
r207 30 42 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=1.94
+ $X2=7.935 $Y2=1.815
r208 30 47 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=7.935 $Y=1.94
+ $X2=7.935 $Y2=2.395
r209 29 39 2.60974 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.71 $Y=2.62
+ $X2=1.71 $Y2=2.777
r210 28 37 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=1.95
r211 28 29 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=2.62
r212 25 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.02
+ $Y=1.775 $X2=8.02 $Y2=1.775
r213 25 27 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=8.032 $Y=1.775
+ $X2=8.032 $Y2=1.94
r214 25 26 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=8.032 $Y=1.775
+ $X2=8.032 $Y2=1.61
r215 22 23 5.53115 $w=3.05e-07 $l=3.5e-08 $layer=POLY_cond $X=1.855 $Y=1.95
+ $X2=1.89 $Y2=1.95
r216 21 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.95 $X2=1.71 $Y2=1.95
r217 21 22 22.9148 $w=3.05e-07 $l=1.45e-07 $layer=POLY_cond $X=1.71 $Y=1.95
+ $X2=1.855 $Y2=1.95
r218 17 27 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=8.115 $Y=3.235
+ $X2=8.115 $Y2=1.94
r219 13 26 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.045 $Y=0.85
+ $X2=8.045 $Y2=1.61
r220 9 19 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.925 $Y=0.85
+ $X2=1.925 $Y2=1.295
r221 3 22 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=2.115
+ $X2=1.855 $Y2=1.95
r222 3 5 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.855 $Y=2.115
+ $X2=1.855 $Y2=3.235
r223 2 23 10.4756 $w=2.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.785
+ $X2=1.89 $Y2=1.95
r224 1 19 38.6248 $w=2.2e-07 $l=1.1e-07 $layer=POLY_cond $X=1.89 $Y=1.405
+ $X2=1.89 $Y2=1.295
r225 1 2 110.842 $w=2.2e-07 $l=3.8e-07 $layer=POLY_cond $X=1.89 $Y=1.405
+ $X2=1.89 $Y2=1.785
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_432_424# 1 3 11 15 18 22 23 24 25 28
+ 29 30 32 35 41
c109 41 0 1.72079e-19 $X=3.795 $Y=0.755
c110 30 0 1.07085e-19 $X=2.855 $Y=2.705
c111 11 0 1.32807e-19 $X=2.285 $Y=0.85
r112 41 43 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=3.795 $Y=0.755
+ $X2=3.895 $Y2=0.755
r113 35 37 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=3.895 $Y=2.955
+ $X2=3.895 $Y2=3.635
r114 33 35 2.03372 $w=3.38e-07 $l=6e-08 $layer=LI1_cond $X=3.895 $Y=2.895
+ $X2=3.895 $Y2=2.955
r115 31 41 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.795 $Y=0.935
+ $X2=3.795 $Y2=0.755
r116 31 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.795 $Y=0.935
+ $X2=3.795 $Y2=1.2
r117 29 33 7.85115 $w=1.7e-07 $l=2.61534e-07 $layer=LI1_cond $X=3.725 $Y=2.705
+ $X2=3.895 $Y2=2.895
r118 29 30 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.725 $Y=2.705
+ $X2=2.855 $Y2=2.705
r119 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=2.62
+ $X2=2.855 $Y2=2.705
r120 27 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.77 $Y=2.37
+ $X2=2.77 $Y2=2.62
r121 26 40 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.38 $Y=2.285
+ $X2=2.295 $Y2=2.325
r122 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.685 $Y=2.285
+ $X2=2.77 $Y2=2.37
r123 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.685 $Y=2.285
+ $X2=2.38 $Y2=2.285
r124 23 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=1.285
+ $X2=3.795 $Y2=1.2
r125 23 24 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.71 $Y=1.285
+ $X2=2.38 $Y2=1.285
r126 22 40 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=2.2
+ $X2=2.295 $Y2=2.325
r127 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=1.37
+ $X2=2.38 $Y2=1.285
r128 21 22 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.295 $Y=1.37
+ $X2=2.295 $Y2=2.2
r129 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=2.285 $X2=2.295 $Y2=2.285
r130 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.285
+ $X2=2.295 $Y2=2.45
r131 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=2.285
+ $X2=2.295 $Y2=2.12
r132 15 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.285 $Y=3.235
+ $X2=2.285 $Y2=2.45
r133 11 19 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=2.285 $Y=0.85
+ $X2=2.285 $Y2=2.12
r134 3 37 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.605 $X2=3.895 $Y2=3.635
r135 3 35 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.605 $X2=3.895 $Y2=2.955
r136 1 43 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.575 $X2=3.895 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%D 3 7 10 14 19
c38 19 0 1.36979e-19 $X=3.295 $Y=1.74
c39 10 0 1.98306e-19 $X=3.295 $Y=1.74
c40 7 0 1.07085e-19 $X=3.235 $Y=3.235
r41 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.295 $Y=1.74
+ $X2=3.295 $Y2=1.74
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.74 $X2=3.295 $Y2=1.74
r43 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.74
+ $X2=3.295 $Y2=1.905
r44 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.74
+ $X2=3.295 $Y2=1.575
r45 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=3.235 $Y=3.235
+ $X2=3.235 $Y2=1.905
r46 3 11 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=3.235 $Y=0.85
+ $X2=3.235 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 67 70 71 72 73 80
c253 73 0 1.48522e-19 $X=6.03 $Y=2.11
c254 72 0 1.37846e-19 $X=6.735 $Y=2.11
c255 71 0 1.48522e-19 $X=3.8 $Y=2.11
c256 70 0 8.87231e-20 $X=5.74 $Y=2.11
c257 55 0 6.91727e-20 $X=5.49 $Y=2.11
c258 54 0 1.81195e-19 $X=5.77 $Y=2.11
c259 48 0 3.67809e-19 $X=4.135 $Y=1.4
c260 44 0 1.89329e-19 $X=4.05 $Y=2.11
c261 37 0 4.3775e-20 $X=5.855 $Y=2.285
c262 34 0 1.46493e-19 $X=5.405 $Y=1.235
c263 25 0 1.36979e-19 $X=3.685 $Y=2.285
r264 73 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.03 $Y=2.11
+ $X2=5.885 $Y2=2.11
r265 72 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.735 $Y=2.11
+ $X2=6.88 $Y2=2.11
r266 72 73 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.735 $Y=2.11
+ $X2=6.03 $Y2=2.11
r267 71 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.8 $Y=2.11
+ $X2=3.655 $Y2=2.11
r268 70 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.74 $Y=2.11
+ $X2=5.885 $Y2=2.11
r269 70 71 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.74 $Y=2.11
+ $X2=3.8 $Y2=2.11
r270 67 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=2.11
+ $X2=5.885 $Y2=2.11
r271 67 69 11.7308 $w=1.82e-07 $l=1.75e-07 $layer=LI1_cond $X=5.87 $Y=2.11
+ $X2=5.87 $Y2=2.285
r272 63 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.655 $Y=2.11
+ $X2=3.655 $Y2=2.11
r273 63 65 11.7308 $w=1.82e-07 $l=1.75e-07 $layer=LI1_cond $X=3.67 $Y=2.11
+ $X2=3.67 $Y2=2.285
r274 57 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.88 $Y=2.11
+ $X2=6.88 $Y2=2.11
r275 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.88 $Y=2.11
+ $X2=6.88 $Y2=2.285
r276 54 67 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.77 $Y=2.11 $X2=5.87
+ $Y2=2.11
r277 54 55 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.77 $Y=2.11
+ $X2=5.49 $Y2=2.11
r278 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.405 $Y=2.025
+ $X2=5.49 $Y2=2.11
r279 50 52 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.405 $Y=2.025
+ $X2=5.405 $Y2=1.4
r280 46 48 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.135 $Y=2.025
+ $X2=4.135 $Y2=1.4
r281 45 63 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.77 $Y=2.11 $X2=3.67
+ $Y2=2.11
r282 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.05 $Y=2.11
+ $X2=4.135 $Y2=2.025
r283 44 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.05 $Y=2.11
+ $X2=3.77 $Y2=2.11
r284 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=2.285 $X2=6.88 $Y2=2.285
r285 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.762 $Y=1.205
+ $X2=6.762 $Y2=1.355
r286 37 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.855
+ $Y=2.285 $X2=5.855 $Y2=2.285
r287 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.855 $Y=2.285
+ $X2=5.855 $Y2=2.45
r288 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.4 $X2=5.405 $Y2=1.4
r289 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.4
+ $X2=5.405 $Y2=1.235
r290 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.4 $X2=4.135 $Y2=1.4
r291 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.4
+ $X2=4.135 $Y2=1.235
r292 25 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.285 $X2=3.685 $Y2=2.285
r293 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.285
+ $X2=3.685 $Y2=2.45
r294 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.79 $Y=2.12
+ $X2=6.837 $Y2=2.285
r295 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.79 $Y=2.12
+ $X2=6.79 $Y2=1.355
r296 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.735 $Y=2.45
+ $X2=6.837 $Y2=2.285
r297 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.735 $Y=2.45
+ $X2=6.735 $Y2=3.235
r298 17 40 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.735 $Y=0.85
+ $X2=6.735 $Y2=1.205
r299 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.945 $Y=3.235
+ $X2=5.945 $Y2=2.45
r300 10 34 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.345 $Y=0.85
+ $X2=5.345 $Y2=1.235
r301 7 30 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.195 $Y=0.85
+ $X2=4.195 $Y2=1.235
r302 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.595 $Y=3.235
+ $X2=3.595 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_217_521# 1 3 11 15 17 18 21 22 27 31
+ 35 37 38 41 47 49 55 56 57 62
c164 62 0 7.97351e-20 $X=4.635 $Y=1.37
c165 57 0 1.32807e-19 $X=1.855 $Y=1.37
c166 56 0 2.71143e-19 $X=4.49 $Y=1.37
c167 49 0 1.63455e-19 $X=1.68 $Y=1.61
c168 47 0 1.5821e-19 $X=4.725 $Y=2.285
c169 41 0 1.63226e-19 $X=1.71 $Y=0.755
c170 37 0 1.95862e-19 $X=1.565 $Y=1.61
c171 31 0 6.36774e-20 $X=4.985 $Y=3.235
c172 22 0 1.89329e-19 $X=4.63 $Y=2.285
c173 21 0 6.91727e-20 $X=4.91 $Y=2.285
c174 15 0 6.36774e-20 $X=4.555 $Y=3.235
r175 57 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.37
+ $X2=1.71 $Y2=1.37
r176 56 62 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.49 $Y=1.37
+ $X2=4.635 $Y2=1.37
r177 56 57 2.53719 $w=1.7e-07 $l=2.635e-06 $layer=MET1_cond $X=4.49 $Y=1.37
+ $X2=1.855 $Y2=1.37
r178 53 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.37
+ $X2=4.635 $Y2=1.37
r179 53 55 5.43564 $w=2.02e-07 $l=9e-08 $layer=LI1_cond $X=4.635 $Y=1.345
+ $X2=4.725 $Y2=1.345
r180 49 50 8.57418 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.68 $Y=1.61
+ $X2=1.68 $Y2=1.455
r181 45 55 1.74864 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.725 $Y=1.455
+ $X2=4.725 $Y2=1.345
r182 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.725 $Y=1.455
+ $X2=4.725 $Y2=2.285
r183 44 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.37
+ $X2=1.71 $Y2=1.37
r184 44 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.37
+ $X2=1.71 $Y2=1.455
r185 41 44 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.71 $Y=0.755
+ $X2=1.71 $Y2=1.37
r186 37 49 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=1.61
+ $X2=1.68 $Y2=1.61
r187 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.565 $Y=1.61
+ $X2=1.295 $Y2=1.61
r188 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.695
+ $X2=1.295 $Y2=1.61
r189 33 35 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=1.21 $Y=1.695
+ $X2=1.21 $Y2=3.295
r190 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.985 $Y=2.42
+ $X2=4.985 $Y2=3.235
r191 25 27 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.985 $Y=1.265
+ $X2=4.985 $Y2=0.85
r192 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=2.285 $X2=4.725 $Y2=2.285
r193 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=2.285
+ $X2=4.725 $Y2=2.285
r194 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=2.285
+ $X2=4.985 $Y2=2.42
r195 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=2.285
+ $X2=4.725 $Y2=2.285
r196 20 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=1.4 $X2=4.725 $Y2=1.4
r197 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.63 $Y=1.4
+ $X2=4.725 $Y2=1.4
r198 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.91 $Y=1.4
+ $X2=4.985 $Y2=1.265
r199 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.91 $Y=1.4
+ $X2=4.725 $Y2=1.4
r200 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.63 $Y2=2.285
r201 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.555 $Y2=3.235
r202 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.265
+ $X2=4.63 $Y2=1.4
r203 9 11 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.555 $Y=1.265
+ $X2=4.555 $Y2=0.85
r204 3 35 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.605 $X2=1.21 $Y2=3.295
r205 1 41 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.575 $X2=1.71 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_704_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 50 54 59 63 67 69 70 75
c212 70 0 2.2497e-19 $X=6.05 $Y=1.725
c213 59 0 1.36413e-19 $X=7.22 $Y=2.62
c214 44 0 2.26569e-19 $X=5.885 $Y=1.725
c215 34 0 1.69503e-19 $X=3.715 $Y=1.28
c216 24 0 1.48522e-19 $X=5.345 $Y=3.235
c217 18 0 1.48522e-19 $X=4.195 $Y=3.235
r218 70 72 0.116207 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=6.05 $Y=1.725
+ $X2=5.885 $Y2=1.725
r219 69 75 0.0841272 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=6.835 $Y=1.725
+ $X2=6.95 $Y2=1.725
r220 69 70 0.755863 $w=1.7e-07 $l=7.85e-07 $layer=MET1_cond $X=6.835 $Y=1.725
+ $X2=6.05 $Y2=1.725
r221 65 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=2.705
+ $X2=7.22 $Y2=2.705
r222 62 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.95 $Y=1.725
+ $X2=6.95 $Y2=1.725
r223 62 63 16.1867 $w=1.83e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=1.717
+ $X2=7.22 $Y2=1.717
r224 59 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.62
+ $X2=7.22 $Y2=2.705
r225 58 63 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=7.22 $Y=1.81
+ $X2=7.22 $Y2=1.717
r226 58 59 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=7.22 $Y=1.81
+ $X2=7.22 $Y2=2.62
r227 54 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.95 $Y=2.955
+ $X2=6.95 $Y2=3.635
r228 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=2.79
+ $X2=6.95 $Y2=2.705
r229 52 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=2.79
+ $X2=6.95 $Y2=2.955
r230 48 62 1.22693 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=6.95 $Y=1.625
+ $X2=6.95 $Y2=1.717
r231 48 50 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.95 $Y=1.625
+ $X2=6.95 $Y2=0.755
r232 44 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.885 $Y=1.725
+ $X2=5.885 $Y2=1.725
r233 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=1.725 $X2=5.885 $Y2=1.725
r234 39 41 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=5.885 $Y=1.725
+ $X2=5.885 $Y2=1.85
r235 39 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.725
+ $X2=5.885 $Y2=1.56
r236 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.595 $Y=1.28
+ $X2=3.715 $Y2=1.28
r237 30 40 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.945 $Y=0.85
+ $X2=5.945 $Y2=1.56
r238 27 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=1.85
+ $X2=5.345 $Y2=1.85
r239 26 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.75 $Y=1.85
+ $X2=5.885 $Y2=1.85
r240 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.75 $Y=1.85
+ $X2=5.42 $Y2=1.85
r241 22 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.345 $Y=1.925
+ $X2=5.345 $Y2=1.85
r242 22 24 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=5.345 $Y=1.925
+ $X2=5.345 $Y2=3.235
r243 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=1.85
+ $X2=4.195 $Y2=1.85
r244 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=1.85
+ $X2=5.345 $Y2=1.85
r245 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.27 $Y=1.85 $X2=4.27
+ $Y2=1.85
r246 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=1.925
+ $X2=4.195 $Y2=1.85
r247 16 18 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=4.195 $Y=1.925
+ $X2=4.195 $Y2=3.235
r248 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=1.85
+ $X2=4.195 $Y2=1.85
r249 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.12 $Y=1.85
+ $X2=3.79 $Y2=1.85
r250 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=1.775
+ $X2=3.79 $Y2=1.85
r251 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.715 $Y=1.355
+ $X2=3.715 $Y2=1.28
r252 12 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.715 $Y=1.355
+ $X2=3.715 $Y2=1.775
r253 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.205
+ $X2=3.595 $Y2=1.28
r254 9 11 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=3.595 $Y=1.205
+ $X2=3.595 $Y2=0.85
r255 3 56 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=2.605 $X2=6.95 $Y2=3.635
r256 3 54 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=2.605 $X2=6.95 $Y2=2.955
r257 1 50 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.575 $X2=6.95 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1246_89# 1 3 11 15 23 26 28 32 33 35
+ 36 37 38 40 47 51 53 55 60 63 64 65 69 71
c211 47 0 1.63226e-19 $X=8.26 $Y=0.755
c212 40 0 1.6261e-19 $X=6.365 $Y=1.71
c213 37 0 8.77106e-20 $X=9.47 $Y=2.375
c214 33 0 3.77772e-20 $X=9.382 $Y=1.545
c215 32 0 2.20654e-19 $X=9.38 $Y=1.71
c216 11 0 1.35097e-19 $X=6.305 $Y=0.85
r217 67 69 0.105038 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=6.365 $Y=2.48
+ $X2=6.515 $Y2=2.48
r218 64 71 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.235 $Y=1.71
+ $X2=9.38 $Y2=1.71
r219 64 65 1.79096 $w=1.7e-07 $l=1.86e-06 $layer=MET1_cond $X=9.235 $Y=1.71
+ $X2=7.375 $Y2=1.71
r220 62 65 0.0706952 $w=1.7e-07 $l=1.14782e-07 $layer=MET1_cond $X=7.305
+ $Y=1.795 $X2=7.375 $Y2=1.71
r221 62 63 0.736385 $w=1.4e-07 $l=5.95e-07 $layer=MET1_cond $X=7.305 $Y=1.795
+ $X2=7.305 $Y2=2.39
r222 60 63 0.0709685 $w=1.75e-07 $l=1.80222e-07 $layer=MET1_cond $X=7.165
+ $Y=2.482 $X2=7.305 $Y2=2.39
r223 60 69 0.588306 $w=1.75e-07 $l=6.5e-07 $layer=MET1_cond $X=7.165 $Y=2.482
+ $X2=6.515 $Y2=2.482
r224 55 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.38 $Y=1.71
+ $X2=9.38 $Y2=1.71
r225 53 55 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.845 $Y=1.71
+ $X2=9.38 $Y2=1.71
r226 49 53 5.37722 $w=2.41e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=1.795
+ $X2=8.845 $Y2=1.71
r227 49 51 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=8.76 $Y=1.795
+ $X2=8.76 $Y2=3.295
r228 45 49 25.3112 $w=2.41e-07 $l=6.89202e-07 $layer=LI1_cond $X=8.26 $Y=1.345
+ $X2=8.76 $Y2=1.795
r229 45 47 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.26 $Y=1.345
+ $X2=8.26 $Y2=0.755
r230 43 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.365 $Y=2.48
+ $X2=6.365 $Y2=2.48
r231 40 43 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.365 $Y=1.71
+ $X2=6.365 $Y2=2.48
r232 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=2.375
+ $X2=9.47 $Y2=2.525
r233 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.47 $Y=1.23 $X2=9.47
+ $Y2=1.38
r234 34 37 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.445 $Y=1.875
+ $X2=9.445 $Y2=2.375
r235 33 36 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.445 $Y=1.545
+ $X2=9.445 $Y2=1.38
r236 32 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.38
+ $Y=1.71 $X2=9.38 $Y2=1.71
r237 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=1.71
+ $X2=9.382 $Y2=1.875
r238 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.382 $Y=1.71
+ $X2=9.382 $Y2=1.545
r239 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=1.71 $X2=6.365 $Y2=1.71
r240 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.71
+ $X2=6.365 $Y2=1.875
r241 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.71
+ $X2=6.365 $Y2=1.545
r242 26 38 228.147 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=9.495 $Y=3.235
+ $X2=9.495 $Y2=2.525
r243 23 35 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.495 $Y=0.85
+ $X2=9.495 $Y2=1.23
r244 15 30 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=6.305 $Y=3.235
+ $X2=6.305 $Y2=1.875
r245 11 29 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.305 $Y=0.85
+ $X2=6.305 $Y2=1.545
r246 3 51 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=8.62
+ $Y=2.605 $X2=8.76 $Y2=3.295
r247 1 47 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=8.12
+ $Y=0.575 $X2=8.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1084_115# 1 3 10 11 13 16 20 26 30 32
+ 33 36 40 43 49 52 53 54 55 62
c177 55 0 2.81591e-19 $X=5.89 $Y=1.37
c178 53 0 1.5821e-19 $X=5.21 $Y=1.37
c179 49 0 1.71621e-19 $X=5.645 $Y=0.755
c180 30 0 1.57671e-19 $X=5.065 $Y=1.37
c181 16 0 6.36774e-20 $X=7.685 $Y=3.235
r182 55 60 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=5.89 $Y=1.37
+ $X2=5.745 $Y2=1.34
r183 54 62 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=1.37
+ $X2=7.595 $Y2=1.37
r184 54 55 1.5021 $w=1.7e-07 $l=1.56e-06 $layer=MET1_cond $X=7.45 $Y=1.37
+ $X2=5.89 $Y2=1.37
r185 53 57 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.21 $Y=1.37
+ $X2=5.065 $Y2=1.37
r186 52 60 0.0886454 $w=2.23e-07 $l=1.59295e-07 $layer=MET1_cond $X=5.6 $Y=1.37
+ $X2=5.745 $Y2=1.34
r187 52 53 0.375524 $w=1.7e-07 $l=3.9e-07 $layer=MET1_cond $X=5.6 $Y=1.37
+ $X2=5.21 $Y2=1.37
r188 49 51 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=5.652 $Y=0.755
+ $X2=5.652 $Y2=1.035
r189 43 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=1.37
+ $X2=7.595 $Y2=1.37
r190 43 46 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.595 $Y=1.37
+ $X2=7.595 $Y2=2.285
r191 40 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=1.34
r192 40 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=1.035
r193 34 36 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=5.645 $Y=2.79
+ $X2=5.645 $Y2=3.295
r194 32 34 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.475 $Y=2.705
+ $X2=5.645 $Y2=2.79
r195 32 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.475 $Y=2.705
+ $X2=5.15 $Y2=2.705
r196 30 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.065 $Y=1.37
+ $X2=5.065 $Y2=1.37
r197 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=2.62
+ $X2=5.15 $Y2=2.705
r198 28 30 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.065 $Y=2.62
+ $X2=5.065 $Y2=1.37
r199 25 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=2.285 $X2=7.595 $Y2=2.285
r200 25 26 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=2.285
+ $X2=7.685 $Y2=2.285
r201 22 25 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=2.285
+ $X2=7.595 $Y2=2.285
r202 18 20 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=7.505 $Y=1.29
+ $X2=7.685 $Y2=1.29
r203 14 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.685 $Y=2.42
+ $X2=7.685 $Y2=2.285
r204 14 16 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=7.685 $Y=2.42
+ $X2=7.685 $Y2=3.235
r205 11 20 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.685 $Y=1.21
+ $X2=7.685 $Y2=1.29
r206 11 13 115.68 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.685 $Y=1.21
+ $X2=7.685 $Y2=0.85
r207 10 22 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.505 $Y=2.15
+ $X2=7.505 $Y2=2.285
r208 9 18 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.505 $Y=1.37
+ $X2=7.505 $Y2=1.29
r209 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.505 $Y=1.37
+ $X2=7.505 $Y2=2.15
r210 3 36 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=5.42
+ $Y=2.605 $X2=5.645 $Y2=3.295
r211 1 49 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=5.42
+ $Y=0.575 $X2=5.645 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c83 44 0 8.77106e-20 $X=9.285 $Y=2.48
c84 35 0 9.99996e-20 $X=9.78 $Y=2.285
c85 34 0 8.31638e-20 $X=9.365 $Y=1.37
c86 33 0 1.20654e-19 $X=9.78 $Y=1.37
c87 27 0 1.09867e-19 $X=9.28 $Y=2.48
c88 18 0 1.98165e-19 $X=9.865 $Y=1.915
r89 42 44 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=9.28 $Y=2.48
+ $X2=9.285 $Y2=2.48
r90 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.865 $Y=2.2
+ $X2=9.865 $Y2=1.915
r91 37 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.865 $Y=1.455
+ $X2=9.865 $Y2=1.915
r92 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=2.285
+ $X2=9.865 $Y2=2.2
r93 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=2.285
+ $X2=9.365 $Y2=2.285
r94 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.37
+ $X2=9.865 $Y2=1.455
r95 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.78 $Y=1.37
+ $X2=9.365 $Y2=1.37
r96 29 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.28 $Y=2.955
+ $X2=9.28 $Y2=3.635
r97 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=2.48
+ $X2=9.28 $Y2=2.48
r98 27 29 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=9.28 $Y=2.48
+ $X2=9.28 $Y2=2.955
r99 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=2.37
+ $X2=9.365 $Y2=2.285
r100 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.28 $Y=2.37
+ $X2=9.28 $Y2=2.48
r101 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=1.285
+ $X2=9.365 $Y2=1.37
r102 21 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.28 $Y=1.285
+ $X2=9.28 $Y2=0.755
r103 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.865
+ $Y=1.915 $X2=9.865 $Y2=1.915
r104 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=1.915
+ $X2=9.865 $Y2=2.08
r105 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=1.915
+ $X2=9.865 $Y2=1.75
r106 15 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.925 $Y=3.235
+ $X2=9.925 $Y2=2.08
r107 11 19 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=9.925 $Y=0.85
+ $X2=9.925 $Y2=1.75
r108 3 31 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=2.605 $X2=9.28 $Y2=3.635
r109 3 29 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=2.605 $X2=9.28 $Y2=2.955
r110 1 23 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.575 $X2=9.28 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_300_521# 1 2 11 13 14 17
c20 1 0 1.5152e-19 $X=1.5 $Y=2.605
r21 15 17 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.5 $Y=3.275 $X2=2.5
+ $Y2=3.295
r22 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=3.19
+ $X2=2.5 $Y2=3.275
r23 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.415 $Y=3.19
+ $X2=1.725 $Y2=3.19
r24 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.275
+ $X2=1.725 $Y2=3.19
r25 9 11 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.64 $Y=3.275 $X2=1.64
+ $Y2=3.295
r26 2 17 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=2.605 $X2=2.5 $Y2=3.295
r27 1 11 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.605 $X2=1.64 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%A_1469_521# 1 2 11 13 14 17
r20 15 17 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.33 $Y=3.27
+ $X2=8.33 $Y2=3.295
r21 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.245 $Y=3.185
+ $X2=8.33 $Y2=3.27
r22 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.245 $Y=3.185
+ $X2=7.555 $Y2=3.185
r23 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=3.27
+ $X2=7.555 $Y2=3.185
r24 9 11 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.47 $Y=3.27 $X2=7.47
+ $Y2=3.295
r25 2 17 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=2.605 $X2=8.33 $Y2=3.295
r26 1 11 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=2.605 $X2=7.47 $Y2=3.295
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFSR_1%Q 1 3 11 15 22 25 29 32
r19 27 29 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=2.61
+ $X2=10.255 $Y2=2.61
r20 23 25 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.14 $Y=1.035
+ $X2=10.255 $Y2=1.035
r21 22 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=2.525
+ $X2=10.255 $Y2=2.61
r22 21 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.255 $Y=1.12
+ $X2=10.255 $Y2=1.035
r23 21 22 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=10.255 $Y=1.12
+ $X2=10.255 $Y2=2.525
r24 17 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=10.14 $Y=2.955
+ $X2=10.14 $Y2=3.635
r25 15 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.14 $Y=2.85
+ $X2=10.14 $Y2=2.85
r26 15 17 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=10.14 $Y=2.85
+ $X2=10.14 $Y2=2.955
r27 13 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=2.695
+ $X2=10.14 $Y2=2.61
r28 13 15 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.14 $Y=2.695
+ $X2=10.14 $Y2=2.85
r29 9 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.14 $Y=0.95
+ $X2=10.14 $Y2=1.035
r30 9 11 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.14 $Y=0.95
+ $X2=10.14 $Y2=0.755
r31 3 19 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=10
+ $Y=2.605 $X2=10.14 $Y2=3.635
r32 3 17 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=10
+ $Y=2.605 $X2=10.14 $Y2=2.955
r33 1 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=10 $Y=0.575
+ $X2=10.14 $Y2=0.755
.ends

