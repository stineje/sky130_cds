* File: sky130_osu_sc_18T_hs__nor2_1.pex.spice
* Created: Fri Nov 12 13:51:48 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__NOR2_1%GND 1 2 21 25 27 35 41 44
r27 41 44 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r28 33 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r29 27 33 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.305
r30 23 25 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r31 21 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r32 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r33 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r34 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r35 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r36 2 35 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r37 1 25 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NOR2_1%VDD 1 13 15 21 29 32
r18 29 32 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r19 26 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r20 21 24 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.05 $Y=4.135
+ $X2=1.05 $Y2=5.835
r21 19 26 4.25596 $w=1.7e-07 $l=2.13185e-07 $layer=LI1_cond $X=1.05 $Y=6.355
+ $X2=1.197 $Y2=6.507
r22 19 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=6.355
+ $X2=1.05 $Y2=5.835
r23 15 26 3.30228 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=0.965 $Y=6.507
+ $X2=1.197 $Y2=6.507
r24 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=6.507
+ $X2=0.34 $Y2=6.507
r25 13 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r26 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r27 1 24 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.91
+ $Y=3.085 $X2=1.05 $Y2=5.835
r28 1 21 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.91
+ $Y=3.085 $X2=1.05 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NOR2_1%B 3 7 10 13 19 22
r49 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.65 $Y=2.96
+ $X2=0.65 $Y2=2.96
r50 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.65 $Y=2.175
+ $X2=0.65 $Y2=2.96
r51 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=2.09
+ $X2=0.65 $Y2=2.175
r52 13 15 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.565 $Y=2.09
+ $X2=0.415 $Y2=2.09
r53 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=2.09 $X2=0.415 $Y2=2.09
r54 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.09
+ $X2=0.415 $Y2=2.255
r55 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.09
+ $X2=0.415 $Y2=1.925
r56 7 12 1194.74 $w=1.5e-07 $l=2.33e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.255
r57 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=1.925
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NOR2_1%A 3 7 10 14 20
r36 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=3.33
+ $X2=0.99 $Y2=3.33
r37 14 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.99 $Y=2.755
+ $X2=0.99 $Y2=3.33
r38 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.755 $X2=0.99 $Y2=2.755
r39 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.755
+ $X2=0.942 $Y2=2.92
r40 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.755
+ $X2=0.942 $Y2=2.59
r41 7 11 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.59
r42 3 12 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=0.835 $Y=4.585
+ $X2=0.835 $Y2=2.92
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NOR2_1%Y 1 3 10 18 23 24 28 34
r41 26 28 0.519956 $w=1.7e-07 $l=5.4e-07 $layer=MET1_cond $X=0.69 $Y=2.505
+ $X2=0.69 $Y2=1.965
r42 25 34 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.48
r43 25 28 0.356266 $w=1.7e-07 $l=3.7e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.965
r44 24 31 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=2.59
+ $X2=0.26 $Y2=2.59
r45 23 26 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=0.605 $Y=2.59
+ $X2=0.69 $Y2=2.505
r46 23 24 0.192576 $w=1.7e-07 $l=2e-07 $layer=MET1_cond $X=0.605 $Y=2.59
+ $X2=0.405 $Y2=2.59
r47 21 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.48
r48 18 21 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.69 $Y=0.825
+ $X2=0.69 $Y2=1.48
r49 13 15 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r50 10 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.59
+ $X2=0.26 $Y2=2.59
r51 10 13 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=0.26 $Y=2.59
+ $X2=0.26 $Y2=3.455
r52 3 15 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r53 3 13 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r54 1 18 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

