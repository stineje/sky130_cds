* File: sky130_osu_sc_15T_ms__buf_1.pex.spice
* Created: Fri Nov 12 14:41:22 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__BUF_1%GND 1 17 19 26 36 39
r27 36 39 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r28 28 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r29 24 34 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r30 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.74
r31 19 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r32 17 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r33 17 28 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r34 17 19 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r35 1 26 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__BUF_1%VDD 1 13 15 21 27 32 35
r21 32 35 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r22 27 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r23 25 30 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=0.69 $Y2=5.397
r24 25 27 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=5.397
+ $X2=1.02 $Y2=5.397
r25 21 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=3.895
+ $X2=0.69 $Y2=4.575
r26 19 30 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=5.397
r27 19 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.69 $Y=5.245
+ $X2=0.69 $Y2=4.575
r28 15 30 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.69 $Y2=5.397
r29 15 17 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=5.397
+ $X2=0.34 $Y2=5.397
r30 13 27 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r31 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r32 1 24 400 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.575
r33 1 21 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__BUF_1%A 3 7 10 14 20
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.07
+ $X2=0.635 $Y2=3.07
r41 14 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=2.22
+ $X2=0.635 $Y2=3.07
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.22 $X2=0.635 $Y2=2.22
r43 10 12 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.22
+ $X2=0.585 $Y2=2.385
r44 10 11 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.22
+ $X2=0.585 $Y2=2.055
r45 7 12 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=0.475 $Y=3.825
+ $X2=0.475 $Y2=2.385
r46 3 11 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__BUF_1%A_27_115# 1 3 11 13 15 17 22 26 30 34 38
+ 40 43
r55 39 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.675
+ $X2=0.26 $Y2=1.675
r56 38 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.675
+ $X2=0.965 $Y2=1.675
r57 38 39 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.675
+ $X2=0.345 $Y2=1.675
r58 34 36 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=4.575
r59 32 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.76 $X2=0.26
+ $Y2=1.675
r60 32 34 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=0.26 $Y=1.76
+ $X2=0.26 $Y2=3.215
r61 28 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.59 $X2=0.26
+ $Y2=1.675
r62 28 30 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.74
r63 24 26 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.675
+ $X2=1.18 $Y2=2.675
r64 21 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.675 $X2=0.965 $Y2=1.675
r65 21 22 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=1.18 $Y2=1.675
r66 18 21 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.965 $Y2=1.675
r67 17 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.6 $X2=1.18
+ $Y2=2.675
r68 16 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.84
+ $X2=1.18 $Y2=1.675
r69 16 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=1.84
+ $X2=1.18 $Y2=2.6
r70 13 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=2.675
r71 13 15 345.433 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.905 $Y=2.75
+ $X2=0.905 $Y2=3.825
r72 9 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.905 $Y2=1.675
r73 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.905 $Y2=0.945
r74 3 36 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r75 3 34 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.215
r76 1 30 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__BUF_1%Y 1 3 10 16 26 29 32
r33 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.585
+ $X2=1.12 $Y2=2.7
r34 24 26 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.12 $Y=2.585
+ $X2=1.12 $Y2=2.015
r35 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=1.22
r36 23 26 0.65476 $w=1.7e-07 $l=6.8e-07 $layer=MET1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=2.015
r37 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.12 $Y=3.215
+ $X2=1.12 $Y2=4.575
r38 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.7 $X2=1.12
+ $Y2=2.7
r39 16 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.12 $Y=2.7
+ $X2=1.12 $Y2=3.215
r40 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.22
+ $X2=1.12 $Y2=1.22
r41 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.12 $Y=0.74
+ $X2=1.12 $Y2=1.22
r42 3 21 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r43 3 19 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.215
r44 1 10 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.74
.ends

