* File: sky130_osu_sc_18T_ms__dffs_1.pxi.spice
* Created: Fri Nov 12 14:02:58 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%GND N_GND_M1000_d N_GND_M1001_s N_GND_M1022_d
+ N_GND_M1008_d N_GND_M1027_d N_GND_M1010_d N_GND_M1014_b N_GND_c_2_p
+ N_GND_c_20_p N_GND_c_21_p N_GND_c_42_p N_GND_c_22_p N_GND_c_61_p N_GND_c_23_p
+ N_GND_c_6_p N_GND_c_7_p N_GND_c_142_p N_GND_c_143_p GND N_GND_c_3_p
+ PM_SKY130_OSU_SC_18T_MS__DFFS_1%GND
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%VDD N_VDD_M1026_s N_VDD_M1017_d N_VDD_M1002_s
+ N_VDD_M1023_d N_VDD_M1009_d N_VDD_M1020_s N_VDD_M1021_d N_VDD_M1011_d
+ N_VDD_M1026_b N_VDD_c_194_p N_VDD_c_195_p N_VDD_c_203_p N_VDD_c_204_p
+ N_VDD_c_212_p N_VDD_c_238_p N_VDD_c_222_p N_VDD_c_226_p N_VDD_c_227_p
+ N_VDD_c_228_p N_VDD_c_198_p N_VDD_c_199_p N_VDD_c_268_p N_VDD_c_269_p
+ N_VDD_c_284_p VDD N_VDD_c_196_p PM_SKY130_OSU_SC_18T_MS__DFFS_1%VDD
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%SN N_SN_M1014_g N_SN_M1026_g N_SN_c_301_n
+ N_SN_M1027_g N_SN_M1021_g N_SN_c_306_n N_SN_c_307_n N_SN_c_309_n N_SN_c_310_n
+ N_SN_c_312_n N_SN_c_320_n SN N_SN_c_321_n PM_SKY130_OSU_SC_18T_MS__DFFS_1%SN
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_152_89# N_A_152_89#_M1024_d
+ N_A_152_89#_M1025_d N_A_152_89#_M1000_g N_A_152_89#_M1017_g
+ N_A_152_89#_c_433_n N_A_152_89#_c_434_n N_A_152_89#_c_435_n
+ N_A_152_89#_c_438_n N_A_152_89#_c_450_n N_A_152_89#_c_453_n
+ N_A_152_89#_c_440_n N_A_152_89#_c_441_n N_A_152_89#_c_454_n
+ N_A_152_89#_c_466_n PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_152_89#
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%D N_D_M1001_g N_D_M1002_g N_D_c_518_n
+ N_D_c_519_n D PM_SKY130_OSU_SC_18T_MS__DFFS_1%D
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%CK N_CK_M1025_g N_CK_M1018_g N_CK_M1012_g
+ N_CK_M1005_g N_CK_M1004_g N_CK_c_554_n N_CK_M1006_g N_CK_c_555_n N_CK_c_556_n
+ N_CK_c_557_n N_CK_c_558_n N_CK_c_561_n N_CK_c_562_n N_CK_c_565_n N_CK_c_566_n
+ N_CK_c_570_n N_CK_c_571_n N_CK_c_572_n N_CK_c_573_n N_CK_c_574_n N_CK_c_575_n
+ N_CK_c_576_n N_CK_c_577_n N_CK_c_578_n N_CK_c_579_n N_CK_c_580_n N_CK_c_581_n
+ N_CK_c_582_n CK PM_SKY130_OSU_SC_18T_MS__DFFS_1%CK
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_27_115# N_A_27_115#_M1014_s
+ N_A_27_115#_M1026_d N_A_27_115#_M1022_g N_A_27_115#_M1023_g
+ N_A_27_115#_c_776_n N_A_27_115#_c_778_n N_A_27_115#_c_779_n
+ N_A_27_115#_c_780_n N_A_27_115#_M1015_g N_A_27_115#_M1016_g
+ N_A_27_115#_c_785_n N_A_27_115#_c_811_n N_A_27_115#_c_815_n
+ N_A_27_115#_c_788_n N_A_27_115#_c_789_n N_A_27_115#_c_790_n
+ N_A_27_115#_c_792_n N_A_27_115#_c_793_n N_A_27_115#_c_827_n
+ PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_27_115#
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_428_89# N_A_428_89#_M1004_d
+ N_A_428_89#_M1006_d N_A_428_89#_c_899_n N_A_428_89#_M1024_g
+ N_A_428_89#_c_902_n N_A_428_89#_c_903_n N_A_428_89#_c_904_n
+ N_A_428_89#_M1019_g N_A_428_89#_c_906_n N_A_428_89#_M1013_g
+ N_A_428_89#_c_908_n N_A_428_89#_c_909_n N_A_428_89#_M1003_g
+ N_A_428_89#_c_910_n N_A_428_89#_c_911_n N_A_428_89#_c_912_n
+ N_A_428_89#_c_913_n N_A_428_89#_c_914_n N_A_428_89#_c_917_n
+ N_A_428_89#_c_919_n N_A_428_89#_c_923_n N_A_428_89#_c_933_n
+ N_A_428_89#_c_924_n N_A_428_89#_c_925_n N_A_428_89#_c_926_n
+ N_A_428_89#_c_938_n PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_428_89#
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_970_89# N_A_970_89#_M1007_s
+ N_A_970_89#_M1020_d N_A_970_89#_M1008_g N_A_970_89#_M1009_g
+ N_A_970_89#_M1010_g N_A_970_89#_M1011_g N_A_970_89#_c_1092_n
+ N_A_970_89#_c_1093_n N_A_970_89#_c_1094_n N_A_970_89#_c_1095_n
+ N_A_970_89#_c_1100_n N_A_970_89#_c_1101_n N_A_970_89#_c_1102_n
+ N_A_970_89#_c_1103_n N_A_970_89#_c_1104_n N_A_970_89#_c_1130_n
+ N_A_970_89#_c_1132_n N_A_970_89#_c_1107_n N_A_970_89#_c_1108_n
+ N_A_970_89#_c_1109_n N_A_970_89#_c_1110_n N_A_970_89#_c_1111_n
+ N_A_970_89#_c_1112_n N_A_970_89#_c_1113_n
+ PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_970_89#
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_808_115# N_A_808_115#_M1012_d
+ N_A_808_115#_M1013_d N_A_808_115#_M1007_g N_A_808_115#_M1020_g
+ N_A_808_115#_c_1255_n N_A_808_115#_c_1256_n N_A_808_115#_c_1280_n
+ N_A_808_115#_c_1281_n N_A_808_115#_c_1297_n N_A_808_115#_c_1325_n
+ N_A_808_115#_c_1257_n N_A_808_115#_c_1270_n N_A_808_115#_c_1260_n
+ N_A_808_115#_c_1261_n N_A_808_115#_c_1263_n N_A_808_115#_c_1264_n
+ PM_SKY130_OSU_SC_18T_MS__DFFS_1%A_808_115#
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%QN N_QN_M1010_s N_QN_M1011_s N_QN_M1028_g
+ N_QN_M1029_g N_QN_c_1383_n N_QN_c_1384_n N_QN_c_1388_n N_QN_c_1389_n
+ N_QN_c_1390_n N_QN_c_1391_n N_QN_c_1392_n N_QN_c_1393_n QN
+ PM_SKY130_OSU_SC_18T_MS__DFFS_1%QN
x_PM_SKY130_OSU_SC_18T_MS__DFFS_1%Q N_Q_M1028_d N_Q_M1029_d N_Q_c_1464_n
+ N_Q_c_1468_n N_Q_c_1466_n N_Q_c_1467_n N_Q_c_1472_n Q
+ PM_SKY130_OSU_SC_18T_MS__DFFS_1%Q
cc_1 N_GND_M1014_b N_SN_M1014_g 0.0366893f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_SN_M1014_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_SN_M1014_g 0.00468827f $X=7.815 $Y=0.19 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1014_b N_SN_M1026_g 0.0715368f $X=-0.05 $Y=0 $X2=0.475 $Y2=5.085
cc_5 N_GND_M1014_b N_SN_c_301_n 0.0172063f $X=-0.05 $Y=0 $X2=6.665 $Y2=1.425
cc_6 N_GND_c_6_p N_SN_c_301_n 0.00606474f $X=6.795 $Y=0.152 $X2=6.665 $Y2=1.425
cc_7 N_GND_c_7_p N_SN_c_301_n 0.00713292f $X=6.88 $Y=0.825 $X2=6.665 $Y2=1.425
cc_8 N_GND_c_3_p N_SN_c_301_n 0.00468827f $X=7.815 $Y=0.19 $X2=6.665 $Y2=1.425
cc_9 N_GND_M1014_b N_SN_M1021_g 0.0790728f $X=-0.05 $Y=0 $X2=6.735 $Y2=5.085
cc_10 N_GND_M1014_b N_SN_c_306_n 0.047507f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.85
cc_11 N_GND_M1014_b N_SN_c_307_n 0.0414397f $X=-0.05 $Y=0 $X2=6.735 $Y2=1.59
cc_12 N_GND_c_7_p N_SN_c_307_n 0.0016316f $X=6.88 $Y=0.825 $X2=6.735 $Y2=1.59
cc_13 N_GND_M1014_b N_SN_c_309_n 0.0129875f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.48
cc_14 N_GND_M1014_b N_SN_c_310_n 0.0028593f $X=-0.05 $Y=0 $X2=6.86 $Y2=1.48
cc_15 N_GND_c_7_p N_SN_c_310_n 0.00557352f $X=6.88 $Y=0.825 $X2=6.86 $Y2=1.48
cc_16 N_GND_M1001_s N_SN_c_312_n 0.00506021f $X=1.515 $Y=0.575 $X2=6.715
+ $Y2=1.48
cc_17 N_GND_M1022_d N_SN_c_312_n 0.0109039f $X=3.25 $Y=0.575 $X2=6.715 $Y2=1.48
cc_18 N_GND_M1008_d N_SN_c_312_n 0.00557645f $X=5 $Y=0.575 $X2=6.715 $Y2=1.48
cc_19 N_GND_M1014_b N_SN_c_312_n 0.0397781f $X=-0.05 $Y=0 $X2=6.715 $Y2=1.48
cc_20 N_GND_c_20_p N_SN_c_312_n 0.00484697f $X=1.05 $Y=0.825 $X2=6.715 $Y2=1.48
cc_21 N_GND_c_21_p N_SN_c_312_n 0.0120854f $X=1.64 $Y=0.825 $X2=6.715 $Y2=1.48
cc_22 N_GND_c_22_p N_SN_c_312_n 0.00558854f $X=3.39 $Y=0.825 $X2=6.715 $Y2=1.48
cc_23 N_GND_c_23_p N_SN_c_312_n 0.0119903f $X=5.14 $Y=0.825 $X2=6.715 $Y2=1.48
cc_24 N_GND_M1014_b N_SN_c_320_n 0.0119644f $X=-0.05 $Y=0 $X2=0.465 $Y2=1.48
cc_25 N_GND_M1014_b N_SN_c_321_n 0.00737611f $X=-0.05 $Y=0 $X2=6.86 $Y2=1.48
cc_26 N_GND_c_7_p N_SN_c_321_n 0.00500768f $X=6.88 $Y=0.825 $X2=6.86 $Y2=1.48
cc_27 N_GND_M1014_b N_A_152_89#_M1000_g 0.0578472f $X=-0.05 $Y=0 $X2=0.835
+ $Y2=0.945
cc_28 N_GND_c_2_p N_A_152_89#_M1000_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835
+ $Y2=0.945
cc_29 N_GND_c_20_p N_A_152_89#_M1000_g 0.00713292f $X=1.05 $Y=0.825 $X2=0.835
+ $Y2=0.945
cc_30 N_GND_c_21_p N_A_152_89#_M1000_g 0.00829768f $X=1.64 $Y=0.825 $X2=0.835
+ $Y2=0.945
cc_31 N_GND_c_3_p N_A_152_89#_M1000_g 0.00468827f $X=7.815 $Y=0.19 $X2=0.835
+ $Y2=0.945
cc_32 N_GND_M1014_b N_A_152_89#_M1017_g 0.0275072f $X=-0.05 $Y=0 $X2=0.905
+ $Y2=5.085
cc_33 N_GND_M1014_b N_A_152_89#_c_433_n 0.0440769f $X=-0.05 $Y=0 $X2=1.03
+ $Y2=2.305
cc_34 N_GND_M1014_b N_A_152_89#_c_434_n 0.0125993f $X=-0.05 $Y=0 $X2=1.03
+ $Y2=2.305
cc_35 N_GND_M1014_b N_A_152_89#_c_435_n 0.0257852f $X=-0.05 $Y=0 $X2=2.33
+ $Y2=1.765
cc_36 N_GND_c_20_p N_A_152_89#_c_435_n 2.45692e-19 $X=1.05 $Y=0.825 $X2=2.33
+ $Y2=1.765
cc_37 N_GND_c_21_p N_A_152_89#_c_435_n 0.00673409f $X=1.64 $Y=0.825 $X2=2.33
+ $Y2=1.765
cc_38 N_GND_M1014_b N_A_152_89#_c_438_n 0.00378473f $X=-0.05 $Y=0 $X2=1.115
+ $Y2=1.765
cc_39 N_GND_c_20_p N_A_152_89#_c_438_n 0.00216341f $X=1.05 $Y=0.825 $X2=1.115
+ $Y2=1.765
cc_40 N_GND_M1014_b N_A_152_89#_c_440_n 0.00198494f $X=-0.05 $Y=0 $X2=2.415
+ $Y2=1.68
cc_41 N_GND_M1014_b N_A_152_89#_c_441_n 0.00313975f $X=-0.05 $Y=0 $X2=2.515
+ $Y2=0.825
cc_42 N_GND_c_42_p N_A_152_89#_c_441_n 0.0149461f $X=3.305 $Y=0.152 $X2=2.515
+ $Y2=0.825
cc_43 N_GND_c_3_p N_A_152_89#_c_441_n 0.00958198f $X=7.815 $Y=0.19 $X2=2.515
+ $Y2=0.825
cc_44 N_GND_M1014_b N_D_M1001_g 0.0421748f $X=-0.05 $Y=0 $X2=1.855 $Y2=1.075
cc_45 N_GND_c_21_p N_D_M1001_g 0.0071489f $X=1.64 $Y=0.825 $X2=1.855 $Y2=1.075
cc_46 N_GND_c_42_p N_D_M1001_g 0.00606474f $X=3.305 $Y=0.152 $X2=1.855 $Y2=1.075
cc_47 N_GND_c_3_p N_D_M1001_g 0.00468827f $X=7.815 $Y=0.19 $X2=1.855 $Y2=1.075
cc_48 N_GND_M1014_b N_D_M1002_g 0.0367665f $X=-0.05 $Y=0 $X2=1.855 $Y2=4.585
cc_49 N_GND_M1014_b N_D_c_518_n 0.0305253f $X=-0.05 $Y=0 $X2=1.915 $Y2=2.22
cc_50 N_GND_M1014_b N_D_c_519_n 0.00311208f $X=-0.05 $Y=0 $X2=1.915 $Y2=2.22
cc_51 N_GND_M1014_b D 0.01184f $X=-0.05 $Y=0 $X2=1.915 $Y2=2.22
cc_52 N_GND_M1014_b N_CK_c_554_n 0.0311248f $X=-0.05 $Y=0 $X2=5.355 $Y2=2.93
cc_53 N_GND_M1014_b N_CK_c_555_n 0.0444827f $X=-0.05 $Y=0 $X2=5.41 $Y2=2.6
cc_54 N_GND_M1014_b N_CK_c_556_n 0.0244095f $X=-0.05 $Y=0 $X2=2.275 $Y2=2.765
cc_55 N_GND_M1014_b N_CK_c_557_n 0.0254608f $X=-0.05 $Y=0 $X2=2.755 $Y2=1.85
cc_56 N_GND_M1014_b N_CK_c_558_n 0.0173906f $X=-0.05 $Y=0 $X2=2.755 $Y2=1.685
cc_57 N_GND_c_42_p N_CK_c_558_n 0.00606474f $X=3.305 $Y=0.152 $X2=2.755
+ $Y2=1.685
cc_58 N_GND_c_3_p N_CK_c_558_n 0.00468827f $X=7.815 $Y=0.19 $X2=2.755 $Y2=1.685
cc_59 N_GND_M1014_b N_CK_c_561_n 0.0252285f $X=-0.05 $Y=0 $X2=4.025 $Y2=1.85
cc_60 N_GND_M1014_b N_CK_c_562_n 0.0175305f $X=-0.05 $Y=0 $X2=4.025 $Y2=1.685
cc_61 N_GND_c_61_p N_CK_c_562_n 0.00606474f $X=5.055 $Y=0.152 $X2=4.025
+ $Y2=1.685
cc_62 N_GND_c_3_p N_CK_c_562_n 0.00468827f $X=7.815 $Y=0.19 $X2=4.025 $Y2=1.685
cc_63 N_GND_M1014_b N_CK_c_565_n 0.0233827f $X=-0.05 $Y=0 $X2=4.505 $Y2=2.765
cc_64 N_GND_M1014_b N_CK_c_566_n 0.0206446f $X=-0.05 $Y=0 $X2=5.382 $Y2=1.685
cc_65 N_GND_c_23_p N_CK_c_566_n 0.00356864f $X=5.14 $Y=0.825 $X2=5.382 $Y2=1.685
cc_66 N_GND_c_6_p N_CK_c_566_n 0.00606474f $X=6.795 $Y=0.152 $X2=5.382 $Y2=1.685
cc_67 N_GND_c_3_p N_CK_c_566_n 0.00468827f $X=7.815 $Y=0.19 $X2=5.382 $Y2=1.685
cc_68 N_GND_M1014_b N_CK_c_570_n 0.0128304f $X=-0.05 $Y=0 $X2=5.382 $Y2=1.835
cc_69 N_GND_M1014_b N_CK_c_571_n 0.00609317f $X=-0.05 $Y=0 $X2=2.67 $Y2=2.59
cc_70 N_GND_M1014_b N_CK_c_572_n 0.00921066f $X=-0.05 $Y=0 $X2=2.755 $Y2=1.85
cc_71 N_GND_M1014_b N_CK_c_573_n 0.00838835f $X=-0.05 $Y=0 $X2=4.025 $Y2=1.85
cc_72 N_GND_M1014_b N_CK_c_574_n 0.00543853f $X=-0.05 $Y=0 $X2=4.42 $Y2=2.59
cc_73 N_GND_M1014_b N_CK_c_575_n 5.00459e-19 $X=-0.05 $Y=0 $X2=4.11 $Y2=2.59
cc_74 N_GND_M1014_b N_CK_c_576_n 6.58573e-19 $X=-0.05 $Y=0 $X2=5.5 $Y2=2.59
cc_75 N_GND_M1014_b N_CK_c_577_n 0.00276905f $X=-0.05 $Y=0 $X2=2.275 $Y2=2.59
cc_76 N_GND_M1014_b N_CK_c_578_n 0.00265612f $X=-0.05 $Y=0 $X2=4.505 $Y2=2.59
cc_77 N_GND_M1014_b N_CK_c_579_n 0.0345662f $X=-0.05 $Y=0 $X2=4.36 $Y2=2.59
cc_78 N_GND_M1014_b N_CK_c_580_n 0.00714094f $X=-0.05 $Y=0 $X2=2.42 $Y2=2.59
cc_79 N_GND_M1014_b N_CK_c_581_n 0.0181831f $X=-0.05 $Y=0 $X2=5.355 $Y2=2.59
cc_80 N_GND_M1014_b N_CK_c_582_n 0.0041728f $X=-0.05 $Y=0 $X2=4.65 $Y2=2.59
cc_81 N_GND_M1014_b CK 0.00236135f $X=-0.05 $Y=0 $X2=5.5 $Y2=2.59
cc_82 N_GND_M1014_b N_A_27_115#_M1022_g 0.0171814f $X=-0.05 $Y=0 $X2=3.175
+ $Y2=1.075
cc_83 N_GND_c_42_p N_A_27_115#_M1022_g 0.00606474f $X=3.305 $Y=0.152 $X2=3.175
+ $Y2=1.075
cc_84 N_GND_c_22_p N_A_27_115#_M1022_g 0.00354579f $X=3.39 $Y=0.825 $X2=3.175
+ $Y2=1.075
cc_85 N_GND_c_3_p N_A_27_115#_M1022_g 0.00468827f $X=7.815 $Y=0.19 $X2=3.175
+ $Y2=1.075
cc_86 N_GND_M1014_b N_A_27_115#_c_776_n 0.0240953f $X=-0.05 $Y=0 $X2=3.53
+ $Y2=1.85
cc_87 N_GND_c_22_p N_A_27_115#_c_776_n 8.07204e-19 $X=3.39 $Y=0.825 $X2=3.53
+ $Y2=1.85
cc_88 N_GND_M1014_b N_A_27_115#_c_778_n 0.0105855f $X=-0.05 $Y=0 $X2=3.25
+ $Y2=1.85
cc_89 N_GND_M1014_b N_A_27_115#_c_779_n 0.0232417f $X=-0.05 $Y=0 $X2=3.53
+ $Y2=2.765
cc_90 N_GND_M1014_b N_A_27_115#_c_780_n 0.0105265f $X=-0.05 $Y=0 $X2=3.25
+ $Y2=2.765
cc_91 N_GND_M1014_b N_A_27_115#_M1015_g 0.0163216f $X=-0.05 $Y=0 $X2=3.605
+ $Y2=1.075
cc_92 N_GND_c_22_p N_A_27_115#_M1015_g 0.00354579f $X=3.39 $Y=0.825 $X2=3.605
+ $Y2=1.075
cc_93 N_GND_c_61_p N_A_27_115#_M1015_g 0.00606474f $X=5.055 $Y=0.152 $X2=3.605
+ $Y2=1.075
cc_94 N_GND_c_3_p N_A_27_115#_M1015_g 0.00468827f $X=7.815 $Y=0.19 $X2=3.605
+ $Y2=1.075
cc_95 N_GND_M1014_b N_A_27_115#_c_785_n 0.00155645f $X=-0.05 $Y=0 $X2=0.26
+ $Y2=0.825
cc_96 N_GND_c_2_p N_A_27_115#_c_785_n 0.00728471f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_97 N_GND_c_3_p N_A_27_115#_c_785_n 0.00474053f $X=7.815 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_98 N_GND_M1014_b N_A_27_115#_c_788_n 0.0155204f $X=-0.05 $Y=0 $X2=0.69
+ $Y2=1.85
cc_99 N_GND_M1014_b N_A_27_115#_c_789_n 0.00871176f $X=-0.05 $Y=0 $X2=3.345
+ $Y2=2.765
cc_100 N_GND_M1014_b N_A_27_115#_c_790_n 0.00245573f $X=-0.05 $Y=0 $X2=3.345
+ $Y2=1.85
cc_101 N_GND_c_22_p N_A_27_115#_c_790_n 0.00177942f $X=3.39 $Y=0.825 $X2=3.345
+ $Y2=1.85
cc_102 N_GND_M1014_b N_A_27_115#_c_792_n 0.0341069f $X=-0.05 $Y=0 $X2=3.11
+ $Y2=1.85
cc_103 N_GND_M1014_b N_A_27_115#_c_793_n 0.0023707f $X=-0.05 $Y=0 $X2=0.835
+ $Y2=1.85
cc_104 N_GND_M1014_b N_A_428_89#_c_899_n 0.0173059f $X=-0.05 $Y=0 $X2=2.215
+ $Y2=1.685
cc_105 N_GND_c_42_p N_A_428_89#_c_899_n 0.00606474f $X=3.305 $Y=0.152 $X2=2.215
+ $Y2=1.685
cc_106 N_GND_c_3_p N_A_428_89#_c_899_n 0.00468827f $X=7.815 $Y=0.19 $X2=2.215
+ $Y2=1.685
cc_107 N_GND_M1014_b N_A_428_89#_c_902_n 0.0203057f $X=-0.05 $Y=0 $X2=2.335
+ $Y2=2.225
cc_108 N_GND_M1014_b N_A_428_89#_c_903_n 0.0187566f $X=-0.05 $Y=0 $X2=2.74
+ $Y2=2.3
cc_109 N_GND_M1014_b N_A_428_89#_c_904_n 0.00755029f $X=-0.05 $Y=0 $X2=2.41
+ $Y2=2.3
cc_110 N_GND_M1014_b N_A_428_89#_M1019_g 0.032457f $X=-0.05 $Y=0 $X2=2.815
+ $Y2=4.585
cc_111 N_GND_M1014_b N_A_428_89#_c_906_n 0.0559794f $X=-0.05 $Y=0 $X2=3.89
+ $Y2=2.3
cc_112 N_GND_M1014_b N_A_428_89#_M1013_g 0.0319667f $X=-0.05 $Y=0 $X2=3.965
+ $Y2=4.585
cc_113 N_GND_M1014_b N_A_428_89#_c_908_n 0.0270462f $X=-0.05 $Y=0 $X2=4.37
+ $Y2=2.3
cc_114 N_GND_M1014_b N_A_428_89#_c_909_n 0.0125754f $X=-0.05 $Y=0 $X2=4.445
+ $Y2=2.225
cc_115 N_GND_M1014_b N_A_428_89#_c_910_n 0.0141451f $X=-0.05 $Y=0 $X2=2.335
+ $Y2=1.76
cc_116 N_GND_M1014_b N_A_428_89#_c_911_n 0.00426512f $X=-0.05 $Y=0 $X2=2.815
+ $Y2=2.3
cc_117 N_GND_M1014_b N_A_428_89#_c_912_n 0.00426512f $X=-0.05 $Y=0 $X2=3.965
+ $Y2=2.3
cc_118 N_GND_M1014_b N_A_428_89#_c_913_n 0.0256431f $X=-0.05 $Y=0 $X2=4.505
+ $Y2=1.85
cc_119 N_GND_M1014_b N_A_428_89#_c_914_n 0.01755f $X=-0.05 $Y=0 $X2=4.505
+ $Y2=1.685
cc_120 N_GND_c_61_p N_A_428_89#_c_914_n 0.00606474f $X=5.055 $Y=0.152 $X2=4.505
+ $Y2=1.685
cc_121 N_GND_c_3_p N_A_428_89#_c_914_n 0.00468827f $X=7.815 $Y=0.19 $X2=4.505
+ $Y2=1.685
cc_122 N_GND_M1014_b N_A_428_89#_c_917_n 0.0116005f $X=-0.05 $Y=0 $X2=5.485
+ $Y2=1.85
cc_123 N_GND_c_23_p N_A_428_89#_c_917_n 0.00564434f $X=5.14 $Y=0.825 $X2=5.485
+ $Y2=1.85
cc_124 N_GND_M1014_b N_A_428_89#_c_919_n 0.00549177f $X=-0.05 $Y=0 $X2=5.57
+ $Y2=0.825
cc_125 N_GND_c_23_p N_A_428_89#_c_919_n 4.65312e-19 $X=5.14 $Y=0.825 $X2=5.57
+ $Y2=0.825
cc_126 N_GND_c_6_p N_A_428_89#_c_919_n 0.00747016f $X=6.795 $Y=0.152 $X2=5.57
+ $Y2=0.825
cc_127 N_GND_c_3_p N_A_428_89#_c_919_n 0.00476261f $X=7.815 $Y=0.19 $X2=5.57
+ $Y2=0.825
cc_128 N_GND_M1014_b N_A_428_89#_c_923_n 0.0046852f $X=-0.05 $Y=0 $X2=5.57
+ $Y2=2.165
cc_129 N_GND_M1014_b N_A_428_89#_c_924_n 0.0131399f $X=-0.05 $Y=0 $X2=5.845
+ $Y2=3.1
cc_130 N_GND_M1014_b N_A_428_89#_c_925_n 8.79856e-19 $X=-0.05 $Y=0 $X2=5.57
+ $Y2=1.85
cc_131 N_GND_M1014_b N_A_428_89#_c_926_n 0.0128476f $X=-0.05 $Y=0 $X2=5.845
+ $Y2=2.25
cc_132 N_GND_M1014_b N_A_970_89#_M1008_g 0.0319752f $X=-0.05 $Y=0 $X2=4.925
+ $Y2=1.075
cc_133 N_GND_c_61_p N_A_970_89#_M1008_g 0.00606474f $X=5.055 $Y=0.152 $X2=4.925
+ $Y2=1.075
cc_134 N_GND_c_23_p N_A_970_89#_M1008_g 0.00360474f $X=5.14 $Y=0.825 $X2=4.925
+ $Y2=1.075
cc_135 N_GND_c_3_p N_A_970_89#_M1008_g 0.00468827f $X=7.815 $Y=0.19 $X2=4.925
+ $Y2=1.075
cc_136 N_GND_M1014_b N_A_970_89#_M1009_g 0.0330331f $X=-0.05 $Y=0 $X2=4.925
+ $Y2=4.585
cc_137 N_GND_M1014_b N_A_970_89#_c_1092_n 0.0263191f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=2.19
cc_138 N_GND_M1014_b N_A_970_89#_c_1093_n 0.0292185f $X=-0.05 $Y=0 $X2=7.57
+ $Y2=2.19
cc_139 N_GND_M1014_b N_A_970_89#_c_1094_n 0.0154776f $X=-0.05 $Y=0 $X2=7.572
+ $Y2=2.025
cc_140 N_GND_M1014_b N_A_970_89#_c_1095_n 0.0170508f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=1.65
cc_141 N_GND_c_7_p N_A_970_89#_c_1095_n 0.00380101f $X=6.88 $Y=0.825 $X2=7.66
+ $Y2=1.65
cc_142 N_GND_c_142_p N_A_970_89#_c_1095_n 0.00606474f $X=7.815 $Y=0.152 $X2=7.66
+ $Y2=1.65
cc_143 N_GND_c_143_p N_A_970_89#_c_1095_n 0.00354579f $X=7.9 $Y=0.825 $X2=7.66
+ $Y2=1.65
cc_144 N_GND_c_3_p N_A_970_89#_c_1095_n 0.00468827f $X=7.815 $Y=0.19 $X2=7.66
+ $Y2=1.65
cc_145 N_GND_M1014_b N_A_970_89#_c_1100_n 0.0140996f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=1.8
cc_146 N_GND_M1014_b N_A_970_89#_c_1101_n 0.0365245f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=2.855
cc_147 N_GND_M1014_b N_A_970_89#_c_1102_n 0.00495925f $X=-0.05 $Y=0 $X2=7.66
+ $Y2=3.005
cc_148 N_GND_M1014_b N_A_970_89#_c_1103_n 0.00396219f $X=-0.05 $Y=0 $X2=4.985
+ $Y2=2.19
cc_149 N_GND_M1014_b N_A_970_89#_c_1104_n 0.00155645f $X=-0.05 $Y=0 $X2=6.09
+ $Y2=0.825
cc_150 N_GND_c_6_p N_A_970_89#_c_1104_n 0.00750025f $X=6.795 $Y=0.152 $X2=6.09
+ $Y2=0.825
cc_151 N_GND_c_3_p N_A_970_89#_c_1104_n 0.00474053f $X=7.815 $Y=0.19 $X2=6.09
+ $Y2=0.825
cc_152 N_GND_M1014_b N_A_970_89#_c_1107_n 0.0109395f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=2.105
cc_153 N_GND_M1014_b N_A_970_89#_c_1108_n 0.0140059f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=4.815
cc_154 N_GND_M1014_b N_A_970_89#_c_1109_n 0.0189667f $X=-0.05 $Y=0 $X2=7.57
+ $Y2=2.19
cc_155 N_GND_M1014_b N_A_970_89#_c_1110_n 0.00193448f $X=-0.05 $Y=0 $X2=6.52
+ $Y2=2.19
cc_156 N_GND_M1014_b N_A_970_89#_c_1111_n 0.0581721f $X=-0.05 $Y=0 $X2=7.425
+ $Y2=2.19
cc_157 N_GND_M1014_b N_A_970_89#_c_1112_n 0.0017195f $X=-0.05 $Y=0 $X2=5.13
+ $Y2=2.19
cc_158 N_GND_M1014_b N_A_970_89#_c_1113_n 0.00173636f $X=-0.05 $Y=0 $X2=7.57
+ $Y2=2.19
cc_159 N_GND_M1014_b N_A_808_115#_M1007_g 0.0367887f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=0.945
cc_160 N_GND_c_6_p N_A_808_115#_M1007_g 0.00606474f $X=6.795 $Y=0.152 $X2=6.305
+ $Y2=0.945
cc_161 N_GND_c_3_p N_A_808_115#_M1007_g 0.00468827f $X=7.815 $Y=0.19 $X2=6.305
+ $Y2=0.945
cc_162 N_GND_M1014_b N_A_808_115#_M1020_g 0.0548413f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=5.085
cc_163 N_GND_M1014_b N_A_808_115#_c_1255_n 0.0460049f $X=-0.05 $Y=0 $X2=6.305
+ $Y2=1.85
cc_164 N_GND_M1014_b N_A_808_115#_c_1256_n 0.0112983f $X=-0.05 $Y=0 $X2=3.685
+ $Y2=1.85
cc_165 N_GND_M1014_b N_A_808_115#_c_1257_n 0.00313975f $X=-0.05 $Y=0 $X2=4.265
+ $Y2=0.825
cc_166 N_GND_c_61_p N_A_808_115#_c_1257_n 0.014959f $X=5.055 $Y=0.152 $X2=4.265
+ $Y2=0.825
cc_167 N_GND_c_3_p N_A_808_115#_c_1257_n 0.00958198f $X=7.815 $Y=0.19 $X2=4.265
+ $Y2=0.825
cc_168 N_GND_M1014_b N_A_808_115#_c_1260_n 0.00161958f $X=-0.05 $Y=0 $X2=6.1
+ $Y2=1.85
cc_169 N_GND_M1014_b N_A_808_115#_c_1261_n 0.0204013f $X=-0.05 $Y=0 $X2=5.955
+ $Y2=1.85
cc_170 N_GND_c_23_p N_A_808_115#_c_1261_n 5.03331e-19 $X=5.14 $Y=0.825 $X2=5.955
+ $Y2=1.85
cc_171 N_GND_M1014_b N_A_808_115#_c_1263_n 0.00120467f $X=-0.05 $Y=0 $X2=3.83
+ $Y2=1.85
cc_172 N_GND_M1014_b N_A_808_115#_c_1264_n 6.71961e-19 $X=-0.05 $Y=0 $X2=6.1
+ $Y2=1.85
cc_173 N_GND_M1014_b N_QN_M1028_g 0.0561552f $X=-0.05 $Y=0 $X2=8.115 $Y2=1.075
cc_174 N_GND_c_143_p N_QN_M1028_g 0.00354579f $X=7.9 $Y=0.825 $X2=8.115
+ $Y2=1.075
cc_175 N_GND_c_3_p N_QN_M1028_g 0.00468827f $X=7.815 $Y=0.19 $X2=8.115 $Y2=1.075
cc_176 N_GND_M1014_b N_QN_M1029_g 0.0186095f $X=-0.05 $Y=0 $X2=8.115 $Y2=4.585
cc_177 N_GND_M1014_b N_QN_c_1383_n 0.0291912f $X=-0.05 $Y=0 $X2=8.055 $Y2=2.395
cc_178 N_GND_M1014_b N_QN_c_1384_n 0.00514305f $X=-0.05 $Y=0 $X2=7.47 $Y2=0.825
cc_179 N_GND_c_7_p N_QN_c_1384_n 0.0186519f $X=6.88 $Y=0.825 $X2=7.47 $Y2=0.825
cc_180 N_GND_c_142_p N_QN_c_1384_n 0.00757793f $X=7.815 $Y=0.152 $X2=7.47
+ $Y2=0.825
cc_181 N_GND_c_3_p N_QN_c_1384_n 0.00476261f $X=7.815 $Y=0.19 $X2=7.47 $Y2=0.825
cc_182 N_GND_M1014_b N_QN_c_1388_n 0.00138285f $X=-0.05 $Y=0 $X2=7.47 $Y2=2.96
cc_183 N_GND_M1014_b N_QN_c_1389_n 0.0171269f $X=-0.05 $Y=0 $X2=7.97 $Y2=1.85
cc_184 N_GND_M1014_b N_QN_c_1390_n 0.00371251f $X=-0.05 $Y=0 $X2=7.555 $Y2=1.85
cc_185 N_GND_M1014_b N_QN_c_1391_n 0.0176115f $X=-0.05 $Y=0 $X2=7.97 $Y2=2.765
cc_186 N_GND_M1014_b N_QN_c_1392_n 0.00426693f $X=-0.05 $Y=0 $X2=7.555 $Y2=2.765
cc_187 N_GND_M1014_b N_QN_c_1393_n 0.0034889f $X=-0.05 $Y=0 $X2=8.055 $Y2=2.395
cc_188 N_GND_M1014_b QN 0.0029781f $X=-0.05 $Y=0 $X2=7.475 $Y2=2.96
cc_189 N_GND_M1014_b N_Q_c_1464_n 0.00913846f $X=-0.05 $Y=0 $X2=8.33 $Y2=0.825
cc_190 N_GND_c_3_p N_Q_c_1464_n 0.00476261f $X=7.815 $Y=0.19 $X2=8.33 $Y2=0.825
cc_191 N_GND_M1014_b N_Q_c_1466_n 0.0625704f $X=-0.05 $Y=0 $X2=8.445 $Y2=3.16
cc_192 N_GND_M1014_b N_Q_c_1467_n 0.0140324f $X=-0.05 $Y=0 $X2=8.445 $Y2=1.515
cc_193 N_VDD_M1026_b N_SN_M1026_g 0.107741f $X=-0.05 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_194 N_VDD_c_194_p N_SN_M1026_g 0.00713292f $X=0.26 $Y=4.815 $X2=0.475
+ $Y2=5.085
cc_195 N_VDD_c_195_p N_SN_M1026_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475
+ $Y2=5.085
cc_196 N_VDD_c_196_p N_SN_M1026_g 0.00468827f $X=7.815 $Y=6.47 $X2=0.475
+ $Y2=5.085
cc_197 N_VDD_M1026_b N_SN_M1021_g 0.0872322f $X=-0.05 $Y=2.905 $X2=6.735
+ $Y2=5.085
cc_198 N_VDD_c_198_p N_SN_M1021_g 0.00606474f $X=6.865 $Y=6.507 $X2=6.735
+ $Y2=5.085
cc_199 N_VDD_c_199_p N_SN_M1021_g 0.00713292f $X=6.95 $Y=4.815 $X2=6.735
+ $Y2=5.085
cc_200 N_VDD_c_196_p N_SN_M1021_g 0.00468827f $X=7.815 $Y=6.47 $X2=6.735
+ $Y2=5.085
cc_201 N_VDD_M1026_b N_A_152_89#_M1017_g 0.0915939f $X=-0.05 $Y=2.905 $X2=0.905
+ $Y2=5.085
cc_202 N_VDD_c_195_p N_A_152_89#_M1017_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905
+ $Y2=5.085
cc_203 N_VDD_c_203_p N_A_152_89#_M1017_g 0.00713292f $X=1.12 $Y=4.815 $X2=0.905
+ $Y2=5.085
cc_204 N_VDD_c_204_p N_A_152_89#_M1017_g 0.026288f $X=1.64 $Y=3.795 $X2=0.905
+ $Y2=5.085
cc_205 N_VDD_c_196_p N_A_152_89#_M1017_g 0.00468827f $X=7.815 $Y=6.47 $X2=0.905
+ $Y2=5.085
cc_206 N_VDD_M1026_b N_A_152_89#_c_434_n 0.00286294f $X=-0.05 $Y=2.905 $X2=1.03
+ $Y2=2.305
cc_207 N_VDD_M1002_s N_A_152_89#_c_450_n 0.0125004f $X=1.515 $Y=3.085 $X2=2.345
+ $Y2=3.185
cc_208 N_VDD_M1026_b N_A_152_89#_c_450_n 0.0286398f $X=-0.05 $Y=2.905 $X2=2.345
+ $Y2=3.185
cc_209 N_VDD_c_204_p N_A_152_89#_c_450_n 0.00952036f $X=1.64 $Y=3.795 $X2=2.345
+ $Y2=3.185
cc_210 N_VDD_M1026_b N_A_152_89#_c_453_n 0.00545748f $X=-0.05 $Y=2.905 $X2=1.115
+ $Y2=3.185
cc_211 N_VDD_M1026_b N_A_152_89#_c_454_n 0.00313975f $X=-0.05 $Y=2.905 $X2=2.515
+ $Y2=3.455
cc_212 N_VDD_c_212_p N_A_152_89#_c_454_n 0.0149461f $X=3.305 $Y=6.507 $X2=2.515
+ $Y2=3.455
cc_213 N_VDD_c_196_p N_A_152_89#_c_454_n 0.00958198f $X=7.815 $Y=6.47 $X2=2.515
+ $Y2=3.455
cc_214 N_VDD_M1026_b N_D_M1002_g 0.0222869f $X=-0.05 $Y=2.905 $X2=1.855
+ $Y2=4.585
cc_215 N_VDD_c_204_p N_D_M1002_g 0.00713292f $X=1.64 $Y=3.795 $X2=1.855
+ $Y2=4.585
cc_216 N_VDD_c_212_p N_D_M1002_g 0.00606474f $X=3.305 $Y=6.507 $X2=1.855
+ $Y2=4.585
cc_217 N_VDD_c_196_p N_D_M1002_g 0.00468827f $X=7.815 $Y=6.47 $X2=1.855
+ $Y2=4.585
cc_218 N_VDD_M1026_b N_CK_M1025_g 0.020128f $X=-0.05 $Y=2.905 $X2=2.215
+ $Y2=4.585
cc_219 N_VDD_c_212_p N_CK_M1025_g 0.00606474f $X=3.305 $Y=6.507 $X2=2.215
+ $Y2=4.585
cc_220 N_VDD_c_196_p N_CK_M1025_g 0.00468827f $X=7.815 $Y=6.47 $X2=2.215
+ $Y2=4.585
cc_221 N_VDD_M1026_b N_CK_M1005_g 0.020128f $X=-0.05 $Y=2.905 $X2=4.565
+ $Y2=4.585
cc_222 N_VDD_c_222_p N_CK_M1005_g 0.00606474f $X=5.055 $Y=6.507 $X2=4.565
+ $Y2=4.585
cc_223 N_VDD_c_196_p N_CK_M1005_g 0.00468827f $X=7.815 $Y=6.47 $X2=4.565
+ $Y2=4.585
cc_224 N_VDD_M1026_b N_CK_c_554_n 0.00774555f $X=-0.05 $Y=2.905 $X2=5.355
+ $Y2=2.93
cc_225 N_VDD_M1026_b N_CK_M1006_g 0.0214648f $X=-0.05 $Y=2.905 $X2=5.355
+ $Y2=4.585
cc_226 N_VDD_c_226_p N_CK_M1006_g 0.00354579f $X=5.14 $Y=3.455 $X2=5.355
+ $Y2=4.585
cc_227 N_VDD_c_227_p N_CK_M1006_g 0.00606474f $X=6.005 $Y=6.507 $X2=5.355
+ $Y2=4.585
cc_228 N_VDD_c_228_p N_CK_M1006_g 0.00603096f $X=6.09 $Y=4.815 $X2=5.355
+ $Y2=4.585
cc_229 N_VDD_c_196_p N_CK_M1006_g 0.00468827f $X=7.815 $Y=6.47 $X2=5.355
+ $Y2=4.585
cc_230 N_VDD_M1026_b N_CK_c_556_n 0.00487135f $X=-0.05 $Y=2.905 $X2=2.275
+ $Y2=2.765
cc_231 N_VDD_M1026_b N_CK_c_565_n 0.00487051f $X=-0.05 $Y=2.905 $X2=4.505
+ $Y2=2.765
cc_232 N_VDD_M1026_b N_CK_c_576_n 0.00302835f $X=-0.05 $Y=2.905 $X2=5.5 $Y2=2.59
cc_233 N_VDD_M1026_b N_CK_c_577_n 6.42499e-19 $X=-0.05 $Y=2.905 $X2=2.275
+ $Y2=2.59
cc_234 N_VDD_M1026_b N_CK_c_578_n 0.0022456f $X=-0.05 $Y=2.905 $X2=4.505
+ $Y2=2.59
cc_235 N_VDD_c_226_p N_CK_c_581_n 0.00634153f $X=5.14 $Y=3.455 $X2=5.355
+ $Y2=2.59
cc_236 N_VDD_M1026_b N_A_27_115#_M1023_g 0.0192219f $X=-0.05 $Y=2.905 $X2=3.175
+ $Y2=4.585
cc_237 N_VDD_c_212_p N_A_27_115#_M1023_g 0.00606474f $X=3.305 $Y=6.507 $X2=3.175
+ $Y2=4.585
cc_238 N_VDD_c_238_p N_A_27_115#_M1023_g 0.00354579f $X=3.39 $Y=3.795 $X2=3.175
+ $Y2=4.585
cc_239 N_VDD_c_196_p N_A_27_115#_M1023_g 0.00468827f $X=7.815 $Y=6.47 $X2=3.175
+ $Y2=4.585
cc_240 N_VDD_c_238_p N_A_27_115#_c_779_n 8.24975e-19 $X=3.39 $Y=3.795 $X2=3.53
+ $Y2=2.765
cc_241 N_VDD_M1026_b N_A_27_115#_M1016_g 0.0181098f $X=-0.05 $Y=2.905 $X2=3.605
+ $Y2=4.585
cc_242 N_VDD_c_238_p N_A_27_115#_M1016_g 0.00354579f $X=3.39 $Y=3.795 $X2=3.605
+ $Y2=4.585
cc_243 N_VDD_c_222_p N_A_27_115#_M1016_g 0.00606474f $X=5.055 $Y=6.507 $X2=3.605
+ $Y2=4.585
cc_244 N_VDD_c_196_p N_A_27_115#_M1016_g 0.00468827f $X=7.815 $Y=6.47 $X2=3.605
+ $Y2=4.585
cc_245 N_VDD_M1026_b N_A_27_115#_c_788_n 0.0289135f $X=-0.05 $Y=2.905 $X2=0.69
+ $Y2=1.85
cc_246 N_VDD_c_195_p N_A_27_115#_c_788_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69
+ $Y2=1.85
cc_247 N_VDD_c_196_p N_A_27_115#_c_788_n 0.00475776f $X=7.815 $Y=6.47 $X2=0.69
+ $Y2=1.85
cc_248 N_VDD_M1026_b N_A_27_115#_c_789_n 0.00424346f $X=-0.05 $Y=2.905 $X2=3.345
+ $Y2=2.765
cc_249 N_VDD_c_238_p N_A_27_115#_c_789_n 0.004428f $X=3.39 $Y=3.795 $X2=3.345
+ $Y2=2.765
cc_250 N_VDD_M1026_b N_A_428_89#_M1019_g 0.0215131f $X=-0.05 $Y=2.905 $X2=2.815
+ $Y2=4.585
cc_251 N_VDD_c_212_p N_A_428_89#_M1019_g 0.00606474f $X=3.305 $Y=6.507 $X2=2.815
+ $Y2=4.585
cc_252 N_VDD_c_196_p N_A_428_89#_M1019_g 0.00468827f $X=7.815 $Y=6.47 $X2=2.815
+ $Y2=4.585
cc_253 N_VDD_M1026_b N_A_428_89#_M1013_g 0.0214821f $X=-0.05 $Y=2.905 $X2=3.965
+ $Y2=4.585
cc_254 N_VDD_c_222_p N_A_428_89#_M1013_g 0.00606474f $X=5.055 $Y=6.507 $X2=3.965
+ $Y2=4.585
cc_255 N_VDD_c_196_p N_A_428_89#_M1013_g 0.00468827f $X=7.815 $Y=6.47 $X2=3.965
+ $Y2=4.585
cc_256 N_VDD_M1026_b N_A_428_89#_c_933_n 0.00156053f $X=-0.05 $Y=2.905 $X2=5.57
+ $Y2=3.455
cc_257 N_VDD_c_227_p N_A_428_89#_c_933_n 0.00747016f $X=6.005 $Y=6.507 $X2=5.57
+ $Y2=3.455
cc_258 N_VDD_c_228_p N_A_428_89#_c_933_n 0.064932f $X=6.09 $Y=4.815 $X2=5.57
+ $Y2=3.455
cc_259 N_VDD_c_196_p N_A_428_89#_c_933_n 0.00476261f $X=7.815 $Y=6.47 $X2=5.57
+ $Y2=3.455
cc_260 N_VDD_M1026_b N_A_428_89#_c_924_n 0.00560125f $X=-0.05 $Y=2.905 $X2=5.845
+ $Y2=3.1
cc_261 N_VDD_M1026_b N_A_428_89#_c_938_n 0.0139078f $X=-0.05 $Y=2.905 $X2=5.845
+ $Y2=3.185
cc_262 N_VDD_M1026_b N_A_970_89#_M1009_g 0.0197647f $X=-0.05 $Y=2.905 $X2=4.925
+ $Y2=4.585
cc_263 N_VDD_c_222_p N_A_970_89#_M1009_g 0.00606474f $X=5.055 $Y=6.507 $X2=4.925
+ $Y2=4.585
cc_264 N_VDD_c_226_p N_A_970_89#_M1009_g 0.00354579f $X=5.14 $Y=3.455 $X2=4.925
+ $Y2=4.585
cc_265 N_VDD_c_196_p N_A_970_89#_M1009_g 0.00468827f $X=7.815 $Y=6.47 $X2=4.925
+ $Y2=4.585
cc_266 N_VDD_M1026_b N_A_970_89#_c_1102_n 0.0266934f $X=-0.05 $Y=2.905 $X2=7.66
+ $Y2=3.005
cc_267 N_VDD_c_199_p N_A_970_89#_c_1102_n 0.00603096f $X=6.95 $Y=4.815 $X2=7.66
+ $Y2=3.005
cc_268 N_VDD_c_268_p N_A_970_89#_c_1102_n 0.00606474f $X=7.815 $Y=6.507 $X2=7.66
+ $Y2=3.005
cc_269 N_VDD_c_269_p N_A_970_89#_c_1102_n 0.00354579f $X=7.9 $Y=4.475 $X2=7.66
+ $Y2=3.005
cc_270 N_VDD_c_196_p N_A_970_89#_c_1102_n 0.00468827f $X=7.815 $Y=6.47 $X2=7.66
+ $Y2=3.005
cc_271 N_VDD_M1026_b N_A_970_89#_c_1108_n 0.0294479f $X=-0.05 $Y=2.905 $X2=6.52
+ $Y2=4.815
cc_272 N_VDD_c_198_p N_A_970_89#_c_1108_n 0.00734006f $X=6.865 $Y=6.507 $X2=6.52
+ $Y2=4.815
cc_273 N_VDD_c_196_p N_A_970_89#_c_1108_n 0.00475776f $X=7.815 $Y=6.47 $X2=6.52
+ $Y2=4.815
cc_274 N_VDD_M1026_b N_A_808_115#_M1020_g 0.0852884f $X=-0.05 $Y=2.905 $X2=6.305
+ $Y2=5.085
cc_275 N_VDD_c_228_p N_A_808_115#_M1020_g 0.00713292f $X=6.09 $Y=4.815 $X2=6.305
+ $Y2=5.085
cc_276 N_VDD_c_198_p N_A_808_115#_M1020_g 0.00606474f $X=6.865 $Y=6.507
+ $X2=6.305 $Y2=5.085
cc_277 N_VDD_c_196_p N_A_808_115#_M1020_g 0.00468827f $X=7.815 $Y=6.47 $X2=6.305
+ $Y2=5.085
cc_278 N_VDD_M1026_b N_A_808_115#_c_1256_n 0.00168314f $X=-0.05 $Y=2.905
+ $X2=3.685 $Y2=1.85
cc_279 N_VDD_M1026_b N_A_808_115#_c_1270_n 0.00313975f $X=-0.05 $Y=2.905
+ $X2=4.265 $Y2=3.795
cc_280 N_VDD_c_222_p N_A_808_115#_c_1270_n 0.014959f $X=5.055 $Y=6.507 $X2=4.265
+ $Y2=3.795
cc_281 N_VDD_c_196_p N_A_808_115#_c_1270_n 0.00958198f $X=7.815 $Y=6.47
+ $X2=4.265 $Y2=3.795
cc_282 N_VDD_M1026_b N_QN_M1029_g 0.0248218f $X=-0.05 $Y=2.905 $X2=8.115
+ $Y2=4.585
cc_283 N_VDD_c_269_p N_QN_M1029_g 0.00354579f $X=7.9 $Y=4.475 $X2=8.115
+ $Y2=4.585
cc_284 N_VDD_c_284_p N_QN_M1029_g 0.00606474f $X=7.815 $Y=6.47 $X2=8.115
+ $Y2=4.585
cc_285 N_VDD_c_196_p N_QN_M1029_g 0.00468827f $X=7.815 $Y=6.47 $X2=8.115
+ $Y2=4.585
cc_286 N_VDD_M1026_b N_QN_c_1388_n 0.00648064f $X=-0.05 $Y=2.905 $X2=7.47
+ $Y2=2.96
cc_287 N_VDD_c_199_p N_QN_c_1388_n 0.064932f $X=6.95 $Y=4.815 $X2=7.47 $Y2=2.96
cc_288 N_VDD_c_268_p N_QN_c_1388_n 0.00757793f $X=7.815 $Y=6.507 $X2=7.47
+ $Y2=2.96
cc_289 N_VDD_c_196_p N_QN_c_1388_n 0.00476261f $X=7.815 $Y=6.47 $X2=7.47
+ $Y2=2.96
cc_290 N_VDD_M1026_b QN 0.0110667f $X=-0.05 $Y=2.905 $X2=7.475 $Y2=2.96
cc_291 N_VDD_M1026_b N_Q_c_1468_n 0.00156053f $X=-0.05 $Y=2.905 $X2=8.33
+ $Y2=4.475
cc_292 N_VDD_c_284_p N_Q_c_1468_n 0.00757793f $X=7.815 $Y=6.47 $X2=8.33
+ $Y2=4.475
cc_293 N_VDD_c_196_p N_Q_c_1468_n 0.00476261f $X=7.815 $Y=6.47 $X2=8.33
+ $Y2=4.475
cc_294 N_VDD_M1026_b N_Q_c_1466_n 0.0117744f $X=-0.05 $Y=2.905 $X2=8.445
+ $Y2=3.16
cc_295 N_VDD_M1026_b N_Q_c_1472_n 0.0093035f $X=-0.05 $Y=2.905 $X2=8.33
+ $Y2=3.287
cc_296 N_VDD_M1026_b Q 0.00503768f $X=-0.05 $Y=2.905 $X2=8.325 $Y2=3.33
cc_297 N_SN_c_312_n N_A_152_89#_M1024_d 0.00558831f $X=6.715 $Y=1.48 $X2=2.29
+ $Y2=0.575
cc_298 N_SN_M1014_g N_A_152_89#_M1000_g 0.0617259f $X=0.475 $Y=0.945 $X2=0.835
+ $Y2=0.945
cc_299 N_SN_c_309_n N_A_152_89#_M1000_g 5.71653e-19 $X=0.32 $Y=1.48 $X2=0.835
+ $Y2=0.945
cc_300 N_SN_c_312_n N_A_152_89#_M1000_g 0.0100323f $X=6.715 $Y=1.48 $X2=0.835
+ $Y2=0.945
cc_301 N_SN_M1026_g N_A_152_89#_M1017_g 0.0825015f $X=0.475 $Y=5.085 $X2=0.905
+ $Y2=5.085
cc_302 N_SN_c_306_n N_A_152_89#_c_433_n 0.0617259f $X=0.32 $Y=1.85 $X2=1.03
+ $Y2=2.305
cc_303 N_SN_c_312_n N_A_152_89#_c_435_n 0.0293336f $X=6.715 $Y=1.48 $X2=2.33
+ $Y2=1.765
cc_304 N_SN_c_312_n N_A_152_89#_c_438_n 0.00320514f $X=6.715 $Y=1.48 $X2=1.115
+ $Y2=1.765
cc_305 N_SN_c_312_n N_A_152_89#_c_440_n 0.0151351f $X=6.715 $Y=1.48 $X2=2.415
+ $Y2=1.68
cc_306 N_SN_c_312_n N_A_152_89#_c_466_n 0.0254135f $X=6.715 $Y=1.48 $X2=2.507
+ $Y2=1.415
cc_307 N_SN_c_312_n N_D_M1001_g 0.0116357f $X=6.715 $Y=1.48 $X2=1.855 $Y2=1.075
cc_308 N_SN_c_312_n N_CK_c_557_n 8.06574e-19 $X=6.715 $Y=1.48 $X2=2.755 $Y2=1.85
cc_309 N_SN_c_312_n N_CK_c_558_n 0.0106495f $X=6.715 $Y=1.48 $X2=2.755 $Y2=1.685
cc_310 N_SN_c_312_n N_CK_c_561_n 8.06574e-19 $X=6.715 $Y=1.48 $X2=4.025 $Y2=1.85
cc_311 N_SN_c_312_n N_CK_c_562_n 0.00177838f $X=6.715 $Y=1.48 $X2=4.025
+ $Y2=1.685
cc_312 N_SN_c_312_n N_CK_c_566_n 0.01159f $X=6.715 $Y=1.48 $X2=5.382 $Y2=1.685
cc_313 N_SN_c_312_n N_CK_c_570_n 0.00107886f $X=6.715 $Y=1.48 $X2=5.382
+ $Y2=1.835
cc_314 N_SN_c_312_n N_CK_c_572_n 0.00496158f $X=6.715 $Y=1.48 $X2=2.755 $Y2=1.85
cc_315 N_SN_c_312_n N_CK_c_573_n 0.00118606f $X=6.715 $Y=1.48 $X2=4.025 $Y2=1.85
cc_316 N_SN_c_312_n N_A_27_115#_M1022_g 0.0104272f $X=6.715 $Y=1.48 $X2=3.175
+ $Y2=1.075
cc_317 N_SN_c_312_n N_A_27_115#_c_776_n 2.42482e-19 $X=6.715 $Y=1.48 $X2=3.53
+ $Y2=1.85
cc_318 N_SN_c_312_n N_A_27_115#_M1015_g 0.00491871f $X=6.715 $Y=1.48 $X2=3.605
+ $Y2=1.075
cc_319 N_SN_M1014_g N_A_27_115#_c_811_n 0.0152601f $X=0.475 $Y=0.945 $X2=0.605
+ $Y2=1.08
cc_320 N_SN_c_309_n N_A_27_115#_c_811_n 0.00168015f $X=0.32 $Y=1.48 $X2=0.605
+ $Y2=1.08
cc_321 N_SN_c_312_n N_A_27_115#_c_811_n 0.00543257f $X=6.715 $Y=1.48 $X2=0.605
+ $Y2=1.08
cc_322 N_SN_c_320_n N_A_27_115#_c_811_n 0.00396192f $X=0.465 $Y=1.48 $X2=0.605
+ $Y2=1.08
cc_323 N_SN_c_306_n N_A_27_115#_c_815_n 0.00199006f $X=0.32 $Y=1.85 $X2=0.345
+ $Y2=1.08
cc_324 N_SN_c_309_n N_A_27_115#_c_815_n 0.0057346f $X=0.32 $Y=1.48 $X2=0.345
+ $Y2=1.08
cc_325 N_SN_c_320_n N_A_27_115#_c_815_n 0.00629987f $X=0.465 $Y=1.48 $X2=0.345
+ $Y2=1.08
cc_326 N_SN_M1014_g N_A_27_115#_c_788_n 0.05751f $X=0.475 $Y=0.945 $X2=0.69
+ $Y2=1.85
cc_327 N_SN_c_309_n N_A_27_115#_c_788_n 0.0352919f $X=0.32 $Y=1.48 $X2=0.69
+ $Y2=1.85
cc_328 N_SN_c_312_n N_A_27_115#_c_788_n 0.0203124f $X=6.715 $Y=1.48 $X2=0.69
+ $Y2=1.85
cc_329 N_SN_c_320_n N_A_27_115#_c_788_n 0.00217814f $X=0.465 $Y=1.48 $X2=0.69
+ $Y2=1.85
cc_330 N_SN_c_312_n N_A_27_115#_c_790_n 0.00546464f $X=6.715 $Y=1.48 $X2=3.345
+ $Y2=1.85
cc_331 N_SN_c_312_n N_A_27_115#_c_792_n 0.183238f $X=6.715 $Y=1.48 $X2=3.11
+ $Y2=1.85
cc_332 N_SN_c_306_n N_A_27_115#_c_793_n 0.00336449f $X=0.32 $Y=1.85 $X2=0.835
+ $Y2=1.85
cc_333 N_SN_c_309_n N_A_27_115#_c_793_n 0.00667526f $X=0.32 $Y=1.48 $X2=0.835
+ $Y2=1.85
cc_334 N_SN_c_312_n N_A_27_115#_c_793_n 0.02527f $X=6.715 $Y=1.48 $X2=0.835
+ $Y2=1.85
cc_335 N_SN_c_312_n N_A_27_115#_c_827_n 0.0259207f $X=6.715 $Y=1.48 $X2=3.255
+ $Y2=1.85
cc_336 N_SN_c_312_n N_A_428_89#_M1004_d 0.0042281f $X=6.715 $Y=1.48 $X2=5.43
+ $Y2=0.575
cc_337 N_SN_c_312_n N_A_428_89#_c_899_n 0.0102209f $X=6.715 $Y=1.48 $X2=2.215
+ $Y2=1.685
cc_338 N_SN_c_312_n N_A_428_89#_c_913_n 0.00232964f $X=6.715 $Y=1.48 $X2=4.505
+ $Y2=1.85
cc_339 N_SN_c_312_n N_A_428_89#_c_914_n 0.0103799f $X=6.715 $Y=1.48 $X2=4.505
+ $Y2=1.685
cc_340 N_SN_c_312_n N_A_428_89#_c_917_n 0.0115848f $X=6.715 $Y=1.48 $X2=5.485
+ $Y2=1.85
cc_341 N_SN_c_312_n N_A_428_89#_c_919_n 0.0255624f $X=6.715 $Y=1.48 $X2=5.57
+ $Y2=0.825
cc_342 N_SN_c_312_n N_A_428_89#_c_926_n 4.57217e-19 $X=6.715 $Y=1.48 $X2=5.845
+ $Y2=2.25
cc_343 N_SN_c_312_n N_A_970_89#_M1008_g 0.0100216f $X=6.715 $Y=1.48 $X2=4.925
+ $Y2=1.075
cc_344 N_SN_M1021_g N_A_970_89#_c_1093_n 0.00575596f $X=6.735 $Y=5.085 $X2=7.57
+ $Y2=2.19
cc_345 N_SN_c_307_n N_A_970_89#_c_1095_n 0.00315793f $X=6.735 $Y=1.59 $X2=7.66
+ $Y2=1.65
cc_346 N_SN_c_307_n N_A_970_89#_c_1100_n 0.00149674f $X=6.735 $Y=1.59 $X2=7.66
+ $Y2=1.8
cc_347 N_SN_c_301_n N_A_970_89#_c_1130_n 0.00722422f $X=6.665 $Y=1.425 $X2=6.435
+ $Y2=1.08
cc_348 N_SN_c_312_n N_A_970_89#_c_1130_n 0.00902188f $X=6.715 $Y=1.48 $X2=6.435
+ $Y2=1.08
cc_349 N_SN_c_312_n N_A_970_89#_c_1132_n 0.00539675f $X=6.715 $Y=1.48 $X2=6.175
+ $Y2=1.08
cc_350 N_SN_c_301_n N_A_970_89#_c_1107_n 0.00996282f $X=6.665 $Y=1.425 $X2=6.52
+ $Y2=2.105
cc_351 N_SN_c_307_n N_A_970_89#_c_1107_n 0.01362f $X=6.735 $Y=1.59 $X2=6.52
+ $Y2=2.105
cc_352 N_SN_c_310_n N_A_970_89#_c_1107_n 0.0239974f $X=6.86 $Y=1.48 $X2=6.52
+ $Y2=2.105
cc_353 N_SN_c_312_n N_A_970_89#_c_1107_n 0.0235322f $X=6.715 $Y=1.48 $X2=6.52
+ $Y2=2.105
cc_354 N_SN_c_321_n N_A_970_89#_c_1107_n 0.00211162f $X=6.86 $Y=1.48 $X2=6.52
+ $Y2=2.105
cc_355 N_SN_M1021_g N_A_970_89#_c_1108_n 0.04564f $X=6.735 $Y=5.085 $X2=6.52
+ $Y2=4.815
cc_356 N_SN_M1021_g N_A_970_89#_c_1109_n 0.0140836f $X=6.735 $Y=5.085 $X2=7.57
+ $Y2=2.19
cc_357 N_SN_c_307_n N_A_970_89#_c_1109_n 0.00352021f $X=6.735 $Y=1.59 $X2=7.57
+ $Y2=2.19
cc_358 N_SN_c_310_n N_A_970_89#_c_1109_n 0.00510357f $X=6.86 $Y=1.48 $X2=7.57
+ $Y2=2.19
cc_359 N_SN_c_312_n N_A_970_89#_c_1109_n 9.00052e-19 $X=6.715 $Y=1.48 $X2=7.57
+ $Y2=2.19
cc_360 N_SN_c_321_n N_A_970_89#_c_1109_n 0.00126364f $X=6.86 $Y=1.48 $X2=7.57
+ $Y2=2.19
cc_361 N_SN_M1021_g N_A_970_89#_c_1111_n 0.00852135f $X=6.735 $Y=5.085 $X2=7.425
+ $Y2=2.19
cc_362 N_SN_c_307_n N_A_970_89#_c_1111_n 0.00176046f $X=6.735 $Y=1.59 $X2=7.425
+ $Y2=2.19
cc_363 N_SN_c_310_n N_A_970_89#_c_1111_n 0.00156423f $X=6.86 $Y=1.48 $X2=7.425
+ $Y2=2.19
cc_364 N_SN_c_312_n N_A_970_89#_c_1111_n 0.0209725f $X=6.715 $Y=1.48 $X2=7.425
+ $Y2=2.19
cc_365 N_SN_c_321_n N_A_970_89#_c_1111_n 0.01406f $X=6.86 $Y=1.48 $X2=7.425
+ $Y2=2.19
cc_366 N_SN_M1021_g N_A_970_89#_c_1113_n 7.50694e-19 $X=6.735 $Y=5.085 $X2=7.57
+ $Y2=2.19
cc_367 N_SN_c_312_n N_A_808_115#_M1012_d 0.0051762f $X=6.715 $Y=1.48 $X2=4.04
+ $Y2=0.575
cc_368 N_SN_c_301_n N_A_808_115#_M1007_g 0.074649f $X=6.665 $Y=1.425 $X2=6.305
+ $Y2=0.945
cc_369 N_SN_c_307_n N_A_808_115#_M1007_g 0.0567807f $X=6.735 $Y=1.59 $X2=6.305
+ $Y2=0.945
cc_370 N_SN_c_312_n N_A_808_115#_M1007_g 0.00802725f $X=6.715 $Y=1.48 $X2=6.305
+ $Y2=0.945
cc_371 N_SN_M1021_g N_A_808_115#_c_1255_n 0.0567807f $X=6.735 $Y=5.085 $X2=6.305
+ $Y2=1.85
cc_372 N_SN_c_312_n N_A_808_115#_c_1255_n 0.00412631f $X=6.715 $Y=1.48 $X2=6.305
+ $Y2=1.85
cc_373 N_SN_c_312_n N_A_808_115#_c_1256_n 0.00616681f $X=6.715 $Y=1.48 $X2=3.685
+ $Y2=1.85
cc_374 N_SN_c_312_n N_A_808_115#_c_1280_n 0.0537388f $X=6.715 $Y=1.48 $X2=4.095
+ $Y2=1.43
cc_375 N_SN_c_312_n N_A_808_115#_c_1281_n 0.0129425f $X=6.715 $Y=1.48 $X2=3.77
+ $Y2=1.43
cc_376 N_SN_c_312_n N_A_808_115#_c_1260_n 0.00274558f $X=6.715 $Y=1.48 $X2=6.1
+ $Y2=1.85
cc_377 N_SN_c_312_n N_A_808_115#_c_1261_n 0.176894f $X=6.715 $Y=1.48 $X2=5.955
+ $Y2=1.85
cc_378 N_SN_c_312_n N_A_808_115#_c_1263_n 0.0252354f $X=6.715 $Y=1.48 $X2=3.83
+ $Y2=1.85
cc_379 N_SN_c_312_n N_A_808_115#_c_1264_n 0.02673f $X=6.715 $Y=1.48 $X2=6.1
+ $Y2=1.85
cc_380 N_SN_c_301_n N_QN_c_1384_n 0.00771489f $X=6.665 $Y=1.425 $X2=7.47
+ $Y2=0.825
cc_381 N_SN_M1021_g N_QN_c_1384_n 2.02156e-19 $X=6.735 $Y=5.085 $X2=7.47
+ $Y2=0.825
cc_382 N_SN_c_307_n N_QN_c_1384_n 0.00252942f $X=6.735 $Y=1.59 $X2=7.47
+ $Y2=0.825
cc_383 N_SN_c_310_n N_QN_c_1384_n 0.00977948f $X=6.86 $Y=1.48 $X2=7.47 $Y2=0.825
cc_384 N_SN_c_321_n N_QN_c_1384_n 0.00696569f $X=6.86 $Y=1.48 $X2=7.47 $Y2=0.825
cc_385 N_SN_M1021_g N_QN_c_1388_n 0.0405705f $X=6.735 $Y=5.085 $X2=7.47 $Y2=2.96
cc_386 N_SN_M1021_g N_QN_c_1390_n 0.00458451f $X=6.735 $Y=5.085 $X2=7.555
+ $Y2=1.85
cc_387 N_SN_M1021_g N_QN_c_1392_n 0.00454519f $X=6.735 $Y=5.085 $X2=7.555
+ $Y2=2.765
cc_388 N_SN_M1021_g QN 0.00491824f $X=6.735 $Y=5.085 $X2=7.475 $Y2=2.96
cc_389 N_SN_c_312_n A_386_115# 0.00911585f $X=6.715 $Y=1.48 $X2=1.93 $Y2=0.575
cc_390 N_SN_c_312_n A_578_115# 0.0100396f $X=6.715 $Y=1.48 $X2=2.89 $Y2=0.575
cc_391 N_SN_c_312_n A_736_115# 0.00106636f $X=6.715 $Y=1.48 $X2=3.68 $Y2=0.575
cc_392 N_SN_c_312_n A_928_115# 0.00917995f $X=6.715 $Y=1.48 $X2=4.64 $Y2=0.575
cc_393 N_A_152_89#_c_434_n N_D_M1001_g 0.00508967f $X=1.03 $Y=2.305 $X2=1.855
+ $Y2=1.075
cc_394 N_A_152_89#_c_435_n N_D_M1001_g 0.0123125f $X=2.33 $Y=1.765 $X2=1.855
+ $Y2=1.075
cc_395 N_A_152_89#_c_434_n N_D_M1002_g 0.0129373f $X=1.03 $Y=2.305 $X2=1.855
+ $Y2=4.585
cc_396 N_A_152_89#_c_450_n N_D_M1002_g 0.0211938f $X=2.345 $Y=3.185 $X2=1.855
+ $Y2=4.585
cc_397 N_A_152_89#_c_433_n N_D_c_518_n 0.00628944f $X=1.03 $Y=2.305 $X2=1.915
+ $Y2=2.22
cc_398 N_A_152_89#_c_434_n N_D_c_518_n 0.00131071f $X=1.03 $Y=2.305 $X2=1.915
+ $Y2=2.22
cc_399 N_A_152_89#_c_435_n N_D_c_518_n 0.00207628f $X=2.33 $Y=1.765 $X2=1.915
+ $Y2=2.22
cc_400 N_A_152_89#_c_433_n N_D_c_519_n 0.00168445f $X=1.03 $Y=2.305 $X2=1.915
+ $Y2=2.22
cc_401 N_A_152_89#_c_435_n N_D_c_519_n 0.0086486f $X=2.33 $Y=1.765 $X2=1.915
+ $Y2=2.22
cc_402 N_A_152_89#_c_433_n D 0.00279288f $X=1.03 $Y=2.305 $X2=1.915 $Y2=2.22
cc_403 N_A_152_89#_c_435_n D 0.00200799f $X=2.33 $Y=1.765 $X2=1.915 $Y2=2.22
cc_404 N_A_152_89#_c_450_n N_CK_M1025_g 0.0153421f $X=2.345 $Y=3.185 $X2=2.215
+ $Y2=4.585
cc_405 N_A_152_89#_c_450_n N_CK_c_556_n 0.00150627f $X=2.345 $Y=3.185 $X2=2.275
+ $Y2=2.765
cc_406 N_A_152_89#_c_435_n N_CK_c_557_n 9.45214e-19 $X=2.33 $Y=1.765 $X2=2.755
+ $Y2=1.85
cc_407 N_A_152_89#_c_466_n N_CK_c_557_n 0.00170561f $X=2.507 $Y=1.415 $X2=2.755
+ $Y2=1.85
cc_408 N_A_152_89#_c_440_n N_CK_c_558_n 0.00464203f $X=2.415 $Y=1.68 $X2=2.755
+ $Y2=1.685
cc_409 N_A_152_89#_c_466_n N_CK_c_558_n 0.00545632f $X=2.507 $Y=1.415 $X2=2.755
+ $Y2=1.685
cc_410 N_A_152_89#_c_435_n N_CK_c_571_n 0.0019742f $X=2.33 $Y=1.765 $X2=2.67
+ $Y2=2.59
cc_411 N_A_152_89#_c_450_n N_CK_c_571_n 0.00883015f $X=2.345 $Y=3.185 $X2=2.67
+ $Y2=2.59
cc_412 N_A_152_89#_c_435_n N_CK_c_572_n 0.012316f $X=2.33 $Y=1.765 $X2=2.755
+ $Y2=1.85
cc_413 N_A_152_89#_c_466_n N_CK_c_572_n 5.28119e-19 $X=2.507 $Y=1.415 $X2=2.755
+ $Y2=1.85
cc_414 N_A_152_89#_c_435_n N_CK_c_577_n 0.00224444f $X=2.33 $Y=1.765 $X2=2.275
+ $Y2=2.59
cc_415 N_A_152_89#_c_450_n N_CK_c_577_n 0.0101098f $X=2.345 $Y=3.185 $X2=2.275
+ $Y2=2.59
cc_416 N_A_152_89#_c_450_n N_CK_c_579_n 0.00601583f $X=2.345 $Y=3.185 $X2=4.36
+ $Y2=2.59
cc_417 N_A_152_89#_c_450_n N_CK_c_580_n 0.00409373f $X=2.345 $Y=3.185 $X2=2.42
+ $Y2=2.59
cc_418 N_A_152_89#_M1000_g N_A_27_115#_c_811_n 0.00722422f $X=0.835 $Y=0.945
+ $X2=0.605 $Y2=1.08
cc_419 N_A_152_89#_M1000_g N_A_27_115#_c_788_n 0.0264927f $X=0.835 $Y=0.945
+ $X2=0.69 $Y2=1.85
cc_420 N_A_152_89#_M1017_g N_A_27_115#_c_788_n 0.0274967f $X=0.905 $Y=5.085
+ $X2=0.69 $Y2=1.85
cc_421 N_A_152_89#_c_433_n N_A_27_115#_c_788_n 0.00720273f $X=1.03 $Y=2.305
+ $X2=0.69 $Y2=1.85
cc_422 N_A_152_89#_c_434_n N_A_27_115#_c_788_n 0.0874214f $X=1.03 $Y=2.305
+ $X2=0.69 $Y2=1.85
cc_423 N_A_152_89#_c_438_n N_A_27_115#_c_788_n 0.0124515f $X=1.115 $Y=1.765
+ $X2=0.69 $Y2=1.85
cc_424 N_A_152_89#_c_453_n N_A_27_115#_c_788_n 0.013584f $X=1.115 $Y=3.185
+ $X2=0.69 $Y2=1.85
cc_425 N_A_152_89#_M1000_g N_A_27_115#_c_792_n 0.0065801f $X=0.835 $Y=0.945
+ $X2=3.11 $Y2=1.85
cc_426 N_A_152_89#_c_433_n N_A_27_115#_c_792_n 0.00224331f $X=1.03 $Y=2.305
+ $X2=3.11 $Y2=1.85
cc_427 N_A_152_89#_c_434_n N_A_27_115#_c_792_n 0.00977499f $X=1.03 $Y=2.305
+ $X2=3.11 $Y2=1.85
cc_428 N_A_152_89#_c_435_n N_A_27_115#_c_792_n 0.0532053f $X=2.33 $Y=1.765
+ $X2=3.11 $Y2=1.85
cc_429 N_A_152_89#_c_438_n N_A_27_115#_c_792_n 0.00403513f $X=1.115 $Y=1.765
+ $X2=3.11 $Y2=1.85
cc_430 N_A_152_89#_c_466_n N_A_27_115#_c_792_n 8.61924e-19 $X=2.507 $Y=1.415
+ $X2=3.11 $Y2=1.85
cc_431 N_A_152_89#_M1000_g N_A_27_115#_c_793_n 0.00343239f $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=1.85
cc_432 N_A_152_89#_c_434_n N_A_27_115#_c_793_n 8.0088e-19 $X=1.03 $Y=2.305
+ $X2=0.835 $Y2=1.85
cc_433 N_A_152_89#_c_438_n N_A_27_115#_c_793_n 8.3209e-19 $X=1.115 $Y=1.765
+ $X2=0.835 $Y2=1.85
cc_434 N_A_152_89#_c_435_n N_A_428_89#_c_899_n 0.0022787f $X=2.33 $Y=1.765
+ $X2=2.215 $Y2=1.685
cc_435 N_A_152_89#_c_466_n N_A_428_89#_c_899_n 0.0060945f $X=2.507 $Y=1.415
+ $X2=2.215 $Y2=1.685
cc_436 N_A_152_89#_c_435_n N_A_428_89#_c_902_n 0.00324141f $X=2.33 $Y=1.765
+ $X2=2.335 $Y2=2.225
cc_437 N_A_152_89#_c_435_n N_A_428_89#_c_910_n 0.00993431f $X=2.33 $Y=1.765
+ $X2=2.335 $Y2=1.76
cc_438 N_A_152_89#_c_450_n A_386_617# 0.00732587f $X=2.345 $Y=3.185 $X2=1.93
+ $Y2=3.085
cc_439 N_D_M1002_g N_CK_c_556_n 0.21604f $X=1.855 $Y=4.585 $X2=2.275 $Y2=2.765
cc_440 N_D_c_518_n N_CK_c_572_n 2.89615e-19 $X=1.915 $Y=2.22 $X2=2.755 $Y2=1.85
cc_441 N_D_c_519_n N_CK_c_572_n 0.00478177f $X=1.915 $Y=2.22 $X2=2.755 $Y2=1.85
cc_442 D N_CK_c_572_n 0.00551577f $X=1.915 $Y=2.22 $X2=2.755 $Y2=1.85
cc_443 N_D_M1002_g N_CK_c_577_n 0.00494364f $X=1.855 $Y=4.585 $X2=2.275 $Y2=2.59
cc_444 N_D_M1002_g N_CK_c_580_n 0.00515433f $X=1.855 $Y=4.585 $X2=2.42 $Y2=2.59
cc_445 D N_CK_c_580_n 0.00375733f $X=1.915 $Y=2.22 $X2=2.42 $Y2=2.59
cc_446 N_D_M1001_g N_A_27_115#_c_792_n 0.0030176f $X=1.855 $Y=1.075 $X2=3.11
+ $Y2=1.85
cc_447 N_D_c_518_n N_A_27_115#_c_792_n 7.9412e-19 $X=1.915 $Y=2.22 $X2=3.11
+ $Y2=1.85
cc_448 N_D_c_519_n N_A_27_115#_c_792_n 0.00111625f $X=1.915 $Y=2.22 $X2=3.11
+ $Y2=1.85
cc_449 D N_A_27_115#_c_792_n 0.0353362f $X=1.915 $Y=2.22 $X2=3.11 $Y2=1.85
cc_450 N_D_M1001_g N_A_428_89#_c_899_n 0.0846533f $X=1.855 $Y=1.075 $X2=2.215
+ $Y2=1.685
cc_451 N_D_M1001_g N_A_428_89#_c_902_n 0.00932846f $X=1.855 $Y=1.075 $X2=2.335
+ $Y2=2.225
cc_452 N_D_c_518_n N_A_428_89#_c_902_n 0.0210215f $X=1.915 $Y=2.22 $X2=2.335
+ $Y2=2.225
cc_453 N_D_c_519_n N_A_428_89#_c_902_n 0.00164409f $X=1.915 $Y=2.22 $X2=2.335
+ $Y2=2.225
cc_454 D N_A_428_89#_c_902_n 0.00342011f $X=1.915 $Y=2.22 $X2=2.335 $Y2=2.225
cc_455 D N_A_428_89#_c_904_n 4.62757e-19 $X=1.915 $Y=2.22 $X2=2.41 $Y2=2.3
cc_456 N_CK_c_558_n N_A_27_115#_M1022_g 0.0483944f $X=2.755 $Y=1.685 $X2=3.175
+ $Y2=1.075
cc_457 N_CK_c_572_n N_A_27_115#_M1022_g 0.00109079f $X=2.755 $Y=1.85 $X2=3.175
+ $Y2=1.075
cc_458 N_CK_c_561_n N_A_27_115#_c_776_n 0.0473482f $X=4.025 $Y=1.85 $X2=3.53
+ $Y2=1.85
cc_459 N_CK_c_557_n N_A_27_115#_c_778_n 0.0483944f $X=2.755 $Y=1.85 $X2=3.25
+ $Y2=1.85
cc_460 N_CK_c_579_n N_A_27_115#_c_779_n 0.00772879f $X=4.36 $Y=2.59 $X2=3.53
+ $Y2=2.765
cc_461 N_CK_c_579_n N_A_27_115#_c_780_n 0.00679967f $X=4.36 $Y=2.59 $X2=3.25
+ $Y2=2.765
cc_462 N_CK_c_562_n N_A_27_115#_M1015_g 0.0473482f $X=4.025 $Y=1.685 $X2=3.605
+ $Y2=1.075
cc_463 N_CK_c_573_n N_A_27_115#_M1015_g 3.67139e-19 $X=4.025 $Y=1.85 $X2=3.605
+ $Y2=1.075
cc_464 N_CK_c_557_n N_A_27_115#_c_789_n 7.30049e-19 $X=2.755 $Y=1.85 $X2=3.345
+ $Y2=2.765
cc_465 N_CK_c_571_n N_A_27_115#_c_789_n 0.00401809f $X=2.67 $Y=2.59 $X2=3.345
+ $Y2=2.765
cc_466 N_CK_c_572_n N_A_27_115#_c_789_n 0.0203851f $X=2.755 $Y=1.85 $X2=3.345
+ $Y2=2.765
cc_467 N_CK_c_579_n N_A_27_115#_c_789_n 0.0206884f $X=4.36 $Y=2.59 $X2=3.345
+ $Y2=2.765
cc_468 N_CK_c_557_n N_A_27_115#_c_790_n 7.18106e-19 $X=2.755 $Y=1.85 $X2=3.345
+ $Y2=1.85
cc_469 N_CK_c_572_n N_A_27_115#_c_790_n 0.00742068f $X=2.755 $Y=1.85 $X2=3.345
+ $Y2=1.85
cc_470 N_CK_c_579_n N_A_27_115#_c_790_n 0.00102309f $X=4.36 $Y=2.59 $X2=3.345
+ $Y2=1.85
cc_471 N_CK_c_557_n N_A_27_115#_c_792_n 0.00383172f $X=2.755 $Y=1.85 $X2=3.11
+ $Y2=1.85
cc_472 N_CK_c_571_n N_A_27_115#_c_792_n 0.00443421f $X=2.67 $Y=2.59 $X2=3.11
+ $Y2=1.85
cc_473 N_CK_c_572_n N_A_27_115#_c_792_n 0.0149977f $X=2.755 $Y=1.85 $X2=3.11
+ $Y2=1.85
cc_474 N_CK_c_577_n N_A_27_115#_c_792_n 7.12046e-19 $X=2.275 $Y=2.59 $X2=3.11
+ $Y2=1.85
cc_475 N_CK_c_580_n N_A_27_115#_c_792_n 0.0126164f $X=2.42 $Y=2.59 $X2=3.11
+ $Y2=1.85
cc_476 N_CK_c_557_n N_A_27_115#_c_827_n 3.3031e-19 $X=2.755 $Y=1.85 $X2=3.255
+ $Y2=1.85
cc_477 N_CK_c_572_n N_A_27_115#_c_827_n 0.00143592f $X=2.755 $Y=1.85 $X2=3.255
+ $Y2=1.85
cc_478 N_CK_c_579_n N_A_27_115#_c_827_n 0.0129652f $X=4.36 $Y=2.59 $X2=3.255
+ $Y2=1.85
cc_479 N_CK_c_558_n N_A_428_89#_c_899_n 0.0252931f $X=2.755 $Y=1.685 $X2=2.215
+ $Y2=1.685
cc_480 N_CK_c_572_n N_A_428_89#_c_902_n 0.00613747f $X=2.755 $Y=1.85 $X2=2.335
+ $Y2=2.225
cc_481 N_CK_c_557_n N_A_428_89#_c_903_n 0.0183603f $X=2.755 $Y=1.85 $X2=2.74
+ $Y2=2.3
cc_482 N_CK_c_572_n N_A_428_89#_c_903_n 0.00630484f $X=2.755 $Y=1.85 $X2=2.74
+ $Y2=2.3
cc_483 N_CK_c_579_n N_A_428_89#_c_903_n 0.00613485f $X=4.36 $Y=2.59 $X2=2.74
+ $Y2=2.3
cc_484 N_CK_c_556_n N_A_428_89#_c_904_n 0.00904036f $X=2.275 $Y=2.765 $X2=2.41
+ $Y2=2.3
cc_485 N_CK_c_571_n N_A_428_89#_c_904_n 0.00878348f $X=2.67 $Y=2.59 $X2=2.41
+ $Y2=2.3
cc_486 N_CK_c_577_n N_A_428_89#_c_904_n 0.00109468f $X=2.275 $Y=2.59 $X2=2.41
+ $Y2=2.3
cc_487 N_CK_c_580_n N_A_428_89#_c_904_n 0.00137501f $X=2.42 $Y=2.59 $X2=2.41
+ $Y2=2.3
cc_488 N_CK_M1025_g N_A_428_89#_M1019_g 0.0612221f $X=2.215 $Y=4.585 $X2=2.815
+ $Y2=4.585
cc_489 N_CK_c_556_n N_A_428_89#_M1019_g 0.0128384f $X=2.275 $Y=2.765 $X2=2.815
+ $Y2=4.585
cc_490 N_CK_c_571_n N_A_428_89#_M1019_g 0.0081071f $X=2.67 $Y=2.59 $X2=2.815
+ $Y2=4.585
cc_491 N_CK_c_572_n N_A_428_89#_M1019_g 0.00478024f $X=2.755 $Y=1.85 $X2=2.815
+ $Y2=4.585
cc_492 N_CK_c_577_n N_A_428_89#_M1019_g 0.00184124f $X=2.275 $Y=2.59 $X2=2.815
+ $Y2=4.585
cc_493 N_CK_c_579_n N_A_428_89#_M1019_g 0.00938974f $X=4.36 $Y=2.59 $X2=2.815
+ $Y2=4.585
cc_494 N_CK_c_580_n N_A_428_89#_M1019_g 4.2e-19 $X=2.42 $Y=2.59 $X2=2.815
+ $Y2=4.585
cc_495 N_CK_c_579_n N_A_428_89#_c_906_n 0.00607908f $X=4.36 $Y=2.59 $X2=3.89
+ $Y2=2.3
cc_496 N_CK_M1005_g N_A_428_89#_M1013_g 0.0612221f $X=4.565 $Y=4.585 $X2=3.965
+ $Y2=4.585
cc_497 N_CK_c_565_n N_A_428_89#_M1013_g 0.0118393f $X=4.505 $Y=2.765 $X2=3.965
+ $Y2=4.585
cc_498 N_CK_c_573_n N_A_428_89#_M1013_g 0.00399495f $X=4.025 $Y=1.85 $X2=3.965
+ $Y2=4.585
cc_499 N_CK_c_575_n N_A_428_89#_M1013_g 0.00654233f $X=4.11 $Y=2.59 $X2=3.965
+ $Y2=4.585
cc_500 N_CK_c_578_n N_A_428_89#_M1013_g 0.00128351f $X=4.505 $Y=2.59 $X2=3.965
+ $Y2=4.585
cc_501 N_CK_c_579_n N_A_428_89#_M1013_g 0.00497421f $X=4.36 $Y=2.59 $X2=3.965
+ $Y2=4.585
cc_502 N_CK_c_582_n N_A_428_89#_M1013_g 4.2e-19 $X=4.65 $Y=2.59 $X2=3.965
+ $Y2=4.585
cc_503 N_CK_c_565_n N_A_428_89#_c_908_n 0.00904036f $X=4.505 $Y=2.765 $X2=4.37
+ $Y2=2.3
cc_504 N_CK_c_573_n N_A_428_89#_c_908_n 0.00909647f $X=4.025 $Y=1.85 $X2=4.37
+ $Y2=2.3
cc_505 N_CK_c_574_n N_A_428_89#_c_908_n 0.00924811f $X=4.42 $Y=2.59 $X2=4.37
+ $Y2=2.3
cc_506 N_CK_c_578_n N_A_428_89#_c_908_n 0.00102633f $X=4.505 $Y=2.59 $X2=4.37
+ $Y2=2.3
cc_507 N_CK_c_579_n N_A_428_89#_c_908_n 0.00613485f $X=4.36 $Y=2.59 $X2=4.37
+ $Y2=2.3
cc_508 N_CK_c_582_n N_A_428_89#_c_908_n 0.00137501f $X=4.65 $Y=2.59 $X2=4.37
+ $Y2=2.3
cc_509 N_CK_c_573_n N_A_428_89#_c_909_n 0.00649764f $X=4.025 $Y=1.85 $X2=4.445
+ $Y2=2.225
cc_510 N_CK_c_557_n N_A_428_89#_c_910_n 0.0216263f $X=2.755 $Y=1.85 $X2=2.335
+ $Y2=1.76
cc_511 N_CK_c_577_n N_A_428_89#_c_910_n 2.45465e-19 $X=2.275 $Y=2.59 $X2=2.335
+ $Y2=1.76
cc_512 N_CK_c_572_n N_A_428_89#_c_911_n 0.00568091f $X=2.755 $Y=1.85 $X2=2.815
+ $Y2=2.3
cc_513 N_CK_c_561_n N_A_428_89#_c_912_n 0.0183603f $X=4.025 $Y=1.85 $X2=3.965
+ $Y2=2.3
cc_514 N_CK_c_573_n N_A_428_89#_c_912_n 0.00436024f $X=4.025 $Y=1.85 $X2=3.965
+ $Y2=2.3
cc_515 N_CK_c_561_n N_A_428_89#_c_913_n 0.0220721f $X=4.025 $Y=1.85 $X2=4.505
+ $Y2=1.85
cc_516 N_CK_c_565_n N_A_428_89#_c_913_n 0.00227671f $X=4.505 $Y=2.765 $X2=4.505
+ $Y2=1.85
cc_517 N_CK_c_573_n N_A_428_89#_c_913_n 0.00131283f $X=4.025 $Y=1.85 $X2=4.505
+ $Y2=1.85
cc_518 N_CK_c_578_n N_A_428_89#_c_913_n 5.27321e-19 $X=4.505 $Y=2.59 $X2=4.505
+ $Y2=1.85
cc_519 N_CK_c_582_n N_A_428_89#_c_913_n 8.78837e-19 $X=4.65 $Y=2.59 $X2=4.505
+ $Y2=1.85
cc_520 N_CK_c_562_n N_A_428_89#_c_914_n 0.0268981f $X=4.025 $Y=1.685 $X2=4.505
+ $Y2=1.685
cc_521 N_CK_c_555_n N_A_428_89#_c_917_n 0.00592387f $X=5.41 $Y=2.6 $X2=5.485
+ $Y2=1.85
cc_522 N_CK_c_561_n N_A_428_89#_c_917_n 8.05876e-19 $X=4.025 $Y=1.85 $X2=5.485
+ $Y2=1.85
cc_523 N_CK_c_565_n N_A_428_89#_c_917_n 5.56676e-19 $X=4.505 $Y=2.765 $X2=5.485
+ $Y2=1.85
cc_524 N_CK_c_570_n N_A_428_89#_c_917_n 0.00762848f $X=5.382 $Y=1.835 $X2=5.485
+ $Y2=1.85
cc_525 N_CK_c_573_n N_A_428_89#_c_917_n 0.00853323f $X=4.025 $Y=1.85 $X2=5.485
+ $Y2=1.85
cc_526 N_CK_c_574_n N_A_428_89#_c_917_n 0.00132011f $X=4.42 $Y=2.59 $X2=5.485
+ $Y2=1.85
cc_527 N_CK_c_576_n N_A_428_89#_c_917_n 8.24249e-19 $X=5.5 $Y=2.59 $X2=5.485
+ $Y2=1.85
cc_528 N_CK_c_578_n N_A_428_89#_c_917_n 0.00261697f $X=4.505 $Y=2.59 $X2=5.485
+ $Y2=1.85
cc_529 N_CK_c_579_n N_A_428_89#_c_917_n 3.12599e-19 $X=4.36 $Y=2.59 $X2=5.485
+ $Y2=1.85
cc_530 N_CK_c_581_n N_A_428_89#_c_917_n 0.00341454f $X=5.355 $Y=2.59 $X2=5.485
+ $Y2=1.85
cc_531 N_CK_c_582_n N_A_428_89#_c_917_n 0.00221563f $X=4.65 $Y=2.59 $X2=5.485
+ $Y2=1.85
cc_532 N_CK_c_566_n N_A_428_89#_c_919_n 0.0102351f $X=5.382 $Y=1.685 $X2=5.57
+ $Y2=0.825
cc_533 N_CK_c_570_n N_A_428_89#_c_919_n 0.0022869f $X=5.382 $Y=1.835 $X2=5.57
+ $Y2=0.825
cc_534 N_CK_c_555_n N_A_428_89#_c_923_n 0.00735778f $X=5.41 $Y=2.6 $X2=5.57
+ $Y2=2.165
cc_535 N_CK_c_554_n N_A_428_89#_c_924_n 0.00333903f $X=5.355 $Y=2.93 $X2=5.845
+ $Y2=3.1
cc_536 N_CK_M1006_g N_A_428_89#_c_924_n 0.00495264f $X=5.355 $Y=4.585 $X2=5.845
+ $Y2=3.1
cc_537 N_CK_c_555_n N_A_428_89#_c_924_n 0.00567067f $X=5.41 $Y=2.6 $X2=5.845
+ $Y2=3.1
cc_538 N_CK_c_576_n N_A_428_89#_c_924_n 0.0289277f $X=5.5 $Y=2.59 $X2=5.845
+ $Y2=3.1
cc_539 CK N_A_428_89#_c_924_n 0.00852929f $X=5.5 $Y=2.59 $X2=5.845 $Y2=3.1
cc_540 N_CK_c_555_n N_A_428_89#_c_925_n 0.00114916f $X=5.41 $Y=2.6 $X2=5.57
+ $Y2=1.85
cc_541 N_CK_c_570_n N_A_428_89#_c_925_n 8.09104e-19 $X=5.382 $Y=1.835 $X2=5.57
+ $Y2=1.85
cc_542 N_CK_c_554_n N_A_428_89#_c_926_n 0.00198338f $X=5.355 $Y=2.93 $X2=5.845
+ $Y2=2.25
cc_543 N_CK_c_555_n N_A_428_89#_c_926_n 0.00559872f $X=5.41 $Y=2.6 $X2=5.845
+ $Y2=2.25
cc_544 N_CK_c_576_n N_A_428_89#_c_926_n 0.00661696f $X=5.5 $Y=2.59 $X2=5.845
+ $Y2=2.25
cc_545 CK N_A_428_89#_c_926_n 0.00236431f $X=5.5 $Y=2.59 $X2=5.845 $Y2=2.25
cc_546 N_CK_c_554_n N_A_428_89#_c_938_n 0.00260941f $X=5.355 $Y=2.93 $X2=5.845
+ $Y2=3.185
cc_547 N_CK_c_576_n N_A_428_89#_c_938_n 0.00706443f $X=5.5 $Y=2.59 $X2=5.845
+ $Y2=3.185
cc_548 CK N_A_428_89#_c_938_n 0.00259785f $X=5.5 $Y=2.59 $X2=5.845 $Y2=3.185
cc_549 N_CK_c_555_n N_A_970_89#_M1008_g 0.00697006f $X=5.41 $Y=2.6 $X2=4.925
+ $Y2=1.075
cc_550 N_CK_c_566_n N_A_970_89#_M1008_g 0.0287519f $X=5.382 $Y=1.685 $X2=4.925
+ $Y2=1.075
cc_551 N_CK_c_554_n N_A_970_89#_M1009_g 0.0287701f $X=5.355 $Y=2.93 $X2=4.925
+ $Y2=4.585
cc_552 N_CK_c_555_n N_A_970_89#_M1009_g 0.0175925f $X=5.41 $Y=2.6 $X2=4.925
+ $Y2=4.585
cc_553 N_CK_c_565_n N_A_970_89#_M1009_g 0.214863f $X=4.505 $Y=2.765 $X2=4.925
+ $Y2=4.585
cc_554 N_CK_c_576_n N_A_970_89#_M1009_g 0.0026346f $X=5.5 $Y=2.59 $X2=4.925
+ $Y2=4.585
cc_555 N_CK_c_578_n N_A_970_89#_M1009_g 0.00453616f $X=4.505 $Y=2.59 $X2=4.925
+ $Y2=4.585
cc_556 N_CK_c_581_n N_A_970_89#_M1009_g 0.0114893f $X=5.355 $Y=2.59 $X2=4.925
+ $Y2=4.585
cc_557 N_CK_c_582_n N_A_970_89#_M1009_g 0.00113587f $X=4.65 $Y=2.59 $X2=4.925
+ $Y2=4.585
cc_558 CK N_A_970_89#_M1009_g 3.05655e-19 $X=5.5 $Y=2.59 $X2=4.925 $Y2=4.585
cc_559 N_CK_c_555_n N_A_970_89#_c_1092_n 0.0213116f $X=5.41 $Y=2.6 $X2=4.985
+ $Y2=2.19
cc_560 N_CK_c_581_n N_A_970_89#_c_1092_n 0.00185875f $X=5.355 $Y=2.59 $X2=4.985
+ $Y2=2.19
cc_561 N_CK_c_555_n N_A_970_89#_c_1103_n 9.0669e-19 $X=5.41 $Y=2.6 $X2=4.985
+ $Y2=2.19
cc_562 N_CK_c_581_n N_A_970_89#_c_1103_n 0.00488871f $X=5.355 $Y=2.59 $X2=4.985
+ $Y2=2.19
cc_563 N_CK_c_555_n N_A_970_89#_c_1111_n 0.00431553f $X=5.41 $Y=2.6 $X2=7.425
+ $Y2=2.19
cc_564 N_CK_c_576_n N_A_970_89#_c_1111_n 5.80133e-19 $X=5.5 $Y=2.59 $X2=7.425
+ $Y2=2.19
cc_565 N_CK_c_581_n N_A_970_89#_c_1111_n 0.0179446f $X=5.355 $Y=2.59 $X2=7.425
+ $Y2=2.19
cc_566 CK N_A_970_89#_c_1111_n 0.0240913f $X=5.5 $Y=2.59 $X2=7.425 $Y2=2.19
cc_567 N_CK_c_555_n N_A_970_89#_c_1112_n 8.66236e-19 $X=5.41 $Y=2.6 $X2=5.13
+ $Y2=2.19
cc_568 N_CK_c_581_n N_A_970_89#_c_1112_n 0.0247156f $X=5.355 $Y=2.59 $X2=5.13
+ $Y2=2.19
cc_569 N_CK_c_554_n N_A_808_115#_M1020_g 0.0044653f $X=5.355 $Y=2.93 $X2=6.305
+ $Y2=5.085
cc_570 N_CK_c_570_n N_A_808_115#_c_1255_n 0.00662135f $X=5.382 $Y=1.835
+ $X2=6.305 $Y2=1.85
cc_571 N_CK_c_562_n N_A_808_115#_c_1256_n 0.00554221f $X=4.025 $Y=1.685
+ $X2=3.685 $Y2=1.85
cc_572 N_CK_c_573_n N_A_808_115#_c_1256_n 0.057541f $X=4.025 $Y=1.85 $X2=3.685
+ $Y2=1.85
cc_573 N_CK_c_575_n N_A_808_115#_c_1256_n 0.0116326f $X=4.11 $Y=2.59 $X2=3.685
+ $Y2=1.85
cc_574 N_CK_c_578_n N_A_808_115#_c_1256_n 0.00613815f $X=4.505 $Y=2.59 $X2=3.685
+ $Y2=1.85
cc_575 N_CK_c_579_n N_A_808_115#_c_1256_n 0.020361f $X=4.36 $Y=2.59 $X2=3.685
+ $Y2=1.85
cc_576 N_CK_c_582_n N_A_808_115#_c_1256_n 6.61118e-19 $X=4.65 $Y=2.59 $X2=3.685
+ $Y2=1.85
cc_577 N_CK_c_561_n N_A_808_115#_c_1280_n 0.00227744f $X=4.025 $Y=1.85 $X2=4.095
+ $Y2=1.43
cc_578 N_CK_c_562_n N_A_808_115#_c_1280_n 0.0149609f $X=4.025 $Y=1.685 $X2=4.095
+ $Y2=1.43
cc_579 N_CK_c_573_n N_A_808_115#_c_1280_n 0.0103267f $X=4.025 $Y=1.85 $X2=4.095
+ $Y2=1.43
cc_580 N_CK_c_565_n N_A_808_115#_c_1297_n 0.00150627f $X=4.505 $Y=2.765
+ $X2=4.095 $Y2=3.185
cc_581 N_CK_c_574_n N_A_808_115#_c_1297_n 0.00843004f $X=4.42 $Y=2.59 $X2=4.095
+ $Y2=3.185
cc_582 N_CK_c_575_n N_A_808_115#_c_1297_n 0.00323798f $X=4.11 $Y=2.59 $X2=4.095
+ $Y2=3.185
cc_583 N_CK_c_578_n N_A_808_115#_c_1297_n 0.00103871f $X=4.505 $Y=2.59 $X2=4.095
+ $Y2=3.185
cc_584 N_CK_c_579_n N_A_808_115#_c_1297_n 0.012754f $X=4.36 $Y=2.59 $X2=4.095
+ $Y2=3.185
cc_585 N_CK_c_582_n N_A_808_115#_c_1297_n 0.00146098f $X=4.65 $Y=2.59 $X2=4.095
+ $Y2=3.185
cc_586 N_CK_c_570_n N_A_808_115#_c_1260_n 3.50905e-19 $X=5.382 $Y=1.835 $X2=6.1
+ $Y2=1.85
cc_587 N_CK_c_555_n N_A_808_115#_c_1261_n 0.00128484f $X=5.41 $Y=2.6 $X2=5.955
+ $Y2=1.85
cc_588 N_CK_c_561_n N_A_808_115#_c_1261_n 0.00362401f $X=4.025 $Y=1.85 $X2=5.955
+ $Y2=1.85
cc_589 N_CK_c_570_n N_A_808_115#_c_1261_n 0.00179204f $X=5.382 $Y=1.835
+ $X2=5.955 $Y2=1.85
cc_590 N_CK_c_573_n N_A_808_115#_c_1261_n 0.0127028f $X=4.025 $Y=1.85 $X2=5.955
+ $Y2=1.85
cc_591 N_CK_c_574_n N_A_808_115#_c_1261_n 0.00451177f $X=4.42 $Y=2.59 $X2=5.955
+ $Y2=1.85
cc_592 N_CK_c_578_n N_A_808_115#_c_1261_n 6.39375e-19 $X=4.505 $Y=2.59 $X2=5.955
+ $Y2=1.85
cc_593 N_CK_c_582_n N_A_808_115#_c_1261_n 0.0144351f $X=4.65 $Y=2.59 $X2=5.955
+ $Y2=1.85
cc_594 N_CK_c_561_n N_A_808_115#_c_1263_n 9.79344e-19 $X=4.025 $Y=1.85 $X2=3.83
+ $Y2=1.85
cc_595 N_CK_c_573_n N_A_808_115#_c_1263_n 0.00180575f $X=4.025 $Y=1.85 $X2=3.83
+ $Y2=1.85
cc_596 N_CK_c_579_n N_A_808_115#_c_1263_n 0.0128239f $X=4.36 $Y=2.59 $X2=3.83
+ $Y2=1.85
cc_597 N_A_27_115#_c_792_n N_A_428_89#_c_902_n 0.00253253f $X=3.11 $Y=1.85
+ $X2=2.335 $Y2=2.225
cc_598 N_A_27_115#_c_792_n N_A_428_89#_c_903_n 0.00296105f $X=3.11 $Y=1.85
+ $X2=2.74 $Y2=2.3
cc_599 N_A_27_115#_c_780_n N_A_428_89#_M1019_g 0.215335f $X=3.25 $Y=2.765
+ $X2=2.815 $Y2=4.585
cc_600 N_A_27_115#_c_789_n N_A_428_89#_M1019_g 0.00486364f $X=3.345 $Y=2.765
+ $X2=2.815 $Y2=4.585
cc_601 N_A_27_115#_c_778_n N_A_428_89#_c_906_n 0.0342351f $X=3.25 $Y=1.85
+ $X2=3.89 $Y2=2.3
cc_602 N_A_27_115#_c_780_n N_A_428_89#_c_906_n 0.0307748f $X=3.25 $Y=2.765
+ $X2=3.89 $Y2=2.3
cc_603 N_A_27_115#_c_789_n N_A_428_89#_c_906_n 0.0113171f $X=3.345 $Y=2.765
+ $X2=3.89 $Y2=2.3
cc_604 N_A_27_115#_c_790_n N_A_428_89#_c_906_n 8.69982e-19 $X=3.345 $Y=1.85
+ $X2=3.89 $Y2=2.3
cc_605 N_A_27_115#_c_792_n N_A_428_89#_c_906_n 0.00486036f $X=3.11 $Y=1.85
+ $X2=3.89 $Y2=2.3
cc_606 N_A_27_115#_c_827_n N_A_428_89#_c_906_n 4.12801e-19 $X=3.255 $Y=1.85
+ $X2=3.89 $Y2=2.3
cc_607 N_A_27_115#_c_779_n N_A_428_89#_M1013_g 0.211921f $X=3.53 $Y=2.765
+ $X2=3.965 $Y2=4.585
cc_608 N_A_27_115#_M1022_g N_A_808_115#_c_1256_n 0.001069f $X=3.175 $Y=1.075
+ $X2=3.685 $Y2=1.85
cc_609 N_A_27_115#_M1023_g N_A_808_115#_c_1256_n 9.36754e-19 $X=3.175 $Y=4.585
+ $X2=3.685 $Y2=1.85
cc_610 N_A_27_115#_c_776_n N_A_808_115#_c_1256_n 0.0061959f $X=3.53 $Y=1.85
+ $X2=3.685 $Y2=1.85
cc_611 N_A_27_115#_c_779_n N_A_808_115#_c_1256_n 0.00738718f $X=3.53 $Y=2.765
+ $X2=3.685 $Y2=1.85
cc_612 N_A_27_115#_M1015_g N_A_808_115#_c_1256_n 0.00502021f $X=3.605 $Y=1.075
+ $X2=3.685 $Y2=1.85
cc_613 N_A_27_115#_M1016_g N_A_808_115#_c_1256_n 0.00479454f $X=3.605 $Y=4.585
+ $X2=3.685 $Y2=1.85
cc_614 N_A_27_115#_c_789_n N_A_808_115#_c_1256_n 0.0702347f $X=3.345 $Y=2.765
+ $X2=3.685 $Y2=1.85
cc_615 N_A_27_115#_c_790_n N_A_808_115#_c_1256_n 0.0157315f $X=3.345 $Y=1.85
+ $X2=3.685 $Y2=1.85
cc_616 N_A_27_115#_c_827_n N_A_808_115#_c_1256_n 4.18442e-19 $X=3.255 $Y=1.85
+ $X2=3.685 $Y2=1.85
cc_617 N_A_27_115#_M1022_g N_A_808_115#_c_1281_n 0.00136315f $X=3.175 $Y=1.075
+ $X2=3.77 $Y2=1.43
cc_618 N_A_27_115#_M1015_g N_A_808_115#_c_1281_n 0.0099627f $X=3.605 $Y=1.075
+ $X2=3.77 $Y2=1.43
cc_619 N_A_27_115#_M1023_g N_A_808_115#_c_1325_n 9.13132e-19 $X=3.175 $Y=4.585
+ $X2=3.77 $Y2=3.185
cc_620 N_A_27_115#_M1016_g N_A_808_115#_c_1325_n 0.0096885f $X=3.605 $Y=4.585
+ $X2=3.77 $Y2=3.185
cc_621 N_A_27_115#_c_776_n N_A_808_115#_c_1263_n 0.00229064f $X=3.53 $Y=1.85
+ $X2=3.83 $Y2=1.85
cc_622 N_A_27_115#_c_790_n N_A_808_115#_c_1263_n 0.0012094f $X=3.345 $Y=1.85
+ $X2=3.83 $Y2=1.85
cc_623 N_A_27_115#_c_827_n N_A_808_115#_c_1263_n 0.0241863f $X=3.255 $Y=1.85
+ $X2=3.83 $Y2=1.85
cc_624 N_A_27_115#_c_811_n A_110_115# 0.00433061f $X=0.605 $Y=1.08 $X2=0.55
+ $Y2=0.575
cc_625 N_A_428_89#_c_909_n N_A_970_89#_M1008_g 0.0073696f $X=4.445 $Y=2.225
+ $X2=4.925 $Y2=1.075
cc_626 N_A_428_89#_c_914_n N_A_970_89#_M1008_g 0.0974852f $X=4.505 $Y=1.685
+ $X2=4.925 $Y2=1.075
cc_627 N_A_428_89#_c_917_n N_A_970_89#_M1008_g 0.0107575f $X=5.485 $Y=1.85
+ $X2=4.925 $Y2=1.075
cc_628 N_A_428_89#_c_908_n N_A_970_89#_c_1092_n 0.0073696f $X=4.37 $Y=2.3
+ $X2=4.985 $Y2=2.19
cc_629 N_A_428_89#_c_917_n N_A_970_89#_c_1092_n 0.00290516f $X=5.485 $Y=1.85
+ $X2=4.985 $Y2=2.19
cc_630 N_A_428_89#_c_926_n N_A_970_89#_c_1092_n 4.7338e-19 $X=5.845 $Y=2.25
+ $X2=4.985 $Y2=2.19
cc_631 N_A_428_89#_c_909_n N_A_970_89#_c_1103_n 0.0035305f $X=4.445 $Y=2.225
+ $X2=4.985 $Y2=2.19
cc_632 N_A_428_89#_c_917_n N_A_970_89#_c_1103_n 0.0219931f $X=5.485 $Y=1.85
+ $X2=4.985 $Y2=2.19
cc_633 N_A_428_89#_c_923_n N_A_970_89#_c_1103_n 0.00215086f $X=5.57 $Y=2.165
+ $X2=4.985 $Y2=2.19
cc_634 N_A_428_89#_c_926_n N_A_970_89#_c_1103_n 0.00359729f $X=5.845 $Y=2.25
+ $X2=4.985 $Y2=2.19
cc_635 N_A_428_89#_c_919_n N_A_970_89#_c_1104_n 0.0179204f $X=5.57 $Y=0.825
+ $X2=6.09 $Y2=0.825
cc_636 N_A_428_89#_c_919_n N_A_970_89#_c_1132_n 0.00803359f $X=5.57 $Y=0.825
+ $X2=6.175 $Y2=1.08
cc_637 N_A_428_89#_c_924_n N_A_970_89#_c_1108_n 0.0272317f $X=5.845 $Y=3.1
+ $X2=6.52 $Y2=4.815
cc_638 N_A_428_89#_c_926_n N_A_970_89#_c_1108_n 0.00224409f $X=5.845 $Y=2.25
+ $X2=6.52 $Y2=4.815
cc_639 N_A_428_89#_c_938_n N_A_970_89#_c_1108_n 0.00644034f $X=5.845 $Y=3.185
+ $X2=6.52 $Y2=4.815
cc_640 N_A_428_89#_c_926_n N_A_970_89#_c_1110_n 0.00254232f $X=5.845 $Y=2.25
+ $X2=6.52 $Y2=2.19
cc_641 N_A_428_89#_c_917_n N_A_970_89#_c_1111_n 0.00314603f $X=5.485 $Y=1.85
+ $X2=7.425 $Y2=2.19
cc_642 N_A_428_89#_c_923_n N_A_970_89#_c_1111_n 0.00659876f $X=5.57 $Y=2.165
+ $X2=7.425 $Y2=2.19
cc_643 N_A_428_89#_c_924_n N_A_970_89#_c_1111_n 0.00167455f $X=5.845 $Y=3.1
+ $X2=7.425 $Y2=2.19
cc_644 N_A_428_89#_c_926_n N_A_970_89#_c_1111_n 0.0235843f $X=5.845 $Y=2.25
+ $X2=7.425 $Y2=2.19
cc_645 N_A_428_89#_c_909_n N_A_970_89#_c_1112_n 9.14174e-19 $X=4.445 $Y=2.225
+ $X2=5.13 $Y2=2.19
cc_646 N_A_428_89#_c_917_n N_A_970_89#_c_1112_n 0.0010261f $X=5.485 $Y=1.85
+ $X2=5.13 $Y2=2.19
cc_647 N_A_428_89#_c_923_n N_A_970_89#_c_1112_n 0.00122156f $X=5.57 $Y=2.165
+ $X2=5.13 $Y2=2.19
cc_648 N_A_428_89#_c_926_n N_A_970_89#_c_1112_n 0.00122726f $X=5.845 $Y=2.25
+ $X2=5.13 $Y2=2.19
cc_649 N_A_428_89#_c_919_n N_A_808_115#_M1007_g 0.0107584f $X=5.57 $Y=0.825
+ $X2=6.305 $Y2=0.945
cc_650 N_A_428_89#_c_923_n N_A_808_115#_M1020_g 0.00280704f $X=5.57 $Y=2.165
+ $X2=6.305 $Y2=5.085
cc_651 N_A_428_89#_c_933_n N_A_808_115#_M1020_g 0.0321989f $X=5.57 $Y=3.455
+ $X2=6.305 $Y2=5.085
cc_652 N_A_428_89#_c_924_n N_A_808_115#_M1020_g 0.0115825f $X=5.845 $Y=3.1
+ $X2=6.305 $Y2=5.085
cc_653 N_A_428_89#_c_926_n N_A_808_115#_M1020_g 0.00278359f $X=5.845 $Y=2.25
+ $X2=6.305 $Y2=5.085
cc_654 N_A_428_89#_c_938_n N_A_808_115#_M1020_g 0.00343288f $X=5.845 $Y=3.185
+ $X2=6.305 $Y2=5.085
cc_655 N_A_428_89#_c_919_n N_A_808_115#_c_1255_n 0.00153999f $X=5.57 $Y=0.825
+ $X2=6.305 $Y2=1.85
cc_656 N_A_428_89#_c_923_n N_A_808_115#_c_1255_n 0.00153999f $X=5.57 $Y=2.165
+ $X2=6.305 $Y2=1.85
cc_657 N_A_428_89#_c_925_n N_A_808_115#_c_1255_n 5.35151e-19 $X=5.57 $Y=1.85
+ $X2=6.305 $Y2=1.85
cc_658 N_A_428_89#_c_906_n N_A_808_115#_c_1256_n 0.0124213f $X=3.89 $Y=2.3
+ $X2=3.685 $Y2=1.85
cc_659 N_A_428_89#_M1013_g N_A_808_115#_c_1256_n 0.0111407f $X=3.965 $Y=4.585
+ $X2=3.685 $Y2=1.85
cc_660 N_A_428_89#_c_913_n N_A_808_115#_c_1280_n 0.00174784f $X=4.505 $Y=1.85
+ $X2=4.095 $Y2=1.43
cc_661 N_A_428_89#_c_914_n N_A_808_115#_c_1280_n 0.00205316f $X=4.505 $Y=1.685
+ $X2=4.095 $Y2=1.43
cc_662 N_A_428_89#_c_917_n N_A_808_115#_c_1280_n 0.00436807f $X=5.485 $Y=1.85
+ $X2=4.095 $Y2=1.43
cc_663 N_A_428_89#_M1013_g N_A_808_115#_c_1297_n 0.0162544f $X=3.965 $Y=4.585
+ $X2=4.095 $Y2=3.185
cc_664 N_A_428_89#_c_925_n N_A_808_115#_c_1260_n 0.00755683f $X=5.57 $Y=1.85
+ $X2=6.1 $Y2=1.85
cc_665 N_A_428_89#_c_906_n N_A_808_115#_c_1261_n 0.00156696f $X=3.89 $Y=2.3
+ $X2=5.955 $Y2=1.85
cc_666 N_A_428_89#_c_908_n N_A_808_115#_c_1261_n 0.00244106f $X=4.37 $Y=2.3
+ $X2=5.955 $Y2=1.85
cc_667 N_A_428_89#_c_912_n N_A_808_115#_c_1261_n 5.19983e-19 $X=3.965 $Y=2.3
+ $X2=5.955 $Y2=1.85
cc_668 N_A_428_89#_c_913_n N_A_808_115#_c_1261_n 0.00455939f $X=4.505 $Y=1.85
+ $X2=5.955 $Y2=1.85
cc_669 N_A_428_89#_c_917_n N_A_808_115#_c_1261_n 0.0492477f $X=5.485 $Y=1.85
+ $X2=5.955 $Y2=1.85
cc_670 N_A_428_89#_c_925_n N_A_808_115#_c_1261_n 0.0106815f $X=5.57 $Y=1.85
+ $X2=5.955 $Y2=1.85
cc_671 N_A_428_89#_c_926_n N_A_808_115#_c_1261_n 0.00191587f $X=5.845 $Y=2.25
+ $X2=5.955 $Y2=1.85
cc_672 N_A_428_89#_c_906_n N_A_808_115#_c_1263_n 0.00120486f $X=3.89 $Y=2.3
+ $X2=3.83 $Y2=1.85
cc_673 N_A_428_89#_c_919_n N_A_808_115#_c_1264_n 0.00126742f $X=5.57 $Y=0.825
+ $X2=6.1 $Y2=1.85
cc_674 N_A_428_89#_c_923_n N_A_808_115#_c_1264_n 0.00126742f $X=5.57 $Y=2.165
+ $X2=6.1 $Y2=1.85
cc_675 N_A_970_89#_c_1130_n N_A_808_115#_M1007_g 0.0156439f $X=6.435 $Y=1.08
+ $X2=6.305 $Y2=0.945
cc_676 N_A_970_89#_c_1107_n N_A_808_115#_M1007_g 0.015896f $X=6.52 $Y=2.105
+ $X2=6.305 $Y2=0.945
cc_677 N_A_970_89#_c_1108_n N_A_808_115#_M1020_g 0.0331519f $X=6.52 $Y=4.815
+ $X2=6.305 $Y2=5.085
cc_678 N_A_970_89#_c_1110_n N_A_808_115#_M1020_g 0.00261985f $X=6.52 $Y=2.19
+ $X2=6.305 $Y2=5.085
cc_679 N_A_970_89#_c_1111_n N_A_808_115#_M1020_g 0.0130428f $X=7.425 $Y=2.19
+ $X2=6.305 $Y2=5.085
cc_680 N_A_970_89#_c_1132_n N_A_808_115#_c_1255_n 0.00318645f $X=6.175 $Y=1.08
+ $X2=6.305 $Y2=1.85
cc_681 N_A_970_89#_c_1111_n N_A_808_115#_c_1255_n 0.0041429f $X=7.425 $Y=2.19
+ $X2=6.305 $Y2=1.85
cc_682 N_A_970_89#_c_1130_n N_A_808_115#_c_1260_n 6.3561e-19 $X=6.435 $Y=1.08
+ $X2=6.1 $Y2=1.85
cc_683 N_A_970_89#_c_1132_n N_A_808_115#_c_1260_n 0.00206475f $X=6.175 $Y=1.08
+ $X2=6.1 $Y2=1.85
cc_684 N_A_970_89#_c_1107_n N_A_808_115#_c_1260_n 0.0115453f $X=6.52 $Y=2.105
+ $X2=6.1 $Y2=1.85
cc_685 N_A_970_89#_c_1111_n N_A_808_115#_c_1260_n 0.00483015f $X=7.425 $Y=2.19
+ $X2=6.1 $Y2=1.85
cc_686 N_A_970_89#_M1008_g N_A_808_115#_c_1261_n 0.00231271f $X=4.925 $Y=1.075
+ $X2=5.955 $Y2=1.85
cc_687 N_A_970_89#_c_1092_n N_A_808_115#_c_1261_n 0.00187603f $X=4.985 $Y=2.19
+ $X2=5.955 $Y2=1.85
cc_688 N_A_970_89#_c_1103_n N_A_808_115#_c_1261_n 0.00166223f $X=4.985 $Y=2.19
+ $X2=5.955 $Y2=1.85
cc_689 N_A_970_89#_c_1111_n N_A_808_115#_c_1261_n 0.073586f $X=7.425 $Y=2.19
+ $X2=5.955 $Y2=1.85
cc_690 N_A_970_89#_c_1112_n N_A_808_115#_c_1261_n 0.0289631f $X=5.13 $Y=2.19
+ $X2=5.955 $Y2=1.85
cc_691 N_A_970_89#_c_1107_n N_A_808_115#_c_1264_n 0.00389142f $X=6.52 $Y=2.105
+ $X2=6.1 $Y2=1.85
cc_692 N_A_970_89#_c_1111_n N_A_808_115#_c_1264_n 0.0291144f $X=7.425 $Y=2.19
+ $X2=6.1 $Y2=1.85
cc_693 N_A_970_89#_c_1094_n N_QN_M1028_g 0.0153129f $X=7.572 $Y=2.025 $X2=8.115
+ $Y2=1.075
cc_694 N_A_970_89#_c_1095_n N_QN_M1028_g 0.0391431f $X=7.66 $Y=1.65 $X2=8.115
+ $Y2=1.075
cc_695 N_A_970_89#_c_1109_n N_QN_M1028_g 4.79563e-19 $X=7.57 $Y=2.19 $X2=8.115
+ $Y2=1.075
cc_696 N_A_970_89#_c_1101_n N_QN_M1029_g 0.0102953f $X=7.66 $Y=2.855 $X2=8.115
+ $Y2=4.585
cc_697 N_A_970_89#_c_1102_n N_QN_M1029_g 0.0662174f $X=7.66 $Y=3.005 $X2=8.115
+ $Y2=4.585
cc_698 N_A_970_89#_c_1093_n N_QN_c_1383_n 0.021196f $X=7.57 $Y=2.19 $X2=8.055
+ $Y2=2.395
cc_699 N_A_970_89#_c_1109_n N_QN_c_1383_n 3.0115e-19 $X=7.57 $Y=2.19 $X2=8.055
+ $Y2=2.395
cc_700 N_A_970_89#_c_1113_n N_QN_c_1383_n 4.60229e-19 $X=7.57 $Y=2.19 $X2=8.055
+ $Y2=2.395
cc_701 N_A_970_89#_c_1095_n N_QN_c_1384_n 0.0120685f $X=7.66 $Y=1.65 $X2=7.47
+ $Y2=0.825
cc_702 N_A_970_89#_c_1100_n N_QN_c_1384_n 0.00351772f $X=7.66 $Y=1.8 $X2=7.47
+ $Y2=0.825
cc_703 N_A_970_89#_c_1101_n N_QN_c_1388_n 0.00567875f $X=7.66 $Y=2.855 $X2=7.47
+ $Y2=2.96
cc_704 N_A_970_89#_c_1102_n N_QN_c_1388_n 0.0266189f $X=7.66 $Y=3.005 $X2=7.47
+ $Y2=2.96
cc_705 N_A_970_89#_c_1094_n N_QN_c_1389_n 0.00799433f $X=7.572 $Y=2.025 $X2=7.97
+ $Y2=1.85
cc_706 N_A_970_89#_c_1100_n N_QN_c_1389_n 0.011031f $X=7.66 $Y=1.8 $X2=7.97
+ $Y2=1.85
cc_707 N_A_970_89#_c_1109_n N_QN_c_1389_n 0.0110498f $X=7.57 $Y=2.19 $X2=7.97
+ $Y2=1.85
cc_708 N_A_970_89#_c_1113_n N_QN_c_1389_n 0.00387586f $X=7.57 $Y=2.19 $X2=7.97
+ $Y2=1.85
cc_709 N_A_970_89#_c_1093_n N_QN_c_1390_n 0.00308111f $X=7.57 $Y=2.19 $X2=7.555
+ $Y2=1.85
cc_710 N_A_970_89#_c_1109_n N_QN_c_1390_n 0.0120703f $X=7.57 $Y=2.19 $X2=7.555
+ $Y2=1.85
cc_711 N_A_970_89#_c_1111_n N_QN_c_1390_n 0.0010572f $X=7.425 $Y=2.19 $X2=7.555
+ $Y2=1.85
cc_712 N_A_970_89#_c_1113_n N_QN_c_1390_n 0.00336135f $X=7.57 $Y=2.19 $X2=7.555
+ $Y2=1.85
cc_713 N_A_970_89#_c_1101_n N_QN_c_1391_n 0.016126f $X=7.66 $Y=2.855 $X2=7.97
+ $Y2=2.765
cc_714 N_A_970_89#_c_1102_n N_QN_c_1391_n 0.00248624f $X=7.66 $Y=3.005 $X2=7.97
+ $Y2=2.765
cc_715 N_A_970_89#_c_1109_n N_QN_c_1391_n 0.00426371f $X=7.57 $Y=2.19 $X2=7.97
+ $Y2=2.765
cc_716 N_A_970_89#_c_1113_n N_QN_c_1391_n 0.00253233f $X=7.57 $Y=2.19 $X2=7.97
+ $Y2=2.765
cc_717 N_A_970_89#_c_1093_n N_QN_c_1392_n 0.00265611f $X=7.57 $Y=2.19 $X2=7.555
+ $Y2=2.765
cc_718 N_A_970_89#_c_1109_n N_QN_c_1392_n 0.00471962f $X=7.57 $Y=2.19 $X2=7.555
+ $Y2=2.765
cc_719 N_A_970_89#_c_1111_n N_QN_c_1392_n 9.40773e-19 $X=7.425 $Y=2.19 $X2=7.555
+ $Y2=2.765
cc_720 N_A_970_89#_c_1113_n N_QN_c_1392_n 0.00140341f $X=7.57 $Y=2.19 $X2=7.555
+ $Y2=2.765
cc_721 N_A_970_89#_c_1093_n N_QN_c_1393_n 0.00216137f $X=7.57 $Y=2.19 $X2=8.055
+ $Y2=2.395
cc_722 N_A_970_89#_c_1094_n N_QN_c_1393_n 0.00323473f $X=7.572 $Y=2.025
+ $X2=8.055 $Y2=2.395
cc_723 N_A_970_89#_c_1101_n N_QN_c_1393_n 0.00226435f $X=7.66 $Y=2.855 $X2=8.055
+ $Y2=2.395
cc_724 N_A_970_89#_c_1109_n N_QN_c_1393_n 0.00987106f $X=7.57 $Y=2.19 $X2=8.055
+ $Y2=2.395
cc_725 N_A_970_89#_c_1113_n N_QN_c_1393_n 0.00377439f $X=7.57 $Y=2.19 $X2=8.055
+ $Y2=2.395
cc_726 N_A_970_89#_c_1102_n QN 0.00741861f $X=7.66 $Y=3.005 $X2=7.475 $Y2=2.96
cc_727 N_A_970_89#_c_1108_n QN 0.00570662f $X=6.52 $Y=4.815 $X2=7.475 $Y2=2.96
cc_728 N_A_970_89#_c_1109_n QN 0.00359685f $X=7.57 $Y=2.19 $X2=7.475 $Y2=2.96
cc_729 N_A_970_89#_c_1113_n QN 0.00842298f $X=7.57 $Y=2.19 $X2=7.475 $Y2=2.96
cc_730 N_A_970_89#_c_1102_n Q 0.0011399f $X=7.66 $Y=3.005 $X2=8.325 $Y2=3.33
cc_731 N_A_970_89#_c_1130_n A_1276_115# 0.00433061f $X=6.435 $Y=1.08 $X2=6.38
+ $Y2=0.575
cc_732 N_A_808_115#_c_1297_n A_736_617# 0.00342591f $X=4.095 $Y=3.185 $X2=3.68
+ $Y2=3.085
cc_733 N_A_808_115#_c_1325_n A_736_617# 0.00144354f $X=3.77 $Y=3.185 $X2=3.68
+ $Y2=3.085
cc_734 N_A_808_115#_c_1256_n A_736_115# 9.4749e-19 $X=3.685 $Y=1.85 $X2=3.68
+ $Y2=0.575
cc_735 N_A_808_115#_c_1280_n A_736_115# 0.00337089f $X=4.095 $Y=1.43 $X2=3.68
+ $Y2=0.575
cc_736 N_A_808_115#_c_1281_n A_736_115# 0.00148865f $X=3.77 $Y=1.43 $X2=3.68
+ $Y2=0.575
cc_737 N_QN_M1029_g N_Q_c_1468_n 0.0177846f $X=8.115 $Y=4.585 $X2=8.33 $Y2=4.475
cc_738 N_QN_M1028_g N_Q_c_1466_n 0.0383548f $X=8.115 $Y=1.075 $X2=8.445 $Y2=3.16
cc_739 N_QN_c_1389_n N_Q_c_1466_n 0.0111776f $X=7.97 $Y=1.85 $X2=8.445 $Y2=3.16
cc_740 N_QN_c_1391_n N_Q_c_1466_n 0.0111776f $X=7.97 $Y=2.765 $X2=8.445 $Y2=3.16
cc_741 N_QN_c_1393_n N_Q_c_1466_n 0.0438362f $X=8.055 $Y=2.395 $X2=8.445
+ $Y2=3.16
cc_742 N_QN_M1028_g N_Q_c_1467_n 0.00373219f $X=8.115 $Y=1.075 $X2=8.445
+ $Y2=1.515
cc_743 N_QN_M1029_g N_Q_c_1472_n 0.00613774f $X=8.115 $Y=4.585 $X2=8.33
+ $Y2=3.287
cc_744 N_QN_M1029_g Q 0.0145232f $X=8.115 $Y=4.585 $X2=8.325 $Y2=3.33
cc_745 N_QN_c_1388_n Q 0.00553023f $X=7.47 $Y=2.96 $X2=8.325 $Y2=3.33
cc_746 N_QN_c_1391_n Q 0.00245821f $X=7.97 $Y=2.765 $X2=8.325 $Y2=3.33
