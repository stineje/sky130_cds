* File: sky130_osu_sc_15T_ms__and2_l.pex.spice
* Created: Fri Nov 12 14:40:44 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__AND2_L%GND 1 17 19 26 35 38
r34 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r35 24 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r36 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r37 17 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r38 17 19 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r39 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r40 1 26 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_L%VDD 1 2 17 21 23 30 36 38 41
r25 38 41 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r26 28 36 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r27 28 30 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.235
r28 26 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r29 24 35 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r30 24 26 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r31 23 36 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r32 23 26 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r33 19 35 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r34 19 21 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.235
r35 17 26 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r36 17 35 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r37 2 30 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=3.565 $X2=1.12 $Y2=4.235
r38 1 21 300 $w=1.7e-07 $l=7.29829e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.235
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_L%A 3 7 12 15 23
r28 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=3.07
+ $X2=0.275 $Y2=3.07
r29 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.07
+ $X2=0.27 $Y2=3.07
r30 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.505
+ $X2=0.27 $Y2=3.07
r31 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.505 $X2=0.27 $Y2=2.505
r32 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.505
+ $X2=0.475 $Y2=2.505
r33 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=2.505
r34 5 7 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=4.195
r35 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=2.505
r36 1 3 771.713 $w=1.5e-07 $l=1.505e-06 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_L%B 3 7 10 14 22
r39 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.7
+ $X2=0.955 $Y2=2.7
r40 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.7 $X2=0.95
+ $Y2=2.7
r41 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.165
+ $X2=0.95 $Y2=2.7
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.165 $X2=0.95 $Y2=2.165
r43 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2.33
r44 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2
r45 7 12 956.309 $w=1.5e-07 $l=1.865e-06 $layer=POLY_cond $X=0.905 $Y=4.195
+ $X2=0.905 $Y2=2.33
r46 3 11 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=0.835 $Y=0.835
+ $X2=0.835 $Y2=2
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_L%A_27_115# 1 3 11 15 17 19 20 25 27 28 33
+ 37 39 40 41
r69 40 41 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.985
+ $X2=0.65 $Y2=4.155
r70 35 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=0.61 $Y2=1.675
r71 35 37 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=1.43 $Y2=1.675
r72 33 41 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=4.235 $X2=0.69
+ $Y2=4.155
r73 29 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.76 $X2=0.61
+ $Y2=1.675
r74 29 40 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=3.985
r75 27 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.61 $Y2=1.675
r76 27 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.345 $Y2=1.675
r77 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.345 $Y2=1.675
r78 23 25 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.825
r79 22 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.675 $X2=1.43 $Y2=1.675
r80 19 20 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.55
+ $X2=1.352 $Y2=2.7
r81 17 22 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.412 $Y2=1.675
r82 17 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=2.55
r83 15 20 766.585 $w=1.5e-07 $l=1.495e-06 $layer=POLY_cond $X=1.335 $Y=4.195
+ $X2=1.335 $Y2=2.7
r84 9 22 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.412 $Y2=1.675
r85 9 11 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.835
r86 3 33 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.565 $X2=0.69 $Y2=4.235
r87 1 25 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_L%Y 1 3 10 16 24 27 30
r33 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r34 22 24 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r35 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r36 21 24 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r37 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r38 16 19 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=4.235
r39 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r40 10 13 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.22
r41 3 19 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=3.565 $X2=1.55 $Y2=4.235
r42 1 10 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

