magic
tech sky130A
magscale 1 2
timestamp 1646342132
<< nwell >>
rect 0 1341 255 1342
rect -269 581 1317 1341
<< nmos >>
rect -180 115 -150 315
rect -94 115 -64 315
rect 96 115 126 315
rect 182 115 212 315
rect 254 115 284 315
rect 374 115 404 315
rect 446 115 476 315
rect 532 115 562 315
rect 740 115 770 315
rect 826 115 856 315
rect 1016 115 1046 315
rect 1088 115 1118 315
rect 1188 115 1218 315
<< pmos >>
rect -180 617 -150 1217
rect -108 617 -78 1217
rect 96 617 126 1217
rect 182 617 212 1217
rect 254 617 284 1217
rect 374 617 404 1217
rect 446 617 476 1217
rect 532 617 562 1217
rect 740 617 770 1217
rect 826 617 856 1217
rect 1016 617 1046 1217
rect 1102 617 1132 1217
rect 1188 617 1218 1217
<< ndiff >>
rect -233 267 -180 315
rect -233 131 -225 267
rect -191 131 -180 267
rect -233 115 -180 131
rect -150 267 -94 315
rect -150 131 -139 267
rect -105 131 -94 267
rect -150 115 -94 131
rect -64 267 -11 315
rect -64 131 -53 267
rect -19 131 -11 267
rect -64 115 -11 131
rect 43 267 96 315
rect 43 131 51 267
rect 85 131 96 267
rect 43 115 96 131
rect 126 267 182 315
rect 126 131 137 267
rect 171 131 182 267
rect 126 115 182 131
rect 212 115 254 315
rect 284 267 374 315
rect 284 131 295 267
rect 363 131 374 267
rect 284 115 374 131
rect 404 115 446 315
rect 476 267 532 315
rect 476 131 487 267
rect 521 131 532 267
rect 476 115 532 131
rect 562 267 615 315
rect 562 131 573 267
rect 607 131 615 267
rect 562 115 615 131
rect 687 267 740 315
rect 687 131 695 267
rect 729 131 740 267
rect 687 115 740 131
rect 770 267 826 315
rect 770 131 781 267
rect 815 131 826 267
rect 770 115 826 131
rect 856 267 909 315
rect 856 131 867 267
rect 901 131 909 267
rect 856 115 909 131
rect 963 267 1016 315
rect 963 131 971 267
rect 1005 131 1016 267
rect 963 115 1016 131
rect 1046 115 1088 315
rect 1118 267 1188 315
rect 1118 131 1129 267
rect 1163 131 1188 267
rect 1118 115 1188 131
rect 1218 267 1271 315
rect 1218 131 1229 267
rect 1263 131 1271 267
rect 1218 115 1271 131
<< pdiff >>
rect -233 1201 -180 1217
rect -233 657 -225 1201
rect -191 657 -180 1201
rect -233 617 -180 657
rect -150 617 -108 1217
rect -78 1201 -25 1217
rect -78 793 -67 1201
rect -33 793 -25 1201
rect -78 617 -25 793
rect 43 1201 96 1217
rect 43 725 51 1201
rect 85 725 96 1201
rect 43 617 96 725
rect 126 1201 182 1217
rect 126 725 137 1201
rect 171 725 182 1201
rect 126 617 182 725
rect 212 617 254 1217
rect 284 1201 374 1217
rect 284 657 295 1201
rect 363 657 374 1201
rect 284 617 374 657
rect 404 617 446 1217
rect 476 1201 532 1217
rect 476 657 487 1201
rect 521 657 532 1201
rect 476 617 532 657
rect 562 1201 615 1217
rect 562 657 573 1201
rect 607 657 615 1201
rect 562 617 615 657
rect 687 1201 740 1217
rect 687 657 695 1201
rect 729 657 740 1201
rect 687 617 740 657
rect 770 1201 826 1217
rect 770 657 781 1201
rect 815 657 826 1201
rect 770 617 826 657
rect 856 1201 909 1217
rect 856 657 867 1201
rect 901 657 909 1201
rect 856 617 909 657
rect 963 1201 1016 1217
rect 963 793 971 1201
rect 1005 793 1016 1201
rect 963 617 1016 793
rect 1046 1201 1102 1217
rect 1046 725 1057 1201
rect 1091 725 1102 1201
rect 1046 617 1102 725
rect 1132 1201 1188 1217
rect 1132 725 1143 1201
rect 1177 725 1188 1201
rect 1132 617 1188 725
rect 1218 1201 1271 1217
rect 1218 657 1229 1201
rect 1263 657 1271 1201
rect 1218 617 1271 657
<< ndiffc >>
rect -225 131 -191 267
rect -139 131 -105 267
rect -53 131 -19 267
rect 51 131 85 267
rect 137 131 171 267
rect 295 131 363 267
rect 487 131 521 267
rect 573 131 607 267
rect 695 131 729 267
rect 781 131 815 267
rect 867 131 901 267
rect 971 131 1005 267
rect 1129 131 1163 267
rect 1229 131 1263 267
<< pdiffc >>
rect -225 657 -191 1201
rect -67 793 -33 1201
rect 51 725 85 1201
rect 137 725 171 1201
rect 295 657 363 1201
rect 487 657 521 1201
rect 573 657 607 1201
rect 695 657 729 1201
rect 781 657 815 1201
rect 867 657 901 1201
rect 971 793 1005 1201
rect 1057 725 1091 1201
rect 1143 725 1177 1201
rect 1229 657 1263 1201
<< psubdiff >>
rect -233 27 -209 61
rect -175 27 -151 61
rect -97 27 -73 61
rect -39 27 -15 61
rect 88 27 112 61
rect 146 27 170 61
rect 224 27 248 61
rect 282 27 306 61
rect 360 27 384 61
rect 418 27 442 61
rect 496 27 520 61
rect 554 27 578 61
rect 632 27 656 61
rect 690 27 714 61
rect 768 27 792 61
rect 826 27 850 61
rect 963 27 987 61
rect 1021 27 1045 61
rect 1099 27 1123 61
rect 1157 27 1181 61
<< nsubdiff >>
rect -233 1271 -209 1305
rect -175 1271 -151 1305
rect -97 1271 -73 1305
rect -39 1271 -15 1305
rect 88 1271 112 1305
rect 146 1271 170 1305
rect 224 1271 248 1305
rect 282 1271 306 1305
rect 360 1271 384 1305
rect 418 1271 442 1305
rect 496 1271 520 1305
rect 554 1271 578 1305
rect 632 1271 656 1305
rect 690 1271 714 1305
rect 768 1271 792 1305
rect 826 1271 850 1305
rect 963 1271 987 1305
rect 1021 1271 1045 1305
rect 1099 1271 1123 1305
rect 1157 1271 1181 1305
<< psubdiffcont >>
rect -209 27 -175 61
rect -73 27 -39 61
rect 112 27 146 61
rect 248 27 282 61
rect 384 27 418 61
rect 520 27 554 61
rect 656 27 690 61
rect 792 27 826 61
rect 987 27 1021 61
rect 1123 27 1157 61
<< nsubdiffcont >>
rect -209 1271 -175 1305
rect -73 1271 -39 1305
rect 112 1271 146 1305
rect 248 1271 282 1305
rect 384 1271 418 1305
rect 520 1271 554 1305
rect 656 1271 690 1305
rect 792 1271 826 1305
rect 987 1271 1021 1305
rect 1123 1271 1157 1305
<< poly >>
rect -180 1217 -150 1243
rect -108 1217 -78 1243
rect 96 1217 126 1243
rect 182 1217 212 1243
rect 254 1217 284 1243
rect 374 1217 404 1243
rect 446 1217 476 1243
rect 532 1217 562 1243
rect 740 1217 770 1243
rect 826 1217 856 1243
rect 1016 1217 1046 1243
rect 1102 1217 1132 1243
rect 1188 1217 1218 1243
rect -180 451 -150 617
rect -108 584 -78 617
rect 96 595 126 617
rect -108 568 -35 584
rect -108 534 -79 568
rect -45 534 -35 568
rect -108 518 -35 534
rect 86 561 126 595
rect -204 435 -150 451
rect -204 401 -194 435
rect -160 401 -150 435
rect -204 385 -150 401
rect -180 315 -150 385
rect -94 315 -64 518
rect 86 403 116 561
rect 182 518 212 617
rect 254 586 284 617
rect 374 586 404 617
rect 254 570 308 586
rect 254 536 264 570
rect 298 536 308 570
rect 254 520 308 536
rect 350 570 404 586
rect 350 536 360 570
rect 394 536 404 570
rect 350 520 404 536
rect 158 502 212 518
rect 158 468 168 502
rect 202 468 212 502
rect 350 475 380 520
rect 158 452 212 468
rect 86 387 140 403
rect 86 353 96 387
rect 130 353 140 387
rect 86 337 140 353
rect 96 315 126 337
rect 182 315 212 452
rect 254 445 380 475
rect 446 477 476 617
rect 532 587 562 617
rect 740 601 770 617
rect 532 556 573 587
rect 446 461 500 477
rect 254 315 284 445
rect 446 427 456 461
rect 490 427 500 461
rect 446 411 500 427
rect 350 387 404 403
rect 350 353 360 387
rect 394 353 404 387
rect 350 337 404 353
rect 374 315 404 337
rect 446 315 476 411
rect 543 403 573 556
rect 730 571 770 601
rect 730 477 760 571
rect 826 477 856 617
rect 1016 586 1046 617
rect 963 570 1046 586
rect 963 536 973 570
rect 1007 536 1046 570
rect 963 520 1046 536
rect 705 461 760 477
rect 705 427 715 461
rect 749 427 760 461
rect 705 411 760 427
rect 802 461 856 477
rect 802 427 812 461
rect 846 427 856 461
rect 802 411 856 427
rect 543 387 601 403
rect 543 363 557 387
rect 532 353 557 363
rect 591 353 601 387
rect 532 333 601 353
rect 730 360 760 411
rect 532 315 562 333
rect 730 330 770 360
rect 740 315 770 330
rect 826 315 856 411
rect 1016 315 1046 520
rect 1102 518 1132 617
rect 1188 592 1218 617
rect 1188 562 1225 592
rect 1088 502 1153 518
rect 1088 468 1109 502
rect 1143 468 1153 502
rect 1088 452 1153 468
rect 1088 315 1118 452
rect 1195 420 1225 562
rect 1195 404 1249 420
rect 1195 384 1205 404
rect 1188 370 1205 384
rect 1239 370 1249 404
rect 1188 354 1249 370
rect 1188 315 1218 354
rect -180 89 -150 115
rect -94 89 -64 115
rect 96 89 126 115
rect 182 89 212 115
rect 254 89 284 115
rect 374 89 404 115
rect 446 89 476 115
rect 532 89 562 115
rect 740 89 770 115
rect 826 89 856 115
rect 1016 89 1046 115
rect 1088 89 1118 115
rect 1188 89 1218 115
<< polycont >>
rect -79 534 -45 568
rect -194 401 -160 435
rect 264 536 298 570
rect 360 536 394 570
rect 168 468 202 502
rect 96 353 130 387
rect 456 427 490 461
rect 360 353 394 387
rect 973 536 1007 570
rect 715 427 749 461
rect 812 427 846 461
rect 557 353 591 387
rect 1109 468 1143 502
rect 1205 370 1239 404
<< locali >>
rect -267 1311 1317 1332
rect -267 1271 -209 1311
rect -175 1271 -73 1311
rect -39 1271 112 1311
rect 146 1271 248 1311
rect 282 1271 384 1311
rect 418 1271 520 1311
rect 554 1271 656 1311
rect 690 1271 792 1311
rect 826 1271 987 1311
rect 1021 1271 1123 1311
rect 1157 1271 1317 1311
rect -225 1201 -191 1217
rect -67 1201 -33 1271
rect -67 777 -33 793
rect 51 1201 85 1217
rect 28 725 51 791
rect 28 708 85 725
rect 137 1201 171 1271
rect 137 709 171 725
rect 295 1201 363 1217
rect -225 535 -191 657
rect -147 435 -113 575
rect -79 568 -45 649
rect -79 518 -45 534
rect -210 401 -194 435
rect -160 401 -113 435
rect 28 461 62 708
rect 295 654 363 657
rect -225 267 -191 283
rect -225 61 -191 131
rect 28 296 62 427
rect 96 620 363 654
rect 487 1201 521 1271
rect 487 641 521 657
rect 573 1201 607 1217
rect 96 387 130 620
rect 360 570 394 586
rect 248 536 264 570
rect 298 536 314 570
rect 168 452 202 468
rect 280 387 314 536
rect 360 535 394 536
rect 573 535 607 657
rect 695 1201 729 1217
rect 695 570 729 649
rect 781 1201 815 1271
rect 781 641 815 657
rect 867 1201 901 1217
rect 971 1201 1005 1271
rect 971 777 1005 793
rect 1057 1201 1091 1217
rect 1041 725 1057 743
rect 1041 709 1091 725
rect 1143 1201 1177 1271
rect 1143 709 1177 725
rect 1229 1201 1263 1217
rect 901 657 914 666
rect 867 632 914 657
rect 695 536 846 570
rect 573 471 607 501
rect 440 427 456 461
rect 490 427 506 461
rect 573 437 661 471
rect 812 461 846 536
rect 557 387 591 403
rect 130 353 239 387
rect 280 353 360 387
rect 394 353 557 387
rect 96 337 130 353
rect 205 303 239 353
rect 557 337 591 353
rect 627 303 661 437
rect 699 427 715 461
rect 749 427 765 461
rect 812 387 846 427
rect -139 267 -105 279
rect -139 115 -105 131
rect -53 267 -19 283
rect 28 267 85 296
rect 28 262 51 267
rect -53 61 -19 131
rect 51 115 85 131
rect 137 267 171 283
rect 205 269 363 303
rect 137 61 171 131
rect 295 267 363 269
rect 295 115 363 131
rect 487 267 521 283
rect 487 61 521 131
rect 573 269 661 303
rect 695 353 846 387
rect 880 387 914 632
rect 973 570 1007 649
rect 973 520 1007 536
rect 1041 404 1075 709
rect 1109 502 1143 575
rect 1229 535 1263 657
rect 1109 452 1143 468
rect 1205 404 1239 420
rect 573 267 607 269
rect 573 115 607 131
rect 695 267 729 353
rect 880 319 914 353
rect 867 285 914 319
rect 971 370 1205 404
rect 695 115 729 131
rect 781 267 815 283
rect 781 61 815 131
rect 867 267 901 285
rect 867 115 901 131
rect 971 267 1005 370
rect 1205 354 1239 370
rect 971 115 1005 131
rect 1129 267 1163 283
rect 1129 61 1163 131
rect 1229 267 1263 279
rect 1229 115 1263 131
rect -267 21 -209 61
rect -175 21 -73 61
rect -39 21 112 61
rect 146 21 248 61
rect 282 21 384 61
rect 418 21 520 61
rect 554 21 656 61
rect 690 21 792 61
rect 826 21 987 61
rect 1021 21 1123 61
rect 1157 21 1317 61
rect -267 0 1317 21
<< viali >>
rect -209 1305 -175 1311
rect -209 1277 -175 1305
rect -73 1305 -39 1311
rect -73 1277 -39 1305
rect 112 1305 146 1311
rect 112 1277 146 1305
rect 248 1305 282 1311
rect 248 1277 282 1305
rect 384 1305 418 1311
rect 384 1277 418 1305
rect 520 1305 554 1311
rect 520 1277 554 1305
rect 656 1305 690 1311
rect 656 1277 690 1305
rect 792 1305 826 1311
rect 792 1277 826 1305
rect 987 1305 1021 1311
rect 987 1277 1021 1305
rect 1123 1305 1157 1311
rect 1123 1277 1157 1305
rect -79 649 -45 683
rect -225 501 -191 535
rect -147 575 -113 609
rect 28 427 62 461
rect -139 279 -105 313
rect 264 536 298 570
rect 168 502 202 536
rect 360 501 394 535
rect 695 657 729 683
rect 695 649 729 657
rect 573 501 607 535
rect 456 427 490 461
rect 557 353 591 387
rect 715 427 749 461
rect 973 649 1007 683
rect 1109 575 1143 609
rect 1229 501 1263 535
rect 880 353 914 387
rect 1229 279 1263 313
rect -209 27 -175 55
rect -209 21 -175 27
rect -73 27 -39 55
rect -73 21 -39 27
rect 112 27 146 55
rect 112 21 146 27
rect 248 27 282 55
rect 248 21 282 27
rect 384 27 418 55
rect 384 21 418 27
rect 520 27 554 55
rect 520 21 554 27
rect 656 27 690 55
rect 656 21 690 27
rect 792 27 826 55
rect 792 21 826 27
rect 987 27 1021 55
rect 987 21 1021 27
rect 1123 27 1157 55
rect 1123 21 1157 27
<< metal1 >>
rect -267 1311 1317 1332
rect -267 1277 -209 1311
rect -175 1277 -73 1311
rect -39 1277 112 1311
rect 146 1277 248 1311
rect 282 1277 384 1311
rect 418 1277 520 1311
rect 554 1277 656 1311
rect 690 1277 792 1311
rect 826 1277 987 1311
rect 1021 1277 1123 1311
rect 1157 1277 1317 1311
rect -267 1271 1317 1277
rect -91 683 -33 689
rect -112 649 -79 683
rect -45 649 -33 683
rect -91 643 -33 649
rect 682 683 740 689
rect 961 683 1019 689
rect 682 649 695 683
rect 729 649 973 683
rect 1007 649 1041 683
rect 682 643 740 649
rect 961 643 1019 649
rect -159 609 -101 615
rect 1097 609 1155 615
rect -181 575 -147 609
rect -113 575 -101 609
rect 264 576 314 609
rect -159 569 -101 575
rect 252 575 314 576
rect 1077 575 1109 609
rect 1143 575 1155 609
rect 252 570 310 575
rect -237 535 -179 541
rect 156 536 215 542
rect -142 535 168 536
rect -237 501 -225 535
rect -191 502 168 535
rect 202 502 215 536
rect 252 536 264 570
rect 298 536 310 570
rect 1097 569 1155 575
rect 252 530 310 536
rect 348 535 406 541
rect 561 535 619 541
rect -191 501 215 502
rect -237 495 -179 501
rect -139 319 -105 501
rect 156 496 215 501
rect 348 501 360 535
rect 394 501 573 535
rect 607 501 619 535
rect 348 495 406 501
rect 561 495 619 501
rect 1217 535 1275 541
rect 1217 501 1229 535
rect 1263 501 1275 535
rect 1217 495 1275 501
rect 15 461 74 467
rect 15 427 28 461
rect 62 454 74 461
rect 444 461 503 467
rect 444 454 456 461
rect 62 427 456 454
rect 490 458 503 461
rect 703 461 761 467
rect 703 458 715 461
rect 490 430 715 458
rect 490 427 503 430
rect 15 426 503 427
rect 15 421 74 426
rect 444 421 503 426
rect 703 427 715 430
rect 749 427 761 461
rect 703 421 761 427
rect 543 387 603 393
rect 521 353 557 387
rect 591 353 603 387
rect 543 347 603 353
rect 867 387 927 396
rect 867 353 880 387
rect 914 353 942 387
rect 867 352 942 353
rect 867 344 927 352
rect 1229 319 1263 495
rect -151 313 -93 319
rect -151 279 -139 313
rect -105 279 -93 313
rect -151 273 -93 279
rect 1217 313 1275 319
rect 1217 279 1229 313
rect 1263 279 1275 313
rect 1217 273 1275 279
rect -267 55 1317 61
rect -267 21 -209 55
rect -175 21 -73 55
rect -39 21 112 55
rect 146 21 248 55
rect 282 21 384 55
rect 418 21 520 55
rect 554 21 656 55
rect 690 21 792 55
rect 826 21 987 55
rect 1021 21 1123 55
rect 1157 21 1317 55
rect -267 0 1317 21
<< labels >>
rlabel metal1 -131 592 -131 592 1 SE
port 1 n
rlabel metal1 -62 667 -62 667 1 E
port 2 n
rlabel metal1 574 370 574 370 1 CK
port 3 n
rlabel metal1 1245 443 1245 443 1 ECK
port 4 n
rlabel metal1 -192 44 -192 44 1 gnd
rlabel metal1 -56 44 -56 44 1 gnd
rlabel metal1 129 44 129 44 1 gnd
rlabel metal1 264 42 264 42 1 gnd
rlabel metal1 401 39 401 39 1 gnd
rlabel metal1 537 39 537 39 1 gnd
rlabel metal1 673 40 673 40 1 gnd
rlabel metal1 809 40 809 40 1 gnd
rlabel metal1 1004 40 1004 40 1 gnd
rlabel metal1 1140 40 1140 40 1 gnd
rlabel metal1 -192 1290 -192 1290 1 vdd
rlabel metal1 -55 1291 -55 1291 1 vdd
rlabel metal1 129 1292 129 1292 1 vdd
rlabel metal1 265 1292 265 1292 1 vdd
rlabel metal1 401 1292 401 1292 1 vdd
rlabel metal1 538 1294 538 1294 1 vdd
rlabel metal1 673 1293 673 1293 1 vdd
rlabel metal1 809 1292 809 1292 1 vdd
rlabel metal1 1005 1293 1005 1293 1 vdd
rlabel metal1 1141 1293 1141 1293 1 vdd
rlabel metal1 895 366 895 370 1 Q
port 5 n
rlabel metal1 1126 593 1126 593 1 CKa
port 6 n
<< end >>
