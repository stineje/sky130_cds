* File: sky130_osu_sc_18T_ms__inv_3.pex.spice
* Created: Thu Oct 29 17:29:56 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%GND 1 2 15 19 23 31 32 34 37
r45 34 37 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r46 31 32 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r47 21 32 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r48 21 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.825
r49 17 19 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r50 15 31 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r51 15 27 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r52 15 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.17
+ $X2=1.02 $Y2=0.17
r53 15 17 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r54 15 27 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r55 2 23 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r56 1 19 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%VDD 1 2 13 17 23 32 33 35 38
r33 38 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=6.49
+ $X2=1.02 $Y2=6.49
r34 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.02 $Y2=6.507
r35 32 42 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r36 32 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r37 29 42 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r38 29 31 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r39 23 26 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r40 21 33 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r41 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r42 17 20 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r43 15 31 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r44 15 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r45 13 42 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r46 13 31 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r47 2 26 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r48 2 23 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r49 1 20 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r50 1 17 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 32 33 34 35 37 38 42 45 47
c96 38 0 1.5442e-19 $X=0.535 $Y=2.305
c97 28 0 1.33323e-19 $X=1.335 $Y=2.96
c98 25 0 1.33323e-19 $X=1.335 $Y=1.7
c99 18 0 1.33323e-19 $X=0.905 $Y=2.96
c100 15 0 1.33323e-19 $X=0.905 $Y=1.7
r101 42 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r102 40 45 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=2.39
+ $X2=0.32 $Y2=3.33
r103 38 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.47
r104 38 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=2.305
+ $X2=0.535 $Y2=2.14
r105 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=2.305 $X2=0.535 $Y2=2.305
r106 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.405 $Y=2.305
+ $X2=0.32 $Y2=2.39
r107 35 37 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=2.305
+ $X2=0.535 $Y2=2.305
r108 28 30 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r109 25 27 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.335 $Y=1.7
+ $X2=1.335 $Y2=1.075
r110 24 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.885
+ $X2=0.905 $Y2=2.885
r111 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=1.335 $Y2=2.96
r112 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.885
+ $X2=0.98 $Y2=2.885
r113 22 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.775
+ $X2=0.905 $Y2=1.775
r114 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=1.335 $Y2=1.7
r115 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.775
+ $X2=0.98 $Y2=1.775
r116 18 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=2.885
r117 18 20 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.905 $Y=2.96
+ $X2=0.905 $Y2=4.585
r118 15 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.775
r119 15 17 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.905 $Y=1.7
+ $X2=0.905 $Y2=1.075
r120 14 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.885
+ $X2=0.475 $Y2=2.885
r121 13 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.905 $Y2=2.885
r122 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.885
+ $X2=0.55 $Y2=2.885
r123 12 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.775
+ $X2=0.475 $Y2=1.775
r124 11 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.905 $Y2=1.775
r125 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.775
+ $X2=0.55 $Y2=1.775
r126 8 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=2.885
r127 8 10 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=0.475 $Y=2.96
+ $X2=0.475 $Y2=4.585
r128 7 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.885
r129 7 48 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.81
+ $X2=0.475 $Y2=2.47
r130 4 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=1.775
r131 4 47 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.85
+ $X2=0.475 $Y2=2.14
r132 1 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.775
r133 1 3 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_MS__INV_3%Y 1 2 3 4 13 14 16 18 20 22 23 29 35 37
+ 49
c74 37 0 1.5442e-19 $X=0.69 $Y=0.825
c75 23 0 1.33323e-19 $X=1.55 $Y=2.845
c76 22 0 1.33323e-19 $X=1.55 $Y=1.595
c77 14 0 1.33323e-19 $X=0.69 $Y=2.845
c78 13 0 1.33323e-19 $X=0.69 $Y=1.595
r79 56 58 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r80 44 46 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r81 35 56 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=3.455
r82 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.96
+ $X2=1.55 $Y2=2.96
r83 32 49 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=0.825
r84 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r85 29 44 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=3.455
r86 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.96
+ $X2=0.69 $Y2=2.96
r87 26 37 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=0.825
r88 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.48
r89 23 34 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.845
+ $X2=1.55 $Y2=2.96
r90 22 31 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r91 22 23 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.845
r92 21 28 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.96
+ $X2=0.69 $Y2=2.96
r93 20 34 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=1.55 $Y2=2.96
r94 20 21 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.96
+ $X2=0.835 $Y2=2.96
r95 19 25 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.48
+ $X2=0.69 $Y2=1.48
r96 18 31 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=1.55 $Y2=1.48
r97 18 19 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1.48
+ $X2=0.835 $Y2=1.48
r98 14 28 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.96
r99 14 16 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.845
+ $X2=0.69 $Y2=2.2
r100 13 25 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.48
r101 13 16 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=2.2
r102 4 58 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r103 4 56 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r104 3 46 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r105 3 44 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r106 2 49 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r107 1 37 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

