* File: sky130_osu_sc_18T_hs__ncgate_1.pxi.spice
* Created: Thu Mar 10 17:10:01 2022
* 
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%GND N_GND_M1014_s N_GND_M1024_d
+ N_GND_M1003_d N_GND_M1005_d N_GND_M1022_d N_GND_M1018_s N_GND_M1021_d
+ N_GND_M1014_b N_GND_c_2_p N_GND_c_3_p N_GND_c_14_p N_GND_c_22_p N_GND_c_19_p
+ N_GND_c_33_p N_GND_c_61_p N_GND_c_64_p N_GND_c_109_p N_GND_c_130_p
+ N_GND_c_131_p N_GND_c_79_p N_GND_c_80_p N_GND_c_156_p GND GND GND GND GND GND
+ GND GND GND GND N_GND_c_4_p PM_SKY130_OSU_SC_18T_HS__NCGATE_1%GND
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%VDD N_VDD_M1017_d N_VDD_M1001_d
+ N_VDD_M1004_d N_VDD_M1019_d N_VDD_M1020_d N_VDD_M1011_b N_VDD_c_183_p
+ N_VDD_c_189_p N_VDD_c_199_p N_VDD_c_200_p N_VDD_c_206_p N_VDD_c_229_p
+ N_VDD_c_220_p N_VDD_c_249_p N_VDD_c_233_p N_VDD_c_234_p N_VDD_c_275_p VDD VDD
+ VDD N_VDD_c_184_p PM_SKY130_OSU_SC_18T_HS__NCGATE_1%VDD
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%SE N_SE_M1014_g N_SE_M1011_g N_SE_c_295_n
+ N_SE_c_297_n N_SE_c_299_n SE N_SE_X27_noxref_CONDUCTOR
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%SE
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%E N_E_M1017_g N_E_M1024_g N_E_c_344_n
+ N_E_c_345_n E N_E_X28_noxref_CONDUCTOR PM_SKY130_OSU_SC_18T_HS__NCGATE_1%E
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_86_332# N_A_86_332#_M1025_d
+ N_A_86_332#_M1023_d N_A_86_332#_M1003_g N_A_86_332#_M1001_g
+ N_A_86_332#_c_387_n N_A_86_332#_c_389_n N_A_86_332#_c_394_n
+ N_A_86_332#_c_395_n N_A_86_332#_c_396_n N_A_86_332#_c_397_n
+ N_A_86_332#_c_398_n N_A_86_332#_c_410_n N_A_86_332#_c_458_p
+ N_A_86_332#_c_400_n N_A_86_332#_c_441_p N_A_86_332#_c_423_p
+ N_A_86_332#_c_401_n N_A_86_332#_c_412_n
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_86_332#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_N233_612# N_A_N233_612#_M1014_d
+ N_A_N233_612#_M1011_s N_A_N233_612#_M1002_g N_A_N233_612#_M1000_g
+ N_A_N233_612#_c_475_n N_A_N233_612#_c_476_n N_A_N233_612#_c_477_n
+ N_A_N233_612#_c_480_n N_A_N233_612#_c_481_n N_A_N233_612#_c_482_n
+ N_A_N233_612#_c_483_n N_A_N233_612#_c_484_n N_A_N233_612#_c_485_n
+ N_A_N233_612#_c_488_n PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_N233_612#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_254_515# N_A_254_515#_M1007_d
+ N_A_254_515#_M1006_d N_A_254_515#_M1023_g N_A_254_515#_M1015_g
+ N_A_254_515#_c_574_n N_A_254_515#_c_575_n N_A_254_515#_c_576_n
+ N_A_254_515#_c_579_n N_A_254_515#_c_580_n N_A_254_515#_c_582_n
+ N_A_254_515#_c_583_n N_A_254_515#_c_586_n N_A_254_515#_c_595_n
+ N_A_254_515#_c_587_n N_A_254_515#_c_588_n N_A_254_515#_c_589_n
+ N_A_254_515#_c_590_n N_A_254_515#_c_599_n
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_254_515#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%CK N_CK_M1025_g N_CK_c_703_n N_CK_c_704_n
+ N_CK_M1012_g N_CK_M1007_g N_CK_c_705_n N_CK_M1006_g N_CK_c_706_n N_CK_M1021_g
+ N_CK_M1020_g N_CK_c_712_n N_CK_c_713_n N_CK_c_714_n N_CK_c_718_n N_CK_c_719_n
+ N_CK_c_720_n N_CK_c_721_n N_CK_c_722_n N_CK_c_744_n N_CK_c_723_n N_CK_c_724_n
+ N_CK_c_725_n N_CK_c_726_n CK N_CK_c_727_n PM_SKY130_OSU_SC_18T_HS__NCGATE_1%CK
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_43_110# N_A_43_110#_M1003_s
+ N_A_43_110#_M1001_s N_A_43_110#_M1005_g N_A_43_110#_M1004_g
+ N_A_43_110#_M1022_g N_A_43_110#_M1019_g N_A_43_110#_c_897_n
+ N_A_43_110#_c_898_n N_A_43_110#_c_899_n N_A_43_110#_c_900_n
+ N_A_43_110#_c_904_n N_A_43_110#_c_905_n N_A_43_110#_c_906_n
+ N_A_43_110#_c_907_n N_A_43_110#_c_908_n N_A_43_110#_c_930_n
+ N_A_43_110#_c_912_n N_A_43_110#_c_913_n N_A_43_110#_c_914_n
+ N_A_43_110#_c_934_n N_A_43_110#_c_916_n N_A_43_110#_c_917_n
+ N_A_43_110#_c_918_n N_A_43_110#_c_919_n N_A_43_110#_c_920_n
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_43_110#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_687_110# N_A_687_110#_M1022_s
+ N_A_687_110#_M1019_s N_A_687_110#_M1009_g N_A_687_110#_M1008_g
+ N_A_687_110#_M1018_g N_A_687_110#_M1016_g N_A_687_110#_c_1076_n
+ N_A_687_110#_c_1077_n N_A_687_110#_c_1078_n N_A_687_110#_c_1081_n
+ N_A_687_110#_c_1082_n N_A_687_110#_c_1084_n N_A_687_110#_c_1085_n
+ N_A_687_110#_c_1086_n N_A_687_110#_c_1087_n N_A_687_110#_c_1088_n
+ N_A_687_110#_c_1089_n N_A_687_110#_c_1090_n
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_687_110#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_963_612# N_A_963_612#_M1018_d
+ N_A_963_612#_M1016_s N_A_963_612#_M1013_g N_A_963_612#_M1010_g
+ N_A_963_612#_c_1191_n N_A_963_612#_c_1192_n N_A_963_612#_c_1193_n
+ N_A_963_612#_c_1205_n N_A_963_612#_c_1218_n N_A_963_612#_c_1235_n
+ N_A_963_612#_c_1194_n N_A_963_612#_c_1195_n N_A_963_612#_c_1198_n
+ N_A_963_612#_c_1200_n PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_963_612#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_856_110# N_A_856_110#_M1009_d
+ N_A_856_110#_M1008_d N_A_856_110#_c_1269_n N_A_856_110#_c_1275_n
+ N_A_856_110#_c_1277_n N_A_856_110#_c_1273_n N_A_856_110#_c_1274_n
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%A_856_110#
x_PM_SKY130_OSU_SC_18T_HS__NCGATE_1%ECK N_ECK_M1013_d N_ECK_M1010_d
+ N_ECK_c_1304_n N_ECK_c_1307_n N_ECK_c_1308_n N_ECK_c_1309_n ECK
+ PM_SKY130_OSU_SC_18T_HS__NCGATE_1%ECK
cc_1 N_GND_M1014_b N_SE_M1014_g 0.0397546f $X=-1.345 $Y=-0.025 $X2=-0.825
+ $Y2=1.05
cc_2 N_GND_c_2_p N_SE_M1014_g 0.00713292f $X=-1.039 $Y=0.8 $X2=-0.825 $Y2=1.05
cc_3 N_GND_c_3_p N_SE_M1014_g 0.00606474f $X=-0.265 $Y=0.127 $X2=-0.825 $Y2=1.05
cc_4 N_GND_c_4_p N_SE_M1014_g 0.00468827f $X=5.7 $Y=0.165 $X2=-0.825 $Y2=1.05
cc_5 N_GND_M1014_b N_SE_M1011_g 0.0432223f $X=-1.345 $Y=-0.025 $X2=-0.825
+ $Y2=4.56
cc_6 N_GND_M1014_b N_SE_c_295_n 0.0362021f $X=-1.345 $Y=-0.025 $X2=-0.884
+ $Y2=2.065
cc_7 N_GND_c_2_p N_SE_c_295_n 0.00122211f $X=-1.039 $Y=0.8 $X2=-0.884 $Y2=2.065
cc_8 N_GND_M1014_b N_SE_c_297_n 0.0115466f $X=-1.345 $Y=-0.025 $X2=-0.735
+ $Y2=2.065
cc_9 N_GND_c_2_p N_SE_c_297_n 0.00289632f $X=-1.039 $Y=0.8 $X2=-0.735 $Y2=2.065
cc_10 N_GND_M1014_b N_SE_c_299_n 0.0148611f $X=-1.345 $Y=-0.025 $X2=-0.649
+ $Y2=2.935
cc_11 N_GND_M1014_b N_SE_X27_noxref_CONDUCTOR 5.75357e-19 $X=-1.345 $Y=-0.025
+ $X2=-0.649 $Y2=2.935
cc_12 N_GND_M1014_b N_E_M1024_g 0.0744003f $X=-1.345 $Y=-0.025 $X2=-0.395
+ $Y2=1.05
cc_13 N_GND_c_3_p N_E_M1024_g 0.00606474f $X=-0.265 $Y=0.127 $X2=-0.395 $Y2=1.05
cc_14 N_GND_c_14_p N_E_M1024_g 0.00713292f $X=-0.179 $Y=0.8 $X2=-0.395 $Y2=1.05
cc_15 N_GND_c_4_p N_E_M1024_g 0.00468827f $X=5.7 $Y=0.165 $X2=-0.395 $Y2=1.05
cc_16 N_GND_M1014_b N_E_c_344_n 0.032073f $X=-1.345 $Y=-0.025 $X2=-0.309
+ $Y2=2.73
cc_17 N_GND_M1014_b N_E_c_345_n 0.00121702f $X=-1.345 $Y=-0.025 $X2=-0.309
+ $Y2=2.73
cc_18 N_GND_M1014_b N_A_86_332#_c_387_n 0.030793f $X=-1.345 $Y=-0.025 $X2=0.565
+ $Y2=1.825
cc_19 N_GND_c_19_p N_A_86_332#_c_387_n 3.17551e-19 $X=0.77 $Y=0.8 $X2=0.565
+ $Y2=1.825
cc_20 N_GND_M1014_b N_A_86_332#_c_389_n 0.0184872f $X=-1.345 $Y=-0.025 $X2=0.565
+ $Y2=1.66
cc_21 N_GND_c_14_p N_A_86_332#_c_389_n 0.00458302f $X=-0.179 $Y=0.8 $X2=0.565
+ $Y2=1.66
cc_22 N_GND_c_22_p N_A_86_332#_c_389_n 0.00606474f $X=0.685 $Y=0.127 $X2=0.565
+ $Y2=1.66
cc_23 N_GND_c_19_p N_A_86_332#_c_389_n 0.00354579f $X=0.77 $Y=0.8 $X2=0.565
+ $Y2=1.66
cc_24 N_GND_c_4_p N_A_86_332#_c_389_n 0.00468827f $X=5.7 $Y=0.165 $X2=0.565
+ $Y2=1.66
cc_25 N_GND_M1014_b N_A_86_332#_c_394_n 0.0436632f $X=-1.345 $Y=-0.025 $X2=0.53
+ $Y2=2.78
cc_26 N_GND_M1014_b N_A_86_332#_c_395_n 0.00768983f $X=-1.345 $Y=-0.025 $X2=0.53
+ $Y2=2.95
cc_27 N_GND_M1014_b N_A_86_332#_c_396_n 8.14549e-19 $X=-1.345 $Y=-0.025
+ $X2=0.565 $Y2=1.91
cc_28 N_GND_M1014_b N_A_86_332#_c_397_n 0.00712579f $X=-1.345 $Y=-0.025
+ $X2=0.565 $Y2=3.075
cc_29 N_GND_M1014_b N_A_86_332#_c_398_n 0.00828074f $X=-1.345 $Y=-0.025
+ $X2=1.025 $Y2=1.825
cc_30 N_GND_c_19_p N_A_86_332#_c_398_n 0.00816426f $X=0.77 $Y=0.8 $X2=1.025
+ $Y2=1.825
cc_31 N_GND_M1014_b N_A_86_332#_c_400_n 0.00172671f $X=-1.345 $Y=-0.025 $X2=1.11
+ $Y2=1.74
cc_32 N_GND_M1014_b N_A_86_332#_c_401_n 0.00313975f $X=-1.345 $Y=-0.025
+ $X2=1.645 $Y2=0.8
cc_33 N_GND_c_33_p N_A_86_332#_c_401_n 0.0151591f $X=2.435 $Y=0.127 $X2=1.645
+ $Y2=0.8
cc_34 N_GND_c_4_p N_A_86_332#_c_401_n 0.00958198f $X=5.7 $Y=0.165 $X2=1.645
+ $Y2=0.8
cc_35 N_GND_M1014_b N_A_N233_612#_M1002_g 0.040459f $X=-1.345 $Y=-0.025
+ $X2=0.985 $Y2=1.05
cc_36 N_GND_c_19_p N_A_N233_612#_M1002_g 0.00354579f $X=0.77 $Y=0.8 $X2=0.985
+ $Y2=1.05
cc_37 N_GND_c_33_p N_A_N233_612#_M1002_g 0.00606474f $X=2.435 $Y=0.127 $X2=0.985
+ $Y2=1.05
cc_38 N_GND_c_4_p N_A_N233_612#_M1002_g 0.00468827f $X=5.7 $Y=0.165 $X2=0.985
+ $Y2=1.05
cc_39 N_GND_M1014_b N_A_N233_612#_M1000_g 0.0152798f $X=-1.345 $Y=-0.025
+ $X2=0.985 $Y2=4.56
cc_40 N_GND_M1014_b N_A_N233_612#_c_475_n 0.0294636f $X=-1.345 $Y=-0.025
+ $X2=0.925 $Y2=2.4
cc_41 N_GND_M1014_b N_A_N233_612#_c_476_n 0.0154673f $X=-1.345 $Y=-0.025
+ $X2=-1.039 $Y2=2.565
cc_42 N_GND_M1014_b N_A_N233_612#_c_477_n 0.00155118f $X=-1.345 $Y=-0.025
+ $X2=-0.609 $Y2=0.8
cc_43 N_GND_c_3_p N_A_N233_612#_c_477_n 0.0075556f $X=-0.265 $Y=0.127 $X2=-0.609
+ $Y2=0.8
cc_44 N_GND_c_4_p N_A_N233_612#_c_477_n 0.00475776f $X=5.7 $Y=0.165 $X2=-0.609
+ $Y2=0.8
cc_45 N_GND_M1014_b N_A_N233_612#_c_480_n 0.00123417f $X=-1.345 $Y=-0.025
+ $X2=0.925 $Y2=2.4
cc_46 N_GND_M1014_b N_A_N233_612#_c_481_n 2.54997e-19 $X=-1.345 $Y=-0.025
+ $X2=-0.695 $Y2=2.565
cc_47 N_GND_M1014_b N_A_N233_612#_c_482_n 0.019675f $X=-1.345 $Y=-0.025
+ $X2=-0.895 $Y2=2.565
cc_48 N_GND_M1014_b N_A_N233_612#_c_483_n 0.0195542f $X=-1.345 $Y=-0.025
+ $X2=-0.61 $Y2=2.48
cc_49 N_GND_M1014_b N_A_N233_612#_c_484_n 0.0416807f $X=-1.345 $Y=-0.025
+ $X2=0.78 $Y2=2.565
cc_50 N_GND_M1014_b N_A_N233_612#_c_485_n 0.00257875f $X=-1.345 $Y=-0.025
+ $X2=-0.609 $Y2=1.455
cc_51 N_GND_c_2_p N_A_N233_612#_c_485_n 0.00125659f $X=-1.039 $Y=0.8 $X2=-0.609
+ $Y2=1.455
cc_52 N_GND_c_14_p N_A_N233_612#_c_485_n 0.00125659f $X=-0.179 $Y=0.8 $X2=-0.609
+ $Y2=1.455
cc_53 N_GND_M1014_b N_A_N233_612#_c_488_n 2.07344e-19 $X=-1.345 $Y=-0.025
+ $X2=-0.61 $Y2=2.565
cc_54 N_GND_M1014_b N_A_254_515#_c_574_n 0.019996f $X=-1.345 $Y=-0.025 $X2=1.405
+ $Y2=2.74
cc_55 N_GND_M1014_b N_A_254_515#_c_575_n 0.0303093f $X=-1.345 $Y=-0.025
+ $X2=1.885 $Y2=1.825
cc_56 N_GND_M1014_b N_A_254_515#_c_576_n 0.0175443f $X=-1.345 $Y=-0.025
+ $X2=1.885 $Y2=1.66
cc_57 N_GND_c_33_p N_A_254_515#_c_576_n 0.00606474f $X=2.435 $Y=0.127 $X2=1.885
+ $Y2=1.66
cc_58 N_GND_c_4_p N_A_254_515#_c_576_n 0.00468827f $X=5.7 $Y=0.165 $X2=1.885
+ $Y2=1.66
cc_59 N_GND_M1014_b N_A_254_515#_c_579_n 0.0071877f $X=-1.345 $Y=-0.025
+ $X2=1.485 $Y2=2.655
cc_60 N_GND_M1014_b N_A_254_515#_c_580_n 0.020865f $X=-1.345 $Y=-0.025 $X2=2.865
+ $Y2=1.825
cc_61 N_GND_c_61_p N_A_254_515#_c_580_n 0.00821845f $X=2.52 $Y=0.8 $X2=2.865
+ $Y2=1.825
cc_62 N_GND_M1014_b N_A_254_515#_c_582_n 0.00162414f $X=-1.345 $Y=-0.025
+ $X2=1.57 $Y2=1.825
cc_63 N_GND_M1014_b N_A_254_515#_c_583_n 0.00538063f $X=-1.345 $Y=-0.025
+ $X2=2.95 $Y2=0.8
cc_64 N_GND_c_64_p N_A_254_515#_c_583_n 0.00754714f $X=3.905 $Y=0.127 $X2=2.95
+ $Y2=0.8
cc_65 N_GND_c_4_p N_A_254_515#_c_583_n 0.00476261f $X=5.7 $Y=0.165 $X2=2.95
+ $Y2=0.8
cc_66 N_GND_M1014_b N_A_254_515#_c_586_n 0.0045692f $X=-1.345 $Y=-0.025 $X2=2.95
+ $Y2=2.11
cc_67 N_GND_M1014_b N_A_254_515#_c_587_n 0.0132581f $X=-1.345 $Y=-0.025 $X2=3.22
+ $Y2=3.075
cc_68 N_GND_M1014_b N_A_254_515#_c_588_n 0.00375832f $X=-1.345 $Y=-0.025
+ $X2=1.485 $Y2=2.74
cc_69 N_GND_M1014_b N_A_254_515#_c_589_n 0.00185575f $X=-1.345 $Y=-0.025
+ $X2=2.95 $Y2=1.825
cc_70 N_GND_M1014_b N_A_254_515#_c_590_n 0.0156879f $X=-1.345 $Y=-0.025 $X2=3.22
+ $Y2=2.195
cc_71 N_GND_M1014_b N_CK_M1025_g 0.0458897f $X=-1.345 $Y=-0.025 $X2=1.345
+ $Y2=1.05
cc_72 N_GND_c_33_p N_CK_M1025_g 0.00606474f $X=2.435 $Y=0.127 $X2=1.345 $Y2=1.05
cc_73 N_GND_c_4_p N_CK_M1025_g 0.00468827f $X=5.7 $Y=0.165 $X2=1.345 $Y2=1.05
cc_74 N_GND_M1014_b N_CK_c_703_n 0.032998f $X=-1.345 $Y=-0.025 $X2=1.75
+ $Y2=2.275
cc_75 N_GND_M1014_b N_CK_c_704_n 0.00717301f $X=-1.345 $Y=-0.025 $X2=1.42
+ $Y2=2.275
cc_76 N_GND_M1014_b N_CK_c_705_n 0.0313734f $X=-1.345 $Y=-0.025 $X2=2.735
+ $Y2=2.905
cc_77 N_GND_M1014_b N_CK_c_706_n 0.0458999f $X=-1.345 $Y=-0.025 $X2=2.79
+ $Y2=2.575
cc_78 N_GND_M1014_b N_CK_M1021_g 0.0440597f $X=-1.345 $Y=-0.025 $X2=5.585
+ $Y2=1.05
cc_79 N_GND_c_79_p N_CK_M1021_g 0.00606474f $X=5.715 $Y=0.127 $X2=5.585 $Y2=1.05
cc_80 N_GND_c_80_p N_CK_M1021_g 0.00354579f $X=5.8 $Y=0.8 $X2=5.585 $Y2=1.05
cc_81 N_GND_c_4_p N_CK_M1021_g 0.00468827f $X=5.7 $Y=0.165 $X2=5.585 $Y2=1.05
cc_82 N_GND_M1014_b N_CK_M1020_g 0.0166256f $X=-1.345 $Y=-0.025 $X2=5.585
+ $Y2=4.56
cc_83 N_GND_M1014_b N_CK_c_712_n 0.0203203f $X=-1.345 $Y=-0.025 $X2=1.885
+ $Y2=2.74
cc_84 N_GND_M1014_b N_CK_c_713_n 0.0135787f $X=-1.345 $Y=-0.025 $X2=1.885
+ $Y2=2.575
cc_85 N_GND_M1014_b N_CK_c_714_n 0.0195174f $X=-1.345 $Y=-0.025 $X2=2.762
+ $Y2=1.64
cc_86 N_GND_c_61_p N_CK_c_714_n 0.00354579f $X=2.52 $Y=0.8 $X2=2.762 $Y2=1.64
cc_87 N_GND_c_64_p N_CK_c_714_n 0.00606474f $X=3.905 $Y=0.127 $X2=2.762 $Y2=1.64
cc_88 N_GND_c_4_p N_CK_c_714_n 0.00468827f $X=5.7 $Y=0.165 $X2=2.762 $Y2=1.64
cc_89 N_GND_M1014_b N_CK_c_718_n 0.0140659f $X=-1.345 $Y=-0.025 $X2=2.762
+ $Y2=1.79
cc_90 N_GND_M1014_b N_CK_c_719_n 0.0271998f $X=-1.345 $Y=-0.025 $X2=5.63
+ $Y2=2.36
cc_91 N_GND_M1014_b N_CK_c_720_n 0.00180771f $X=-1.345 $Y=-0.025 $X2=1.885
+ $Y2=2.565
cc_92 N_GND_M1014_b N_CK_c_721_n 7.11312e-19 $X=-1.345 $Y=-0.025 $X2=2.88
+ $Y2=2.565
cc_93 N_GND_M1014_b N_CK_c_722_n 0.00338116f $X=-1.345 $Y=-0.025 $X2=5.63
+ $Y2=2.36
cc_94 N_GND_M1014_b N_CK_c_723_n 0.0171043f $X=-1.345 $Y=-0.025 $X2=2.735
+ $Y2=2.565
cc_95 N_GND_M1014_b N_CK_c_724_n 0.00388969f $X=-1.345 $Y=-0.025 $X2=2.03
+ $Y2=2.565
cc_96 N_GND_M1014_b N_CK_c_725_n 0.0408641f $X=-1.345 $Y=-0.025 $X2=5.485
+ $Y2=2.565
cc_97 N_GND_M1014_b N_CK_c_726_n 0.0011022f $X=-1.345 $Y=-0.025 $X2=3.025
+ $Y2=2.565
cc_98 N_GND_M1014_b N_CK_c_727_n 0.00272833f $X=-1.345 $Y=-0.025 $X2=5.63
+ $Y2=2.565
cc_99 N_GND_M1014_b N_A_43_110#_M1005_g 0.0341436f $X=-1.345 $Y=-0.025 $X2=2.305
+ $Y2=1.05
cc_100 N_GND_c_33_p N_A_43_110#_M1005_g 0.00606474f $X=2.435 $Y=0.127 $X2=2.305
+ $Y2=1.05
cc_101 N_GND_c_61_p N_A_43_110#_M1005_g 0.00354579f $X=2.52 $Y=0.8 $X2=2.305
+ $Y2=1.05
cc_102 N_GND_c_4_p N_A_43_110#_M1005_g 0.00468827f $X=5.7 $Y=0.165 $X2=2.305
+ $Y2=1.05
cc_103 N_GND_M1014_b N_A_43_110#_M1004_g 0.0266205f $X=-1.345 $Y=-0.025
+ $X2=2.305 $Y2=4.56
cc_104 N_GND_M1014_b N_A_43_110#_c_897_n 0.0287113f $X=-1.345 $Y=-0.025
+ $X2=2.365 $Y2=2.195
cc_105 N_GND_M1014_b N_A_43_110#_c_898_n 0.0282897f $X=-1.345 $Y=-0.025 $X2=3.66
+ $Y2=2.195
cc_106 N_GND_M1014_b N_A_43_110#_c_899_n 0.0159661f $X=-1.345 $Y=-0.025
+ $X2=3.662 $Y2=2.03
cc_107 N_GND_M1014_b N_A_43_110#_c_900_n 0.0186694f $X=-1.345 $Y=-0.025 $X2=3.75
+ $Y2=1.625
cc_108 N_GND_c_64_p N_A_43_110#_c_900_n 0.00606474f $X=3.905 $Y=0.127 $X2=3.75
+ $Y2=1.625
cc_109 N_GND_c_109_p N_A_43_110#_c_900_n 0.00354579f $X=3.99 $Y=0.8 $X2=3.75
+ $Y2=1.625
cc_110 N_GND_c_4_p N_A_43_110#_c_900_n 0.00468827f $X=5.7 $Y=0.165 $X2=3.75
+ $Y2=1.625
cc_111 N_GND_M1014_b N_A_43_110#_c_904_n 0.0135442f $X=-1.345 $Y=-0.025 $X2=3.75
+ $Y2=1.775
cc_112 N_GND_M1014_b N_A_43_110#_c_905_n 0.0273935f $X=-1.345 $Y=-0.025 $X2=3.75
+ $Y2=2.83
cc_113 N_GND_M1014_b N_A_43_110#_c_906_n 0.00430539f $X=-1.345 $Y=-0.025
+ $X2=3.75 $Y2=2.98
cc_114 N_GND_M1014_b N_A_43_110#_c_907_n 0.0315687f $X=-1.345 $Y=-0.025
+ $X2=0.225 $Y2=2.195
cc_115 N_GND_M1014_b N_A_43_110#_c_908_n 0.00156053f $X=-1.345 $Y=-0.025
+ $X2=0.34 $Y2=0.8
cc_116 N_GND_c_14_p N_A_43_110#_c_908_n 0.031398f $X=-0.179 $Y=0.8 $X2=0.34
+ $Y2=0.8
cc_117 N_GND_c_22_p N_A_43_110#_c_908_n 0.00757793f $X=0.685 $Y=0.127 $X2=0.34
+ $Y2=0.8
cc_118 N_GND_c_4_p N_A_43_110#_c_908_n 0.00476261f $X=5.7 $Y=0.165 $X2=0.34
+ $Y2=0.8
cc_119 N_GND_M1014_b N_A_43_110#_c_912_n 0.00366408f $X=-1.345 $Y=-0.025
+ $X2=2.365 $Y2=2.195
cc_120 N_GND_M1014_b N_A_43_110#_c_913_n 0.00272681f $X=-1.345 $Y=-0.025
+ $X2=3.66 $Y2=2.195
cc_121 N_GND_M1014_b N_A_43_110#_c_914_n 0.00474188f $X=-1.345 $Y=-0.025
+ $X2=0.34 $Y2=1.37
cc_122 N_GND_c_14_p N_A_43_110#_c_914_n 0.00619665f $X=-0.179 $Y=0.8 $X2=0.34
+ $Y2=1.37
cc_123 N_GND_M1014_b N_A_43_110#_c_916_n 0.0105472f $X=-1.345 $Y=-0.025
+ $X2=3.515 $Y2=2.195
cc_124 N_GND_M1014_b N_A_43_110#_c_917_n 0.00256062f $X=-1.345 $Y=-0.025
+ $X2=2.515 $Y2=2.195
cc_125 N_GND_M1014_b N_A_43_110#_c_918_n 0.0101652f $X=-1.345 $Y=-0.025 $X2=0.37
+ $Y2=2.195
cc_126 N_GND_M1014_b N_A_43_110#_c_919_n 0.0179513f $X=-1.345 $Y=-0.025 $X2=2.22
+ $Y2=2.195
cc_127 N_GND_M1014_b N_A_43_110#_c_920_n 0.00123041f $X=-1.345 $Y=-0.025
+ $X2=3.66 $Y2=2.195
cc_128 N_GND_M1014_b N_A_687_110#_M1009_g 0.0382384f $X=-1.345 $Y=-0.025
+ $X2=4.205 $Y2=1.05
cc_129 N_GND_c_109_p N_A_687_110#_M1009_g 0.00354579f $X=3.99 $Y=0.8 $X2=4.205
+ $Y2=1.05
cc_130 N_GND_c_130_p N_A_687_110#_M1009_g 0.00606474f $X=4.855 $Y=0.127
+ $X2=4.205 $Y2=1.05
cc_131 N_GND_c_131_p N_A_687_110#_M1009_g 0.00463923f $X=4.94 $Y=0.8 $X2=4.205
+ $Y2=1.05
cc_132 N_GND_c_4_p N_A_687_110#_M1009_g 0.00468827f $X=5.7 $Y=0.165 $X2=4.205
+ $Y2=1.05
cc_133 N_GND_M1014_b N_A_687_110#_M1008_g 0.0285283f $X=-1.345 $Y=-0.025
+ $X2=4.205 $Y2=4.56
cc_134 N_GND_M1014_b N_A_687_110#_M1018_g 0.0662302f $X=-1.345 $Y=-0.025
+ $X2=5.155 $Y2=1.05
cc_135 N_GND_c_131_p N_A_687_110#_M1018_g 0.00713292f $X=4.94 $Y=0.8 $X2=5.155
+ $Y2=1.05
cc_136 N_GND_c_79_p N_A_687_110#_M1018_g 0.00606474f $X=5.715 $Y=0.127 $X2=5.155
+ $Y2=1.05
cc_137 N_GND_c_4_p N_A_687_110#_M1018_g 0.00468827f $X=5.7 $Y=0.165 $X2=5.155
+ $Y2=1.05
cc_138 N_GND_M1014_b N_A_687_110#_M1016_g 0.0039012f $X=-1.345 $Y=-0.025
+ $X2=5.155 $Y2=4.56
cc_139 N_GND_M1014_b N_A_687_110#_c_1076_n 0.0289774f $X=-1.345 $Y=-0.025
+ $X2=4.145 $Y2=2.195
cc_140 N_GND_M1014_b N_A_687_110#_c_1077_n 0.0430788f $X=-1.345 $Y=-0.025
+ $X2=5.155 $Y2=2.65
cc_141 N_GND_M1014_b N_A_687_110#_c_1078_n 0.00538086f $X=-1.345 $Y=-0.025
+ $X2=3.56 $Y2=0.8
cc_142 N_GND_c_64_p N_A_687_110#_c_1078_n 0.00745733f $X=3.905 $Y=0.127 $X2=3.56
+ $Y2=0.8
cc_143 N_GND_c_4_p N_A_687_110#_c_1078_n 0.00476261f $X=5.7 $Y=0.165 $X2=3.56
+ $Y2=0.8
cc_144 N_GND_M1014_b N_A_687_110#_c_1081_n 8.75823e-19 $X=-1.345 $Y=-0.025
+ $X2=3.56 $Y2=2.935
cc_145 N_GND_M1014_b N_A_687_110#_c_1082_n 0.00981319f $X=-1.345 $Y=-0.025
+ $X2=4.06 $Y2=1.825
cc_146 N_GND_c_109_p N_A_687_110#_c_1082_n 0.00827205f $X=3.99 $Y=0.8 $X2=4.06
+ $Y2=1.825
cc_147 N_GND_M1014_b N_A_687_110#_c_1084_n 0.00298083f $X=-1.345 $Y=-0.025
+ $X2=3.645 $Y2=1.825
cc_148 N_GND_M1014_b N_A_687_110#_c_1085_n 0.00512756f $X=-1.345 $Y=-0.025
+ $X2=4.06 $Y2=2.74
cc_149 N_GND_M1014_b N_A_687_110#_c_1086_n 0.00247863f $X=-1.345 $Y=-0.025
+ $X2=3.645 $Y2=2.74
cc_150 N_GND_M1014_b N_A_687_110#_c_1087_n 0.0046369f $X=-1.345 $Y=-0.025
+ $X2=4.145 $Y2=2.195
cc_151 N_GND_M1014_b N_A_687_110#_c_1088_n 0.00277707f $X=-1.345 $Y=-0.025
+ $X2=4.95 $Y2=2.65
cc_152 N_GND_M1014_b N_A_687_110#_c_1089_n 0.00492989f $X=-1.345 $Y=-0.025
+ $X2=4.805 $Y2=2.935
cc_153 N_GND_M1014_b N_A_687_110#_c_1090_n 0.00187131f $X=-1.345 $Y=-0.025
+ $X2=3.705 $Y2=2.935
cc_154 N_GND_M1014_b N_A_963_612#_M1013_g 0.0277213f $X=-1.345 $Y=-0.025
+ $X2=6.015 $Y2=1.05
cc_155 N_GND_c_80_p N_A_963_612#_M1013_g 0.00354579f $X=5.8 $Y=0.8 $X2=6.015
+ $Y2=1.05
cc_156 N_GND_c_156_p N_A_963_612#_M1013_g 0.00606474f $X=5.8 $Y=0.127 $X2=6.015
+ $Y2=1.05
cc_157 N_GND_c_4_p N_A_963_612#_M1013_g 0.00468827f $X=5.7 $Y=0.165 $X2=6.015
+ $Y2=1.05
cc_158 N_GND_M1014_b N_A_963_612#_c_1191_n 0.0364586f $X=-1.345 $Y=-0.025
+ $X2=6.05 $Y2=2.075
cc_159 N_GND_M1014_b N_A_963_612#_c_1192_n 0.0466273f $X=-1.345 $Y=-0.025
+ $X2=6.032 $Y2=2.785
cc_160 N_GND_M1014_b N_A_963_612#_c_1193_n 0.0076653f $X=-1.345 $Y=-0.025
+ $X2=6.032 $Y2=2.935
cc_161 N_GND_M1014_b N_A_963_612#_c_1194_n 0.00541552f $X=-1.345 $Y=-0.025
+ $X2=5.29 $Y2=3.52
cc_162 N_GND_M1014_b N_A_963_612#_c_1195_n 0.00710171f $X=-1.345 $Y=-0.025
+ $X2=5.37 $Y2=0.8
cc_163 N_GND_c_79_p N_A_963_612#_c_1195_n 0.0075556f $X=5.715 $Y=0.127 $X2=5.37
+ $Y2=0.8
cc_164 N_GND_c_4_p N_A_963_612#_c_1195_n 0.00475776f $X=5.7 $Y=0.165 $X2=5.37
+ $Y2=0.8
cc_165 N_GND_M1014_b N_A_963_612#_c_1198_n 0.0187633f $X=-1.345 $Y=-0.025
+ $X2=6.11 $Y2=1.91
cc_166 N_GND_c_80_p N_A_963_612#_c_1198_n 0.00702738f $X=5.8 $Y=0.8 $X2=6.11
+ $Y2=1.91
cc_167 N_GND_M1014_b N_A_963_612#_c_1200_n 0.00371235f $X=-1.345 $Y=-0.025
+ $X2=5.33 $Y2=1.91
cc_168 N_GND_M1014_b N_A_856_110#_c_1269_n 0.00156053f $X=-1.345 $Y=-0.025
+ $X2=4.42 $Y2=0.8
cc_169 N_GND_c_130_p N_A_856_110#_c_1269_n 0.00757793f $X=4.855 $Y=0.127
+ $X2=4.42 $Y2=0.8
cc_170 N_GND_c_131_p N_A_856_110#_c_1269_n 0.0358835f $X=4.94 $Y=0.8 $X2=4.42
+ $Y2=0.8
cc_171 N_GND_c_4_p N_A_856_110#_c_1269_n 0.00476261f $X=5.7 $Y=0.165 $X2=4.42
+ $Y2=0.8
cc_172 N_GND_M1014_b N_A_856_110#_c_1273_n 0.0063317f $X=-1.345 $Y=-0.025
+ $X2=4.452 $Y2=1.57
cc_173 N_GND_M1014_b N_A_856_110#_c_1274_n 0.0294549f $X=-1.345 $Y=-0.025
+ $X2=4.452 $Y2=3.135
cc_174 N_GND_M1014_b N_ECK_c_1304_n 0.00156053f $X=-1.345 $Y=-0.025 $X2=6.23
+ $Y2=0.8
cc_175 N_GND_c_156_p N_ECK_c_1304_n 0.00757793f $X=5.8 $Y=0.127 $X2=6.23 $Y2=0.8
cc_176 N_GND_c_4_p N_ECK_c_1304_n 0.00476261f $X=5.7 $Y=0.165 $X2=6.23 $Y2=0.8
cc_177 N_GND_M1014_b N_ECK_c_1307_n 0.016457f $X=-1.345 $Y=-0.025 $X2=6.23
+ $Y2=2.565
cc_178 N_GND_M1014_b N_ECK_c_1308_n 0.039938f $X=-1.345 $Y=-0.025 $X2=6.23
+ $Y2=2.45
cc_179 N_GND_M1014_b N_ECK_c_1309_n 0.0121687f $X=-1.345 $Y=-0.025 $X2=6.23
+ $Y2=1.455
cc_180 N_GND_c_80_p N_ECK_c_1309_n 0.00125659f $X=5.8 $Y=0.8 $X2=6.23 $Y2=1.455
cc_181 N_GND_M1014_b ECK 0.0141689f $X=-1.345 $Y=-0.025 $X2=6.23 $Y2=2.565
cc_182 N_VDD_M1011_b N_SE_M1011_g 0.0246289f $X=-1.345 $Y=2.88 $X2=-0.825
+ $Y2=4.56
cc_183 N_VDD_c_183_p N_SE_M1011_g 0.00606474f $X=-0.335 $Y=6.482 $X2=-0.825
+ $Y2=4.56
cc_184 N_VDD_c_184_p N_SE_M1011_g 0.00468827f $X=5.7 $Y=6.445 $X2=-0.825
+ $Y2=4.56
cc_185 N_VDD_M1011_b N_SE_c_299_n 0.00408216f $X=-1.345 $Y=2.88 $X2=-0.649
+ $Y2=2.935
cc_186 N_VDD_M1011_b N_SE_X27_noxref_CONDUCTOR 0.00838127f $X=-1.345 $Y=2.88
+ $X2=-0.649 $Y2=2.935
cc_187 N_VDD_M1011_b N_E_M1017_g 0.0199366f $X=-1.345 $Y=2.88 $X2=-0.465
+ $Y2=4.56
cc_188 N_VDD_c_183_p N_E_M1017_g 0.00606474f $X=-0.335 $Y=6.482 $X2=-0.465
+ $Y2=4.56
cc_189 N_VDD_c_189_p N_E_M1017_g 0.00713292f $X=-0.249 $Y=4.11 $X2=-0.465
+ $Y2=4.56
cc_190 N_VDD_c_184_p N_E_M1017_g 0.00468827f $X=5.7 $Y=6.445 $X2=-0.465 $Y2=4.56
cc_191 N_VDD_M1011_b N_E_c_344_n 0.007742f $X=-1.345 $Y=2.88 $X2=-0.309 $Y2=2.73
cc_192 N_VDD_M1017_d N_E_c_345_n 0.00499194f $X=-0.39 $Y=3.06 $X2=-0.309
+ $Y2=2.73
cc_193 N_VDD_M1011_b N_E_c_345_n 0.00192816f $X=-1.345 $Y=2.88 $X2=-0.309
+ $Y2=2.73
cc_194 N_VDD_c_189_p N_E_c_345_n 0.00252874f $X=-0.249 $Y=4.11 $X2=-0.309
+ $Y2=2.73
cc_195 N_VDD_M1017_d E 0.00723173f $X=-0.39 $Y=3.06 $X2=-0.305 $Y2=3.3
cc_196 N_VDD_c_189_p E 0.00522047f $X=-0.249 $Y=4.11 $X2=-0.305 $Y2=3.3
cc_197 N_VDD_M1011_b N_A_86_332#_c_395_n 0.02482f $X=-1.345 $Y=2.88 $X2=0.53
+ $Y2=2.95
cc_198 N_VDD_c_189_p N_A_86_332#_c_395_n 0.00742312f $X=-0.249 $Y=4.11 $X2=0.53
+ $Y2=2.95
cc_199 N_VDD_c_199_p N_A_86_332#_c_395_n 0.00606474f $X=0.685 $Y=6.482 $X2=0.53
+ $Y2=2.95
cc_200 N_VDD_c_200_p N_A_86_332#_c_395_n 0.00354579f $X=0.77 $Y=3.77 $X2=0.53
+ $Y2=2.95
cc_201 N_VDD_c_184_p N_A_86_332#_c_395_n 0.00468827f $X=5.7 $Y=6.445 $X2=0.53
+ $Y2=2.95
cc_202 N_VDD_M1011_b N_A_86_332#_c_397_n 0.00184258f $X=-1.345 $Y=2.88 $X2=0.565
+ $Y2=3.075
cc_203 N_VDD_M1001_d N_A_86_332#_c_410_n 0.00445123f $X=0.63 $Y=3.06 $X2=1.475
+ $Y2=3.16
cc_204 N_VDD_c_200_p N_A_86_332#_c_410_n 0.00946335f $X=0.77 $Y=3.77 $X2=1.475
+ $Y2=3.16
cc_205 N_VDD_M1011_b N_A_86_332#_c_412_n 0.00313975f $X=-1.345 $Y=2.88 $X2=1.645
+ $Y2=3.43
cc_206 N_VDD_c_206_p N_A_86_332#_c_412_n 0.0151591f $X=2.435 $Y=6.482 $X2=1.645
+ $Y2=3.43
cc_207 N_VDD_c_184_p N_A_86_332#_c_412_n 0.00958198f $X=5.7 $Y=6.445 $X2=1.645
+ $Y2=3.43
cc_208 N_VDD_M1011_b N_A_N233_612#_M1000_g 0.0197362f $X=-1.345 $Y=2.88
+ $X2=0.985 $Y2=4.56
cc_209 N_VDD_c_200_p N_A_N233_612#_M1000_g 0.00354579f $X=0.77 $Y=3.77 $X2=0.985
+ $Y2=4.56
cc_210 N_VDD_c_206_p N_A_N233_612#_M1000_g 0.00606474f $X=2.435 $Y=6.482
+ $X2=0.985 $Y2=4.56
cc_211 N_VDD_c_184_p N_A_N233_612#_M1000_g 0.00468827f $X=5.7 $Y=6.445 $X2=0.985
+ $Y2=4.56
cc_212 N_VDD_M1011_b N_A_N233_612#_c_476_n 0.00981538f $X=-1.345 $Y=2.88
+ $X2=-1.039 $Y2=2.565
cc_213 N_VDD_c_183_p N_A_N233_612#_c_476_n 0.00736239f $X=-0.335 $Y=6.482
+ $X2=-1.039 $Y2=2.565
cc_214 N_VDD_c_184_p N_A_N233_612#_c_476_n 0.00476261f $X=5.7 $Y=6.445
+ $X2=-1.039 $Y2=2.565
cc_215 N_VDD_M1011_b N_A_254_515#_M1023_g 0.0201267f $X=-1.345 $Y=2.88 $X2=1.345
+ $Y2=4.56
cc_216 N_VDD_c_206_p N_A_254_515#_M1023_g 0.00606474f $X=2.435 $Y=6.482
+ $X2=1.345 $Y2=4.56
cc_217 N_VDD_c_184_p N_A_254_515#_M1023_g 0.00468827f $X=5.7 $Y=6.445 $X2=1.345
+ $Y2=4.56
cc_218 N_VDD_M1011_b N_A_254_515#_c_574_n 0.00444465f $X=-1.345 $Y=2.88
+ $X2=1.405 $Y2=2.74
cc_219 N_VDD_M1011_b N_A_254_515#_c_595_n 0.00156053f $X=-1.345 $Y=2.88 $X2=2.95
+ $Y2=3.43
cc_220 N_VDD_c_220_p N_A_254_515#_c_595_n 0.00754714f $X=3.905 $Y=6.482 $X2=2.95
+ $Y2=3.43
cc_221 N_VDD_c_184_p N_A_254_515#_c_595_n 0.00476261f $X=5.7 $Y=6.445 $X2=2.95
+ $Y2=3.43
cc_222 N_VDD_M1011_b N_A_254_515#_c_587_n 0.00468773f $X=-1.345 $Y=2.88 $X2=3.22
+ $Y2=3.075
cc_223 N_VDD_M1011_b N_A_254_515#_c_599_n 0.0117651f $X=-1.345 $Y=2.88 $X2=3.22
+ $Y2=3.16
cc_224 N_VDD_M1011_b N_CK_M1012_g 0.020128f $X=-1.345 $Y=2.88 $X2=1.945 $Y2=4.56
cc_225 N_VDD_c_206_p N_CK_M1012_g 0.00606474f $X=2.435 $Y=6.482 $X2=1.945
+ $Y2=4.56
cc_226 N_VDD_c_184_p N_CK_M1012_g 0.00468827f $X=5.7 $Y=6.445 $X2=1.945 $Y2=4.56
cc_227 N_VDD_M1011_b N_CK_c_705_n 0.00776576f $X=-1.345 $Y=2.88 $X2=2.735
+ $Y2=2.905
cc_228 N_VDD_M1011_b N_CK_M1006_g 0.0237243f $X=-1.345 $Y=2.88 $X2=2.735
+ $Y2=4.56
cc_229 N_VDD_c_229_p N_CK_M1006_g 0.00354579f $X=2.52 $Y=3.43 $X2=2.735 $Y2=4.56
cc_230 N_VDD_c_220_p N_CK_M1006_g 0.00606474f $X=3.905 $Y=6.482 $X2=2.735
+ $Y2=4.56
cc_231 N_VDD_c_184_p N_CK_M1006_g 0.00468827f $X=5.7 $Y=6.445 $X2=2.735 $Y2=4.56
cc_232 N_VDD_M1011_b N_CK_M1020_g 0.0195137f $X=-1.345 $Y=2.88 $X2=5.585
+ $Y2=4.56
cc_233 N_VDD_c_233_p N_CK_M1020_g 0.00606474f $X=5.715 $Y=6.482 $X2=5.585
+ $Y2=4.56
cc_234 N_VDD_c_234_p N_CK_M1020_g 0.00354579f $X=5.8 $Y=4.11 $X2=5.585 $Y2=4.56
cc_235 N_VDD_c_184_p N_CK_M1020_g 0.00468827f $X=5.7 $Y=6.445 $X2=5.585 $Y2=4.56
cc_236 N_VDD_M1011_b N_CK_c_712_n 0.00484874f $X=-1.345 $Y=2.88 $X2=1.885
+ $Y2=2.74
cc_237 N_VDD_M1011_b N_CK_c_720_n 0.0022456f $X=-1.345 $Y=2.88 $X2=1.885
+ $Y2=2.565
cc_238 N_VDD_M1011_b N_CK_c_721_n 0.00302835f $X=-1.345 $Y=2.88 $X2=2.88
+ $Y2=2.565
cc_239 N_VDD_M1011_b N_CK_c_722_n 0.00153494f $X=-1.345 $Y=2.88 $X2=5.63
+ $Y2=2.36
cc_240 N_VDD_M1020_d N_CK_c_744_n 0.00612903f $X=5.66 $Y=3.06 $X2=5.63 $Y2=2.565
cc_241 N_VDD_c_234_p N_CK_c_744_n 0.00247404f $X=5.8 $Y=4.11 $X2=5.63 $Y2=2.565
cc_242 N_VDD_c_229_p N_CK_c_723_n 0.00634153f $X=2.52 $Y=3.43 $X2=2.735
+ $Y2=2.565
cc_243 N_VDD_M1011_b N_A_43_110#_M1004_g 0.0197647f $X=-1.345 $Y=2.88 $X2=2.305
+ $Y2=4.56
cc_244 N_VDD_c_206_p N_A_43_110#_M1004_g 0.00606474f $X=2.435 $Y=6.482 $X2=2.305
+ $Y2=4.56
cc_245 N_VDD_c_229_p N_A_43_110#_M1004_g 0.00354579f $X=2.52 $Y=3.43 $X2=2.305
+ $Y2=4.56
cc_246 N_VDD_c_184_p N_A_43_110#_M1004_g 0.00468827f $X=5.7 $Y=6.445 $X2=2.305
+ $Y2=4.56
cc_247 N_VDD_M1011_b N_A_43_110#_c_906_n 0.0279523f $X=-1.345 $Y=2.88 $X2=3.75
+ $Y2=2.98
cc_248 N_VDD_c_220_p N_A_43_110#_c_906_n 0.00606474f $X=3.905 $Y=6.482 $X2=3.75
+ $Y2=2.98
cc_249 N_VDD_c_249_p N_A_43_110#_c_906_n 0.00354579f $X=3.99 $Y=3.43 $X2=3.75
+ $Y2=2.98
cc_250 N_VDD_c_184_p N_A_43_110#_c_906_n 0.00468827f $X=5.7 $Y=6.445 $X2=3.75
+ $Y2=2.98
cc_251 N_VDD_M1011_b N_A_43_110#_c_907_n 0.00930728f $X=-1.345 $Y=2.88 $X2=0.225
+ $Y2=2.195
cc_252 N_VDD_M1011_b N_A_43_110#_c_930_n 0.00156053f $X=-1.345 $Y=2.88 $X2=0.34
+ $Y2=4.11
cc_253 N_VDD_c_189_p N_A_43_110#_c_930_n 0.0794385f $X=-0.249 $Y=4.11 $X2=0.34
+ $Y2=4.11
cc_254 N_VDD_c_199_p N_A_43_110#_c_930_n 0.00757793f $X=0.685 $Y=6.482 $X2=0.34
+ $Y2=4.11
cc_255 N_VDD_c_184_p N_A_43_110#_c_930_n 0.00476261f $X=5.7 $Y=6.445 $X2=0.34
+ $Y2=4.11
cc_256 N_VDD_M1011_b N_A_43_110#_c_934_n 0.00962373f $X=-1.345 $Y=2.88 $X2=0.34
+ $Y2=3.77
cc_257 N_VDD_c_189_p N_A_43_110#_c_934_n 0.00355502f $X=-0.249 $Y=4.11 $X2=0.34
+ $Y2=3.77
cc_258 N_VDD_M1011_b N_A_687_110#_M1008_g 0.0256676f $X=-1.345 $Y=2.88 $X2=4.205
+ $Y2=4.56
cc_259 N_VDD_c_249_p N_A_687_110#_M1008_g 0.00354579f $X=3.99 $Y=3.43 $X2=4.205
+ $Y2=4.56
cc_260 N_VDD_c_233_p N_A_687_110#_M1008_g 0.00606474f $X=5.715 $Y=6.482
+ $X2=4.205 $Y2=4.56
cc_261 N_VDD_c_184_p N_A_687_110#_M1008_g 0.00468827f $X=5.7 $Y=6.445 $X2=4.205
+ $Y2=4.56
cc_262 N_VDD_M1011_b N_A_687_110#_M1016_g 0.0258226f $X=-1.345 $Y=2.88 $X2=5.155
+ $Y2=4.56
cc_263 N_VDD_c_233_p N_A_687_110#_M1016_g 0.00606474f $X=5.715 $Y=6.482
+ $X2=5.155 $Y2=4.56
cc_264 N_VDD_c_184_p N_A_687_110#_M1016_g 0.00468827f $X=5.7 $Y=6.445 $X2=5.155
+ $Y2=4.56
cc_265 N_VDD_M1011_b N_A_687_110#_c_1081_n 0.00482437f $X=-1.345 $Y=2.88
+ $X2=3.56 $Y2=2.935
cc_266 N_VDD_c_220_p N_A_687_110#_c_1081_n 0.00745733f $X=3.905 $Y=6.482
+ $X2=3.56 $Y2=2.935
cc_267 N_VDD_c_184_p N_A_687_110#_c_1081_n 0.00476261f $X=5.7 $Y=6.445 $X2=3.56
+ $Y2=2.935
cc_268 N_VDD_c_249_p N_A_687_110#_c_1085_n 0.00435485f $X=3.99 $Y=3.43 $X2=4.06
+ $Y2=2.74
cc_269 N_VDD_M1011_b N_A_687_110#_c_1088_n 0.00272119f $X=-1.345 $Y=2.88
+ $X2=4.95 $Y2=2.65
cc_270 N_VDD_M1011_b N_A_687_110#_c_1089_n 0.0191595f $X=-1.345 $Y=2.88
+ $X2=4.805 $Y2=2.935
cc_271 N_VDD_c_249_p N_A_687_110#_c_1089_n 0.00518939f $X=3.99 $Y=3.43 $X2=4.805
+ $Y2=2.935
cc_272 N_VDD_M1011_b N_A_687_110#_c_1090_n 0.00976168f $X=-1.345 $Y=2.88
+ $X2=3.705 $Y2=2.935
cc_273 N_VDD_M1011_b N_A_963_612#_c_1193_n 0.0267159f $X=-1.345 $Y=2.88
+ $X2=6.032 $Y2=2.935
cc_274 N_VDD_c_234_p N_A_963_612#_c_1193_n 0.00354579f $X=5.8 $Y=4.11 $X2=6.032
+ $Y2=2.935
cc_275 N_VDD_c_275_p N_A_963_612#_c_1193_n 0.00606474f $X=5.8 $Y=6.482 $X2=6.032
+ $Y2=2.935
cc_276 N_VDD_c_184_p N_A_963_612#_c_1193_n 0.00468827f $X=5.7 $Y=6.445 $X2=6.032
+ $Y2=2.935
cc_277 N_VDD_M1011_b N_A_963_612#_c_1205_n 0.00156053f $X=-1.345 $Y=2.88
+ $X2=4.94 $Y2=3.77
cc_278 N_VDD_c_233_p N_A_963_612#_c_1205_n 0.00736239f $X=5.715 $Y=6.482
+ $X2=4.94 $Y2=3.77
cc_279 N_VDD_c_184_p N_A_963_612#_c_1205_n 0.00476261f $X=5.7 $Y=6.445 $X2=4.94
+ $Y2=3.77
cc_280 N_VDD_M1011_b N_A_963_612#_c_1194_n 0.00106577f $X=-1.345 $Y=2.88
+ $X2=5.29 $Y2=3.52
cc_281 N_VDD_M1011_b N_A_856_110#_c_1275_n 0.00514058f $X=-1.345 $Y=2.88
+ $X2=4.42 $Y2=3.305
cc_282 N_VDD_c_249_p N_A_856_110#_c_1275_n 0.00677841f $X=3.99 $Y=3.43 $X2=4.42
+ $Y2=3.305
cc_283 N_VDD_M1011_b N_A_856_110#_c_1277_n 0.00156053f $X=-1.345 $Y=2.88
+ $X2=4.42 $Y2=3.43
cc_284 N_VDD_c_233_p N_A_856_110#_c_1277_n 0.00757793f $X=5.715 $Y=6.482
+ $X2=4.42 $Y2=3.43
cc_285 N_VDD_c_184_p N_A_856_110#_c_1277_n 0.00476261f $X=5.7 $Y=6.445 $X2=4.42
+ $Y2=3.43
cc_286 N_VDD_M1011_b N_A_856_110#_c_1274_n 0.00534142f $X=-1.345 $Y=2.88
+ $X2=4.452 $Y2=3.135
cc_287 N_VDD_M1011_b N_ECK_c_1307_n 0.010295f $X=-1.345 $Y=2.88 $X2=6.23
+ $Y2=2.565
cc_288 N_VDD_c_275_p N_ECK_c_1307_n 0.00757793f $X=5.8 $Y=6.482 $X2=6.23
+ $Y2=2.565
cc_289 N_VDD_c_184_p N_ECK_c_1307_n 0.00476261f $X=5.7 $Y=6.445 $X2=6.23
+ $Y2=2.565
cc_290 N_SE_X27_noxref_CONDUCTOR N_E_M1017_g 0.00231474f $X=-0.649 $Y=2.935
+ $X2=-0.465 $Y2=4.56
cc_291 N_SE_M1014_g N_E_M1024_g 0.060867f $X=-0.825 $Y=1.05 $X2=-0.395 $Y2=1.05
cc_292 N_SE_c_297_n N_E_M1024_g 0.00368334f $X=-0.735 $Y=2.065 $X2=-0.395
+ $Y2=1.05
cc_293 N_SE_c_299_n N_E_M1024_g 0.00800257f $X=-0.649 $Y=2.935 $X2=-0.395
+ $Y2=1.05
cc_294 N_SE_M1011_g N_E_c_344_n 0.217191f $X=-0.825 $Y=4.56 $X2=-0.309 $Y2=2.73
cc_295 N_SE_c_299_n N_E_c_344_n 0.00287728f $X=-0.649 $Y=2.935 $X2=-0.309
+ $Y2=2.73
cc_296 N_SE_X27_noxref_CONDUCTOR N_E_c_344_n 0.00131279f $X=-0.649 $Y=2.935
+ $X2=-0.309 $Y2=2.73
cc_297 N_SE_M1011_g N_E_c_345_n 0.00140064f $X=-0.825 $Y=4.56 $X2=-0.309
+ $Y2=2.73
cc_298 N_SE_c_299_n N_E_c_345_n 0.0302287f $X=-0.649 $Y=2.935 $X2=-0.309
+ $Y2=2.73
cc_299 N_SE_X27_noxref_CONDUCTOR N_E_c_345_n 0.00643447f $X=-0.649 $Y=2.935
+ $X2=-0.309 $Y2=2.73
cc_300 N_SE_M1011_g E 0.00297933f $X=-0.825 $Y=4.56 $X2=-0.305 $Y2=3.3
cc_301 N_SE_X27_noxref_CONDUCTOR E 0.0050603f $X=-0.649 $Y=2.935 $X2=-0.305
+ $Y2=3.3
cc_302 N_SE_M1011_g N_A_N233_612#_c_476_n 0.016616f $X=-0.825 $Y=4.56 $X2=-1.039
+ $Y2=2.565
cc_303 N_SE_c_295_n N_A_N233_612#_c_476_n 0.00138434f $X=-0.884 $Y=2.065
+ $X2=-1.039 $Y2=2.565
cc_304 N_SE_c_297_n N_A_N233_612#_c_476_n 0.00308264f $X=-0.735 $Y=2.065
+ $X2=-1.039 $Y2=2.565
cc_305 N_SE_c_299_n N_A_N233_612#_c_476_n 0.0294278f $X=-0.649 $Y=2.935
+ $X2=-1.039 $Y2=2.565
cc_306 N_SE_X27_noxref_CONDUCTOR N_A_N233_612#_c_476_n 0.00774605f $X=-0.649
+ $Y=2.935 $X2=-1.039 $Y2=2.565
cc_307 N_SE_M1014_g N_A_N233_612#_c_477_n 0.00231637f $X=-0.825 $Y=1.05
+ $X2=-0.609 $Y2=0.8
cc_308 N_SE_c_297_n N_A_N233_612#_c_477_n 0.00336259f $X=-0.735 $Y=2.065
+ $X2=-0.609 $Y2=0.8
cc_309 N_SE_M1011_g N_A_N233_612#_c_481_n 0.00412998f $X=-0.825 $Y=4.56
+ $X2=-0.695 $Y2=2.565
cc_310 N_SE_c_297_n N_A_N233_612#_c_481_n 0.00523952f $X=-0.735 $Y=2.065
+ $X2=-0.695 $Y2=2.565
cc_311 N_SE_c_299_n N_A_N233_612#_c_481_n 0.00526709f $X=-0.649 $Y=2.935
+ $X2=-0.695 $Y2=2.565
cc_312 N_SE_X27_noxref_CONDUCTOR N_A_N233_612#_c_481_n 0.0344998f $X=-0.649
+ $Y=2.935 $X2=-0.695 $Y2=2.565
cc_313 N_SE_M1011_g N_A_N233_612#_c_482_n 0.00327819f $X=-0.825 $Y=4.56
+ $X2=-0.895 $Y2=2.565
cc_314 N_SE_c_295_n N_A_N233_612#_c_482_n 0.00301446f $X=-0.884 $Y=2.065
+ $X2=-0.895 $Y2=2.565
cc_315 N_SE_c_297_n N_A_N233_612#_c_482_n 0.00469337f $X=-0.735 $Y=2.065
+ $X2=-0.895 $Y2=2.565
cc_316 N_SE_c_299_n N_A_N233_612#_c_482_n 0.00157282f $X=-0.649 $Y=2.935
+ $X2=-0.895 $Y2=2.565
cc_317 N_SE_X27_noxref_CONDUCTOR N_A_N233_612#_c_482_n 9.25684e-19 $X=-0.649
+ $Y=2.935 $X2=-0.895 $Y2=2.565
cc_318 N_SE_M1014_g N_A_N233_612#_c_483_n 0.00594872f $X=-0.825 $Y=1.05
+ $X2=-0.61 $Y2=2.48
cc_319 N_SE_c_297_n N_A_N233_612#_c_483_n 0.0124433f $X=-0.735 $Y=2.065
+ $X2=-0.61 $Y2=2.48
cc_320 N_SE_c_299_n N_A_N233_612#_c_483_n 0.0178687f $X=-0.649 $Y=2.935
+ $X2=-0.61 $Y2=2.48
cc_321 N_SE_M1014_g N_A_N233_612#_c_485_n 0.0089989f $X=-0.825 $Y=1.05
+ $X2=-0.609 $Y2=1.455
cc_322 N_SE_c_297_n N_A_N233_612#_c_485_n 0.00244196f $X=-0.735 $Y=2.065
+ $X2=-0.609 $Y2=1.455
cc_323 N_SE_c_299_n N_A_N233_612#_c_488_n 0.0081604f $X=-0.649 $Y=2.935
+ $X2=-0.61 $Y2=2.565
cc_324 N_E_c_344_n N_A_86_332#_c_394_n 0.00466473f $X=-0.309 $Y=2.73 $X2=0.53
+ $Y2=2.78
cc_325 N_E_c_345_n N_A_N233_612#_c_476_n 0.00350166f $X=-0.309 $Y=2.73
+ $X2=-1.039 $Y2=2.565
cc_326 E N_A_N233_612#_c_476_n 0.00623956f $X=-0.305 $Y=3.3 $X2=-1.039 $Y2=2.565
cc_327 N_E_M1024_g N_A_N233_612#_c_477_n 0.00162674f $X=-0.395 $Y=1.05
+ $X2=-0.609 $Y2=0.8
cc_328 N_E_M1024_g N_A_N233_612#_c_483_n 0.013109f $X=-0.395 $Y=1.05 $X2=-0.61
+ $Y2=2.48
cc_329 N_E_M1024_g N_A_N233_612#_c_484_n 0.00815941f $X=-0.395 $Y=1.05 $X2=0.78
+ $Y2=2.565
cc_330 N_E_c_344_n N_A_N233_612#_c_484_n 0.00669754f $X=-0.309 $Y=2.73 $X2=0.78
+ $Y2=2.565
cc_331 N_E_c_345_n N_A_N233_612#_c_484_n 0.0110811f $X=-0.309 $Y=2.73 $X2=0.78
+ $Y2=2.565
cc_332 E N_A_N233_612#_c_484_n 0.0125691f $X=-0.305 $Y=3.3 $X2=0.78 $Y2=2.565
cc_333 N_E_M1024_g N_A_N233_612#_c_485_n 0.00476605f $X=-0.395 $Y=1.05
+ $X2=-0.609 $Y2=1.455
cc_334 N_E_c_344_n N_A_N233_612#_c_488_n 8.16409e-19 $X=-0.309 $Y=2.73 $X2=-0.61
+ $Y2=2.565
cc_335 N_E_M1017_g N_A_43_110#_c_907_n 0.0137937f $X=-0.465 $Y=4.56 $X2=0.225
+ $Y2=2.195
cc_336 N_E_M1024_g N_A_43_110#_c_907_n 0.0254566f $X=-0.395 $Y=1.05 $X2=0.225
+ $Y2=2.195
cc_337 N_E_c_344_n N_A_43_110#_c_907_n 0.00283097f $X=-0.309 $Y=2.73 $X2=0.225
+ $Y2=2.195
cc_338 N_E_c_345_n N_A_43_110#_c_907_n 0.0310495f $X=-0.309 $Y=2.73 $X2=0.225
+ $Y2=2.195
cc_339 E N_A_43_110#_c_907_n 0.00692722f $X=-0.305 $Y=3.3 $X2=0.225 $Y2=2.195
cc_340 N_E_M1024_g N_A_43_110#_c_914_n 0.00130963f $X=-0.395 $Y=1.05 $X2=0.34
+ $Y2=1.37
cc_341 N_E_M1024_g N_A_43_110#_c_918_n 0.00532884f $X=-0.395 $Y=1.05 $X2=0.37
+ $Y2=2.195
cc_342 E A_N150_612# 0.00289505f $X=-0.305 $Y=3.3 $X2=-0.75 $Y2=3.06
cc_343 N_A_86_332#_c_387_n N_A_N233_612#_M1002_g 0.0207333f $X=0.565 $Y=1.825
+ $X2=0.985 $Y2=1.05
cc_344 N_A_86_332#_c_389_n N_A_N233_612#_M1002_g 0.0196577f $X=0.565 $Y=1.66
+ $X2=0.985 $Y2=1.05
cc_345 N_A_86_332#_c_394_n N_A_N233_612#_M1002_g 0.00885564f $X=0.53 $Y=2.78
+ $X2=0.985 $Y2=1.05
cc_346 N_A_86_332#_c_396_n N_A_N233_612#_M1002_g 2.45848e-19 $X=0.565 $Y=1.91
+ $X2=0.985 $Y2=1.05
cc_347 N_A_86_332#_c_397_n N_A_N233_612#_M1002_g 0.00448652f $X=0.565 $Y=3.075
+ $X2=0.985 $Y2=1.05
cc_348 N_A_86_332#_c_398_n N_A_N233_612#_M1002_g 0.0125105f $X=1.025 $Y=1.825
+ $X2=0.985 $Y2=1.05
cc_349 N_A_86_332#_c_400_n N_A_N233_612#_M1002_g 0.00552645f $X=1.11 $Y=1.74
+ $X2=0.985 $Y2=1.05
cc_350 N_A_86_332#_c_423_p N_A_N233_612#_M1002_g 0.00605553f $X=1.195 $Y=1.405
+ $X2=0.985 $Y2=1.05
cc_351 N_A_86_332#_c_394_n N_A_N233_612#_M1000_g 0.00755439f $X=0.53 $Y=2.78
+ $X2=0.985 $Y2=4.56
cc_352 N_A_86_332#_c_395_n N_A_N233_612#_M1000_g 0.0412319f $X=0.53 $Y=2.95
+ $X2=0.985 $Y2=4.56
cc_353 N_A_86_332#_c_397_n N_A_N233_612#_M1000_g 0.00605772f $X=0.565 $Y=3.075
+ $X2=0.985 $Y2=4.56
cc_354 N_A_86_332#_c_410_n N_A_N233_612#_M1000_g 0.0156361f $X=1.475 $Y=3.16
+ $X2=0.985 $Y2=4.56
cc_355 N_A_86_332#_c_394_n N_A_N233_612#_c_475_n 0.0209207f $X=0.53 $Y=2.78
+ $X2=0.925 $Y2=2.4
cc_356 N_A_86_332#_c_397_n N_A_N233_612#_c_475_n 0.00174544f $X=0.565 $Y=3.075
+ $X2=0.925 $Y2=2.4
cc_357 N_A_86_332#_c_398_n N_A_N233_612#_c_475_n 0.00174867f $X=1.025 $Y=1.825
+ $X2=0.925 $Y2=2.4
cc_358 N_A_86_332#_c_410_n N_A_N233_612#_c_475_n 0.00122128f $X=1.475 $Y=3.16
+ $X2=0.925 $Y2=2.4
cc_359 N_A_86_332#_c_394_n N_A_N233_612#_c_480_n 6.09588e-19 $X=0.53 $Y=2.78
+ $X2=0.925 $Y2=2.4
cc_360 N_A_86_332#_c_397_n N_A_N233_612#_c_480_n 0.0263734f $X=0.565 $Y=3.075
+ $X2=0.925 $Y2=2.4
cc_361 N_A_86_332#_c_398_n N_A_N233_612#_c_480_n 0.00476537f $X=1.025 $Y=1.825
+ $X2=0.925 $Y2=2.4
cc_362 N_A_86_332#_c_410_n N_A_N233_612#_c_480_n 0.00315222f $X=1.475 $Y=3.16
+ $X2=0.925 $Y2=2.4
cc_363 N_A_86_332#_c_394_n N_A_N233_612#_c_484_n 0.00470193f $X=0.53 $Y=2.78
+ $X2=0.78 $Y2=2.565
cc_364 N_A_86_332#_c_397_n N_A_N233_612#_c_484_n 0.0192961f $X=0.565 $Y=3.075
+ $X2=0.78 $Y2=2.565
cc_365 N_A_86_332#_c_410_n N_A_N233_612#_c_484_n 0.0164414f $X=1.475 $Y=3.16
+ $X2=0.78 $Y2=2.565
cc_366 N_A_86_332#_c_410_n N_A_254_515#_M1023_g 0.015571f $X=1.475 $Y=3.16
+ $X2=1.345 $Y2=4.56
cc_367 N_A_86_332#_c_410_n N_A_254_515#_c_574_n 0.00158944f $X=1.475 $Y=3.16
+ $X2=1.405 $Y2=2.74
cc_368 N_A_86_332#_c_441_p N_A_254_515#_c_575_n 0.00158944f $X=1.475 $Y=1.405
+ $X2=1.885 $Y2=1.825
cc_369 N_A_86_332#_c_441_p N_A_254_515#_c_580_n 0.0139878f $X=1.475 $Y=1.405
+ $X2=2.865 $Y2=1.825
cc_370 N_A_86_332#_c_398_n N_A_254_515#_c_582_n 0.0132034f $X=1.025 $Y=1.825
+ $X2=1.57 $Y2=1.825
cc_371 N_A_86_332#_c_441_p N_A_254_515#_c_582_n 0.00917449f $X=1.475 $Y=1.405
+ $X2=1.57 $Y2=1.825
cc_372 N_A_86_332#_c_397_n N_A_254_515#_c_588_n 0.00496637f $X=0.565 $Y=3.075
+ $X2=1.485 $Y2=2.74
cc_373 N_A_86_332#_c_410_n N_A_254_515#_c_588_n 0.0153302f $X=1.475 $Y=3.16
+ $X2=1.485 $Y2=2.74
cc_374 N_A_86_332#_c_398_n N_CK_M1025_g 0.00127357f $X=1.025 $Y=1.825 $X2=1.345
+ $Y2=1.05
cc_375 N_A_86_332#_c_400_n N_CK_M1025_g 0.00554866f $X=1.11 $Y=1.74 $X2=1.345
+ $Y2=1.05
cc_376 N_A_86_332#_c_441_p N_CK_M1025_g 0.0165456f $X=1.475 $Y=1.405 $X2=1.345
+ $Y2=1.05
cc_377 N_A_86_332#_c_410_n N_CK_c_712_n 0.0025652f $X=1.475 $Y=3.16 $X2=1.885
+ $Y2=2.74
cc_378 N_A_86_332#_c_410_n N_CK_c_720_n 0.00103871f $X=1.475 $Y=3.16 $X2=1.885
+ $Y2=2.565
cc_379 N_A_86_332#_c_410_n N_CK_c_724_n 0.00257262f $X=1.475 $Y=3.16 $X2=2.03
+ $Y2=2.565
cc_380 N_A_86_332#_c_387_n N_A_43_110#_c_907_n 0.0225182f $X=0.565 $Y=1.825
+ $X2=0.225 $Y2=2.195
cc_381 N_A_86_332#_c_389_n N_A_43_110#_c_907_n 0.00700162f $X=0.565 $Y=1.66
+ $X2=0.225 $Y2=2.195
cc_382 N_A_86_332#_c_395_n N_A_43_110#_c_907_n 0.0128109f $X=0.53 $Y=2.95
+ $X2=0.225 $Y2=2.195
cc_383 N_A_86_332#_c_396_n N_A_43_110#_c_907_n 0.0193917f $X=0.565 $Y=1.91
+ $X2=0.225 $Y2=2.195
cc_384 N_A_86_332#_c_397_n N_A_43_110#_c_907_n 0.0809249f $X=0.565 $Y=3.075
+ $X2=0.225 $Y2=2.195
cc_385 N_A_86_332#_c_458_p N_A_43_110#_c_907_n 0.0133619f $X=0.65 $Y=3.16
+ $X2=0.225 $Y2=2.195
cc_386 N_A_86_332#_c_394_n N_A_43_110#_c_918_n 0.0022955f $X=0.53 $Y=2.78
+ $X2=0.37 $Y2=2.195
cc_387 N_A_86_332#_c_397_n N_A_43_110#_c_918_n 0.00271681f $X=0.565 $Y=3.075
+ $X2=0.37 $Y2=2.195
cc_388 N_A_86_332#_c_387_n N_A_43_110#_c_919_n 0.00127165f $X=0.565 $Y=1.825
+ $X2=2.22 $Y2=2.195
cc_389 N_A_86_332#_c_394_n N_A_43_110#_c_919_n 0.00421591f $X=0.53 $Y=2.78
+ $X2=2.22 $Y2=2.195
cc_390 N_A_86_332#_c_397_n N_A_43_110#_c_919_n 0.0177917f $X=0.565 $Y=3.075
+ $X2=2.22 $Y2=2.195
cc_391 N_A_86_332#_c_398_n N_A_43_110#_c_919_n 0.021201f $X=1.025 $Y=1.825
+ $X2=2.22 $Y2=2.195
cc_392 N_A_86_332#_c_441_p N_A_43_110#_c_919_n 0.00659867f $X=1.475 $Y=1.405
+ $X2=2.22 $Y2=2.195
cc_393 N_A_86_332#_c_410_n A_212_612# 0.0060995f $X=1.475 $Y=3.16 $X2=1.06
+ $Y2=3.06
cc_394 N_A_86_332#_c_400_n A_212_110# 6.51949e-19 $X=1.11 $Y=1.74 $X2=1.06
+ $Y2=0.55
cc_395 N_A_86_332#_c_441_p A_212_110# 9.96211e-19 $X=1.475 $Y=1.405 $X2=1.06
+ $Y2=0.55
cc_396 N_A_86_332#_c_423_p A_212_110# 0.0034593f $X=1.195 $Y=1.405 $X2=1.06
+ $Y2=0.55
cc_397 N_A_N233_612#_M1000_g N_A_254_515#_c_574_n 0.215574f $X=0.985 $Y=4.56
+ $X2=1.405 $Y2=2.74
cc_398 N_A_N233_612#_c_480_n N_A_254_515#_c_574_n 3.50159e-19 $X=0.925 $Y=2.4
+ $X2=1.405 $Y2=2.74
cc_399 N_A_N233_612#_c_484_n N_A_254_515#_c_574_n 0.00162818f $X=0.78 $Y=2.565
+ $X2=1.405 $Y2=2.74
cc_400 N_A_N233_612#_M1002_g N_A_254_515#_c_579_n 0.00234107f $X=0.985 $Y=1.05
+ $X2=1.485 $Y2=2.655
cc_401 N_A_N233_612#_c_475_n N_A_254_515#_c_579_n 0.00185841f $X=0.925 $Y=2.4
+ $X2=1.485 $Y2=2.655
cc_402 N_A_N233_612#_c_480_n N_A_254_515#_c_579_n 0.0124483f $X=0.925 $Y=2.4
+ $X2=1.485 $Y2=2.655
cc_403 N_A_N233_612#_c_484_n N_A_254_515#_c_579_n 0.00655758f $X=0.78 $Y=2.565
+ $X2=1.485 $Y2=2.655
cc_404 N_A_N233_612#_M1000_g N_A_254_515#_c_588_n 0.00165169f $X=0.985 $Y=4.56
+ $X2=1.485 $Y2=2.74
cc_405 N_A_N233_612#_c_484_n N_A_254_515#_c_588_n 0.00103938f $X=0.78 $Y=2.565
+ $X2=1.485 $Y2=2.74
cc_406 N_A_N233_612#_M1002_g N_CK_M1025_g 0.0581908f $X=0.985 $Y=1.05 $X2=1.345
+ $Y2=1.05
cc_407 N_A_N233_612#_c_475_n N_CK_c_704_n 0.0581908f $X=0.925 $Y=2.4 $X2=1.42
+ $Y2=2.275
cc_408 N_A_N233_612#_c_480_n N_CK_c_704_n 4.5169e-19 $X=0.925 $Y=2.4 $X2=1.42
+ $Y2=2.275
cc_409 N_A_N233_612#_c_475_n N_CK_c_713_n 0.00287606f $X=0.925 $Y=2.4 $X2=1.885
+ $Y2=2.575
cc_410 N_A_N233_612#_c_477_n N_A_43_110#_c_907_n 9.77657e-19 $X=-0.609 $Y=0.8
+ $X2=0.225 $Y2=2.195
cc_411 N_A_N233_612#_c_484_n N_A_43_110#_c_907_n 0.020887f $X=0.78 $Y=2.565
+ $X2=0.225 $Y2=2.195
cc_412 N_A_N233_612#_c_485_n N_A_43_110#_c_907_n 0.00241421f $X=-0.609 $Y=1.455
+ $X2=0.225 $Y2=2.195
cc_413 N_A_N233_612#_c_477_n N_A_43_110#_c_914_n 7.79024e-19 $X=-0.609 $Y=0.8
+ $X2=0.34 $Y2=1.37
cc_414 N_A_N233_612#_c_485_n N_A_43_110#_c_914_n 0.00130395f $X=-0.609 $Y=1.455
+ $X2=0.34 $Y2=1.37
cc_415 N_A_N233_612#_c_484_n N_A_43_110#_c_918_n 0.0259204f $X=0.78 $Y=2.565
+ $X2=0.37 $Y2=2.195
cc_416 N_A_N233_612#_M1002_g N_A_43_110#_c_919_n 0.00314369f $X=0.985 $Y=1.05
+ $X2=2.22 $Y2=2.195
cc_417 N_A_N233_612#_c_475_n N_A_43_110#_c_919_n 0.00237496f $X=0.925 $Y=2.4
+ $X2=2.22 $Y2=2.195
cc_418 N_A_N233_612#_c_480_n N_A_43_110#_c_919_n 0.00482511f $X=0.925 $Y=2.4
+ $X2=2.22 $Y2=2.195
cc_419 N_A_N233_612#_c_484_n N_A_43_110#_c_919_n 0.0610643f $X=0.78 $Y=2.565
+ $X2=2.22 $Y2=2.195
cc_420 N_A_254_515#_c_575_n N_CK_M1025_g 0.0122005f $X=1.885 $Y=1.825 $X2=1.345
+ $Y2=1.05
cc_421 N_A_254_515#_c_576_n N_CK_M1025_g 0.0256778f $X=1.885 $Y=1.66 $X2=1.345
+ $Y2=1.05
cc_422 N_A_254_515#_c_579_n N_CK_M1025_g 0.00936286f $X=1.485 $Y=2.655 $X2=1.345
+ $Y2=1.05
cc_423 N_A_254_515#_c_582_n N_CK_M1025_g 0.00439496f $X=1.57 $Y=1.825 $X2=1.345
+ $Y2=1.05
cc_424 N_A_254_515#_c_575_n N_CK_c_703_n 0.0107061f $X=1.885 $Y=1.825 $X2=1.75
+ $Y2=2.275
cc_425 N_A_254_515#_c_579_n N_CK_c_703_n 0.00994433f $X=1.485 $Y=2.655 $X2=1.75
+ $Y2=2.275
cc_426 N_A_254_515#_c_580_n N_CK_c_703_n 0.00524719f $X=2.865 $Y=1.825 $X2=1.75
+ $Y2=2.275
cc_427 N_A_254_515#_c_574_n N_CK_c_704_n 0.0174061f $X=1.405 $Y=2.74 $X2=1.42
+ $Y2=2.275
cc_428 N_A_254_515#_c_579_n N_CK_c_704_n 0.00254254f $X=1.485 $Y=2.655 $X2=1.42
+ $Y2=2.275
cc_429 N_A_254_515#_c_588_n N_CK_c_704_n 9.11794e-19 $X=1.485 $Y=2.74 $X2=1.42
+ $Y2=2.275
cc_430 N_A_254_515#_M1023_g N_CK_M1012_g 0.0612056f $X=1.345 $Y=4.56 $X2=1.945
+ $Y2=4.56
cc_431 N_A_254_515#_c_587_n N_CK_c_705_n 0.00342393f $X=3.22 $Y=3.075 $X2=2.735
+ $Y2=2.905
cc_432 N_A_254_515#_c_590_n N_CK_c_705_n 0.00191755f $X=3.22 $Y=2.195 $X2=2.735
+ $Y2=2.905
cc_433 N_A_254_515#_c_599_n N_CK_c_705_n 0.00260941f $X=3.22 $Y=3.16 $X2=2.735
+ $Y2=2.905
cc_434 N_A_254_515#_c_587_n N_CK_M1006_g 0.00491946f $X=3.22 $Y=3.075 $X2=2.735
+ $Y2=4.56
cc_435 N_A_254_515#_c_580_n N_CK_c_706_n 0.00620802f $X=2.865 $Y=1.825 $X2=2.79
+ $Y2=2.575
cc_436 N_A_254_515#_c_586_n N_CK_c_706_n 0.00735406f $X=2.95 $Y=2.11 $X2=2.79
+ $Y2=2.575
cc_437 N_A_254_515#_c_587_n N_CK_c_706_n 0.00575356f $X=3.22 $Y=3.075 $X2=2.79
+ $Y2=2.575
cc_438 N_A_254_515#_c_589_n N_CK_c_706_n 0.0020984f $X=2.95 $Y=1.825 $X2=2.79
+ $Y2=2.575
cc_439 N_A_254_515#_c_590_n N_CK_c_706_n 0.00257368f $X=3.22 $Y=2.195 $X2=2.79
+ $Y2=2.575
cc_440 N_A_254_515#_c_574_n N_CK_c_712_n 0.0213338f $X=1.405 $Y=2.74 $X2=1.885
+ $Y2=2.74
cc_441 N_A_254_515#_c_575_n N_CK_c_712_n 0.00224211f $X=1.885 $Y=1.825 $X2=1.885
+ $Y2=2.74
cc_442 N_A_254_515#_c_580_n N_CK_c_712_n 2.46382e-19 $X=2.865 $Y=1.825 $X2=1.885
+ $Y2=2.74
cc_443 N_A_254_515#_c_588_n N_CK_c_712_n 0.00102234f $X=1.485 $Y=2.74 $X2=1.885
+ $Y2=2.74
cc_444 N_A_254_515#_c_579_n N_CK_c_713_n 0.00426729f $X=1.485 $Y=2.655 $X2=1.885
+ $Y2=2.575
cc_445 N_A_254_515#_c_583_n N_CK_c_714_n 0.00862611f $X=2.95 $Y=0.8 $X2=2.762
+ $Y2=1.64
cc_446 N_A_254_515#_c_580_n N_CK_c_718_n 0.0111082f $X=2.865 $Y=1.825 $X2=2.762
+ $Y2=1.79
cc_447 N_A_254_515#_c_583_n N_CK_c_718_n 0.00425384f $X=2.95 $Y=0.8 $X2=2.762
+ $Y2=1.79
cc_448 N_A_254_515#_c_589_n N_CK_c_718_n 8.71368e-19 $X=2.95 $Y=1.825 $X2=2.762
+ $Y2=1.79
cc_449 N_A_254_515#_c_574_n N_CK_c_720_n 8.47686e-19 $X=1.405 $Y=2.74 $X2=1.885
+ $Y2=2.565
cc_450 N_A_254_515#_c_575_n N_CK_c_720_n 8.65047e-19 $X=1.885 $Y=1.825 $X2=1.885
+ $Y2=2.565
cc_451 N_A_254_515#_c_579_n N_CK_c_720_n 0.00783596f $X=1.485 $Y=2.655 $X2=1.885
+ $Y2=2.565
cc_452 N_A_254_515#_c_580_n N_CK_c_720_n 0.00210861f $X=2.865 $Y=1.825 $X2=1.885
+ $Y2=2.565
cc_453 N_A_254_515#_c_588_n N_CK_c_720_n 0.00985033f $X=1.485 $Y=2.74 $X2=1.885
+ $Y2=2.565
cc_454 N_A_254_515#_c_580_n N_CK_c_721_n 7.67725e-19 $X=2.865 $Y=1.825 $X2=2.88
+ $Y2=2.565
cc_455 N_A_254_515#_c_587_n N_CK_c_721_n 0.0294301f $X=3.22 $Y=3.075 $X2=2.88
+ $Y2=2.565
cc_456 N_A_254_515#_c_590_n N_CK_c_721_n 0.00560985f $X=3.22 $Y=2.195 $X2=2.88
+ $Y2=2.565
cc_457 N_A_254_515#_c_599_n N_CK_c_721_n 0.00706443f $X=3.22 $Y=3.16 $X2=2.88
+ $Y2=2.565
cc_458 N_A_254_515#_c_579_n N_CK_c_724_n 0.00742331f $X=1.485 $Y=2.655 $X2=2.03
+ $Y2=2.565
cc_459 N_A_254_515#_c_588_n N_CK_c_724_n 7.22629e-19 $X=1.485 $Y=2.74 $X2=2.03
+ $Y2=2.565
cc_460 N_A_254_515#_c_587_n N_CK_c_725_n 0.0154529f $X=3.22 $Y=3.075 $X2=5.485
+ $Y2=2.565
cc_461 N_A_254_515#_c_590_n N_CK_c_725_n 0.00297742f $X=3.22 $Y=2.195 $X2=5.485
+ $Y2=2.565
cc_462 N_A_254_515#_c_599_n N_CK_c_725_n 0.00442383f $X=3.22 $Y=3.16 $X2=5.485
+ $Y2=2.565
cc_463 N_A_254_515#_c_587_n N_CK_c_726_n 0.00247429f $X=3.22 $Y=3.075 $X2=3.025
+ $Y2=2.565
cc_464 N_A_254_515#_c_590_n N_CK_c_726_n 0.00227637f $X=3.22 $Y=2.195 $X2=3.025
+ $Y2=2.565
cc_465 N_A_254_515#_c_599_n N_CK_c_726_n 0.00259785f $X=3.22 $Y=3.16 $X2=3.025
+ $Y2=2.565
cc_466 N_A_254_515#_c_576_n N_A_43_110#_M1005_g 0.0962312f $X=1.885 $Y=1.66
+ $X2=2.305 $Y2=1.05
cc_467 N_A_254_515#_c_579_n N_A_43_110#_M1005_g 0.00249296f $X=1.485 $Y=2.655
+ $X2=2.305 $Y2=1.05
cc_468 N_A_254_515#_c_580_n N_A_43_110#_M1005_g 0.0148268f $X=2.865 $Y=1.825
+ $X2=2.305 $Y2=1.05
cc_469 N_A_254_515#_c_579_n N_A_43_110#_c_897_n 6.23191e-19 $X=1.485 $Y=2.655
+ $X2=2.365 $Y2=2.195
cc_470 N_A_254_515#_c_580_n N_A_43_110#_c_897_n 0.00290043f $X=2.865 $Y=1.825
+ $X2=2.365 $Y2=2.195
cc_471 N_A_254_515#_c_590_n N_A_43_110#_c_897_n 2.7472e-19 $X=3.22 $Y=2.195
+ $X2=2.365 $Y2=2.195
cc_472 N_A_254_515#_c_586_n N_A_43_110#_c_898_n 0.00129872f $X=2.95 $Y=2.11
+ $X2=3.66 $Y2=2.195
cc_473 N_A_254_515#_c_587_n N_A_43_110#_c_898_n 0.00182884f $X=3.22 $Y=3.075
+ $X2=3.66 $Y2=2.195
cc_474 N_A_254_515#_c_590_n N_A_43_110#_c_898_n 6.13768e-19 $X=3.22 $Y=2.195
+ $X2=3.66 $Y2=2.195
cc_475 N_A_254_515#_c_586_n N_A_43_110#_c_899_n 0.00256885f $X=2.95 $Y=2.11
+ $X2=3.662 $Y2=2.03
cc_476 N_A_254_515#_c_589_n N_A_43_110#_c_904_n 8.70096e-19 $X=2.95 $Y=1.825
+ $X2=3.75 $Y2=1.775
cc_477 N_A_254_515#_c_587_n N_A_43_110#_c_905_n 0.00709308f $X=3.22 $Y=3.075
+ $X2=3.75 $Y2=2.83
cc_478 N_A_254_515#_c_579_n N_A_43_110#_c_912_n 0.00297176f $X=1.485 $Y=2.655
+ $X2=2.365 $Y2=2.195
cc_479 N_A_254_515#_c_580_n N_A_43_110#_c_912_n 0.0171514f $X=2.865 $Y=1.825
+ $X2=2.365 $Y2=2.195
cc_480 N_A_254_515#_c_590_n N_A_43_110#_c_912_n 0.00582063f $X=3.22 $Y=2.195
+ $X2=2.365 $Y2=2.195
cc_481 N_A_254_515#_c_590_n N_A_43_110#_c_913_n 0.0111568f $X=3.22 $Y=2.195
+ $X2=3.66 $Y2=2.195
cc_482 N_A_254_515#_c_580_n N_A_43_110#_c_916_n 0.0127136f $X=2.865 $Y=1.825
+ $X2=3.515 $Y2=2.195
cc_483 N_A_254_515#_c_586_n N_A_43_110#_c_916_n 0.00365521f $X=2.95 $Y=2.11
+ $X2=3.515 $Y2=2.195
cc_484 N_A_254_515#_c_587_n N_A_43_110#_c_916_n 6.65649e-19 $X=3.22 $Y=3.075
+ $X2=3.515 $Y2=2.195
cc_485 N_A_254_515#_c_590_n N_A_43_110#_c_916_n 0.0264739f $X=3.22 $Y=2.195
+ $X2=3.515 $Y2=2.195
cc_486 N_A_254_515#_c_580_n N_A_43_110#_c_917_n 0.00713297f $X=2.865 $Y=1.825
+ $X2=2.515 $Y2=2.195
cc_487 N_A_254_515#_c_586_n N_A_43_110#_c_917_n 0.00124859f $X=2.95 $Y=2.11
+ $X2=2.515 $Y2=2.195
cc_488 N_A_254_515#_c_574_n N_A_43_110#_c_919_n 7.03361e-19 $X=1.405 $Y=2.74
+ $X2=2.22 $Y2=2.195
cc_489 N_A_254_515#_c_575_n N_A_43_110#_c_919_n 0.00411095f $X=1.885 $Y=1.825
+ $X2=2.22 $Y2=2.195
cc_490 N_A_254_515#_c_579_n N_A_43_110#_c_919_n 0.0156918f $X=1.485 $Y=2.655
+ $X2=2.22 $Y2=2.195
cc_491 N_A_254_515#_c_580_n N_A_43_110#_c_919_n 0.0253127f $X=2.865 $Y=1.825
+ $X2=2.22 $Y2=2.195
cc_492 N_A_254_515#_c_588_n N_A_43_110#_c_919_n 0.00531735f $X=1.485 $Y=2.74
+ $X2=2.22 $Y2=2.195
cc_493 N_A_254_515#_c_586_n N_A_43_110#_c_920_n 0.00108733f $X=2.95 $Y=2.11
+ $X2=3.66 $Y2=2.195
cc_494 N_A_254_515#_c_587_n N_A_43_110#_c_920_n 0.0014067f $X=3.22 $Y=3.075
+ $X2=3.66 $Y2=2.195
cc_495 N_A_254_515#_c_590_n N_A_43_110#_c_920_n 2.14718e-19 $X=3.22 $Y=2.195
+ $X2=3.66 $Y2=2.195
cc_496 N_A_254_515#_c_583_n N_A_687_110#_c_1078_n 0.0433959f $X=2.95 $Y=0.8
+ $X2=3.56 $Y2=0.8
cc_497 N_A_254_515#_c_595_n N_A_687_110#_c_1081_n 0.101394f $X=2.95 $Y=3.43
+ $X2=3.56 $Y2=2.935
cc_498 N_A_254_515#_c_587_n N_A_687_110#_c_1081_n 0.0163571f $X=3.22 $Y=3.075
+ $X2=3.56 $Y2=2.935
cc_499 N_A_254_515#_c_599_n N_A_687_110#_c_1081_n 0.0134687f $X=3.22 $Y=3.16
+ $X2=3.56 $Y2=2.935
cc_500 N_A_254_515#_c_589_n N_A_687_110#_c_1084_n 0.00821298f $X=2.95 $Y=1.825
+ $X2=3.645 $Y2=1.825
cc_501 N_A_254_515#_c_587_n N_A_687_110#_c_1086_n 0.0141728f $X=3.22 $Y=3.075
+ $X2=3.645 $Y2=2.74
cc_502 N_A_254_515#_c_587_n N_A_687_110#_c_1090_n 0.00864908f $X=3.22 $Y=3.075
+ $X2=3.705 $Y2=2.935
cc_503 N_CK_c_706_n N_A_43_110#_M1005_g 0.00882748f $X=2.79 $Y=2.575 $X2=2.305
+ $Y2=1.05
cc_504 N_CK_c_714_n N_A_43_110#_M1005_g 0.026973f $X=2.762 $Y=1.64 $X2=2.305
+ $Y2=1.05
cc_505 N_CK_c_705_n N_A_43_110#_M1004_g 0.0287701f $X=2.735 $Y=2.905 $X2=2.305
+ $Y2=4.56
cc_506 N_CK_c_706_n N_A_43_110#_M1004_g 0.0162964f $X=2.79 $Y=2.575 $X2=2.305
+ $Y2=4.56
cc_507 N_CK_c_712_n N_A_43_110#_M1004_g 0.214863f $X=1.885 $Y=2.74 $X2=2.305
+ $Y2=4.56
cc_508 N_CK_c_713_n N_A_43_110#_M1004_g 0.00761683f $X=1.885 $Y=2.575 $X2=2.305
+ $Y2=4.56
cc_509 N_CK_c_720_n N_A_43_110#_M1004_g 0.00367682f $X=1.885 $Y=2.565 $X2=2.305
+ $Y2=4.56
cc_510 N_CK_c_721_n N_A_43_110#_M1004_g 0.0026346f $X=2.88 $Y=2.565 $X2=2.305
+ $Y2=4.56
cc_511 N_CK_c_723_n N_A_43_110#_M1004_g 0.0105882f $X=2.735 $Y=2.565 $X2=2.305
+ $Y2=4.56
cc_512 N_CK_c_724_n N_A_43_110#_M1004_g 8.90723e-19 $X=2.03 $Y=2.565 $X2=2.305
+ $Y2=4.56
cc_513 N_CK_c_726_n N_A_43_110#_M1004_g 3.05655e-19 $X=3.025 $Y=2.565 $X2=2.305
+ $Y2=4.56
cc_514 N_CK_c_703_n N_A_43_110#_c_897_n 0.00761683f $X=1.75 $Y=2.275 $X2=2.365
+ $Y2=2.195
cc_515 N_CK_c_706_n N_A_43_110#_c_897_n 0.02116f $X=2.79 $Y=2.575 $X2=2.365
+ $Y2=2.195
cc_516 N_CK_c_723_n N_A_43_110#_c_897_n 0.00186852f $X=2.735 $Y=2.565 $X2=2.365
+ $Y2=2.195
cc_517 N_CK_c_706_n N_A_43_110#_c_898_n 0.00376174f $X=2.79 $Y=2.575 $X2=3.66
+ $Y2=2.195
cc_518 N_CK_c_725_n N_A_43_110#_c_898_n 0.00194637f $X=5.485 $Y=2.565 $X2=3.66
+ $Y2=2.195
cc_519 N_CK_c_705_n N_A_43_110#_c_905_n 0.00460238f $X=2.735 $Y=2.905 $X2=3.75
+ $Y2=2.83
cc_520 N_CK_c_725_n N_A_43_110#_c_905_n 0.00644656f $X=5.485 $Y=2.565 $X2=3.75
+ $Y2=2.83
cc_521 N_CK_c_703_n N_A_43_110#_c_912_n 6.64388e-19 $X=1.75 $Y=2.275 $X2=2.365
+ $Y2=2.195
cc_522 N_CK_c_706_n N_A_43_110#_c_912_n 9.45138e-19 $X=2.79 $Y=2.575 $X2=2.365
+ $Y2=2.195
cc_523 N_CK_c_723_n N_A_43_110#_c_912_n 0.00487271f $X=2.735 $Y=2.565 $X2=2.365
+ $Y2=2.195
cc_524 N_CK_c_706_n N_A_43_110#_c_913_n 2.20146e-19 $X=2.79 $Y=2.575 $X2=3.66
+ $Y2=2.195
cc_525 N_CK_c_725_n N_A_43_110#_c_913_n 0.00227722f $X=5.485 $Y=2.565 $X2=3.66
+ $Y2=2.195
cc_526 N_CK_c_706_n N_A_43_110#_c_916_n 0.00359701f $X=2.79 $Y=2.575 $X2=3.515
+ $Y2=2.195
cc_527 N_CK_c_721_n N_A_43_110#_c_916_n 5.86675e-19 $X=2.88 $Y=2.565 $X2=3.515
+ $Y2=2.195
cc_528 N_CK_c_723_n N_A_43_110#_c_916_n 0.0178163f $X=2.735 $Y=2.565 $X2=3.515
+ $Y2=2.195
cc_529 N_CK_c_725_n N_A_43_110#_c_916_n 0.0377042f $X=5.485 $Y=2.565 $X2=3.515
+ $Y2=2.195
cc_530 N_CK_c_726_n N_A_43_110#_c_916_n 0.0247363f $X=3.025 $Y=2.565 $X2=3.515
+ $Y2=2.195
cc_531 N_CK_c_703_n N_A_43_110#_c_917_n 4.70316e-19 $X=1.75 $Y=2.275 $X2=2.515
+ $Y2=2.195
cc_532 N_CK_c_706_n N_A_43_110#_c_917_n 9.27087e-19 $X=2.79 $Y=2.575 $X2=2.515
+ $Y2=2.195
cc_533 N_CK_c_723_n N_A_43_110#_c_917_n 0.0270759f $X=2.735 $Y=2.565 $X2=2.515
+ $Y2=2.195
cc_534 N_CK_M1025_g N_A_43_110#_c_919_n 0.00255623f $X=1.345 $Y=1.05 $X2=2.22
+ $Y2=2.195
cc_535 N_CK_c_703_n N_A_43_110#_c_919_n 0.00985983f $X=1.75 $Y=2.275 $X2=2.22
+ $Y2=2.195
cc_536 N_CK_c_704_n N_A_43_110#_c_919_n 0.00164908f $X=1.42 $Y=2.275 $X2=2.22
+ $Y2=2.195
cc_537 N_CK_c_720_n N_A_43_110#_c_919_n 9.69764e-19 $X=1.885 $Y=2.565 $X2=2.22
+ $Y2=2.195
cc_538 N_CK_c_723_n N_A_43_110#_c_919_n 0.0147541f $X=2.735 $Y=2.565 $X2=2.22
+ $Y2=2.195
cc_539 N_CK_c_724_n N_A_43_110#_c_919_n 0.0242903f $X=2.03 $Y=2.565 $X2=2.22
+ $Y2=2.195
cc_540 N_CK_c_725_n N_A_43_110#_c_920_n 0.0265966f $X=5.485 $Y=2.565 $X2=3.66
+ $Y2=2.195
cc_541 N_CK_c_725_n N_A_687_110#_M1008_g 0.00440546f $X=5.485 $Y=2.565 $X2=4.205
+ $Y2=4.56
cc_542 N_CK_M1021_g N_A_687_110#_M1018_g 0.0402111f $X=5.585 $Y=1.05 $X2=5.155
+ $Y2=1.05
cc_543 N_CK_c_719_n N_A_687_110#_M1018_g 0.0153344f $X=5.63 $Y=2.36 $X2=5.155
+ $Y2=1.05
cc_544 N_CK_c_722_n N_A_687_110#_M1018_g 0.00130485f $X=5.63 $Y=2.36 $X2=5.155
+ $Y2=1.05
cc_545 N_CK_c_725_n N_A_687_110#_M1018_g 0.00527112f $X=5.485 $Y=2.565 $X2=5.155
+ $Y2=1.05
cc_546 N_CK_c_725_n N_A_687_110#_c_1076_n 0.00130191f $X=5.485 $Y=2.565
+ $X2=4.145 $Y2=2.195
cc_547 N_CK_M1020_g N_A_687_110#_c_1077_n 0.155966f $X=5.585 $Y=4.56 $X2=5.155
+ $Y2=2.65
cc_548 N_CK_c_725_n N_A_687_110#_c_1077_n 0.00552994f $X=5.485 $Y=2.565
+ $X2=5.155 $Y2=2.65
cc_549 N_CK_M1006_g N_A_687_110#_c_1081_n 0.0063972f $X=2.735 $Y=4.56 $X2=3.56
+ $Y2=2.935
cc_550 N_CK_c_725_n N_A_687_110#_c_1082_n 0.00746701f $X=5.485 $Y=2.565 $X2=4.06
+ $Y2=1.825
cc_551 N_CK_c_718_n N_A_687_110#_c_1084_n 8.76784e-19 $X=2.762 $Y=1.79 $X2=3.645
+ $Y2=1.825
cc_552 N_CK_c_725_n N_A_687_110#_c_1085_n 0.00951711f $X=5.485 $Y=2.565 $X2=4.06
+ $Y2=2.74
cc_553 N_CK_c_725_n N_A_687_110#_c_1086_n 0.00301504f $X=5.485 $Y=2.565
+ $X2=3.645 $Y2=2.74
cc_554 N_CK_c_725_n N_A_687_110#_c_1087_n 0.0197525f $X=5.485 $Y=2.565 $X2=4.145
+ $Y2=2.195
cc_555 N_CK_c_725_n N_A_687_110#_c_1088_n 0.0117944f $X=5.485 $Y=2.565 $X2=4.95
+ $Y2=2.65
cc_556 N_CK_c_725_n N_A_687_110#_c_1089_n 0.125093f $X=5.485 $Y=2.565 $X2=4.805
+ $Y2=2.935
cc_557 N_CK_c_725_n N_A_687_110#_c_1090_n 0.0350814f $X=5.485 $Y=2.565 $X2=3.705
+ $Y2=2.935
cc_558 N_CK_M1021_g N_A_963_612#_M1013_g 0.030724f $X=5.585 $Y=1.05 $X2=6.015
+ $Y2=1.05
cc_559 N_CK_M1021_g N_A_963_612#_c_1191_n 0.0119161f $X=5.585 $Y=1.05 $X2=6.05
+ $Y2=2.075
cc_560 N_CK_M1020_g N_A_963_612#_c_1192_n 0.00914307f $X=5.585 $Y=4.56 $X2=6.032
+ $Y2=2.785
cc_561 N_CK_c_719_n N_A_963_612#_c_1192_n 0.0206139f $X=5.63 $Y=2.36 $X2=6.032
+ $Y2=2.785
cc_562 N_CK_c_722_n N_A_963_612#_c_1192_n 0.00374476f $X=5.63 $Y=2.36 $X2=6.032
+ $Y2=2.785
cc_563 N_CK_c_727_n N_A_963_612#_c_1192_n 0.00124193f $X=5.63 $Y=2.565 $X2=6.032
+ $Y2=2.785
cc_564 N_CK_M1020_g N_A_963_612#_c_1193_n 0.0540618f $X=5.585 $Y=4.56 $X2=6.032
+ $Y2=2.935
cc_565 N_CK_c_722_n N_A_963_612#_c_1193_n 0.00341181f $X=5.63 $Y=2.36 $X2=6.032
+ $Y2=2.935
cc_566 N_CK_c_744_n N_A_963_612#_c_1193_n 0.00374181f $X=5.63 $Y=2.565 $X2=6.032
+ $Y2=2.935
cc_567 N_CK_M1020_g N_A_963_612#_c_1218_n 0.00457566f $X=5.585 $Y=4.56 $X2=5.205
+ $Y2=3.605
cc_568 N_CK_M1021_g N_A_963_612#_c_1194_n 0.00429604f $X=5.585 $Y=1.05 $X2=5.29
+ $Y2=3.52
cc_569 N_CK_M1020_g N_A_963_612#_c_1194_n 0.00760546f $X=5.585 $Y=4.56 $X2=5.29
+ $Y2=3.52
cc_570 N_CK_c_719_n N_A_963_612#_c_1194_n 0.00203726f $X=5.63 $Y=2.36 $X2=5.29
+ $Y2=3.52
cc_571 N_CK_c_722_n N_A_963_612#_c_1194_n 0.0810452f $X=5.63 $Y=2.36 $X2=5.29
+ $Y2=3.52
cc_572 N_CK_c_744_n N_A_963_612#_c_1194_n 0.00866797f $X=5.63 $Y=2.565 $X2=5.29
+ $Y2=3.52
cc_573 N_CK_c_725_n N_A_963_612#_c_1194_n 0.0246701f $X=5.485 $Y=2.565 $X2=5.29
+ $Y2=3.52
cc_574 N_CK_c_727_n N_A_963_612#_c_1194_n 0.00183606f $X=5.63 $Y=2.565 $X2=5.29
+ $Y2=3.52
cc_575 N_CK_M1021_g N_A_963_612#_c_1195_n 0.00765999f $X=5.585 $Y=1.05 $X2=5.37
+ $Y2=0.8
cc_576 N_CK_M1021_g N_A_963_612#_c_1198_n 0.0154849f $X=5.585 $Y=1.05 $X2=6.11
+ $Y2=1.91
cc_577 N_CK_c_719_n N_A_963_612#_c_1198_n 0.00276813f $X=5.63 $Y=2.36 $X2=6.11
+ $Y2=1.91
cc_578 N_CK_c_722_n N_A_963_612#_c_1198_n 0.0108125f $X=5.63 $Y=2.36 $X2=6.11
+ $Y2=1.91
cc_579 N_CK_c_725_n N_A_963_612#_c_1198_n 9.91959e-19 $X=5.485 $Y=2.565 $X2=6.11
+ $Y2=1.91
cc_580 N_CK_c_727_n N_A_963_612#_c_1198_n 0.00461695f $X=5.63 $Y=2.565 $X2=6.11
+ $Y2=1.91
cc_581 N_CK_c_725_n N_A_963_612#_c_1200_n 0.00316638f $X=5.485 $Y=2.565 $X2=5.33
+ $Y2=1.91
cc_582 N_CK_c_725_n N_A_856_110#_c_1274_n 0.0193167f $X=5.485 $Y=2.565 $X2=4.452
+ $Y2=3.135
cc_583 N_CK_c_744_n A_1046_612# 0.0116178f $X=5.63 $Y=2.565 $X2=5.23 $Y2=3.06
cc_584 N_CK_c_722_n N_ECK_c_1307_n 0.0215696f $X=5.63 $Y=2.36 $X2=6.23 $Y2=2.565
cc_585 N_CK_c_744_n N_ECK_c_1307_n 0.00659455f $X=5.63 $Y=2.565 $X2=6.23
+ $Y2=2.565
cc_586 N_CK_c_727_n N_ECK_c_1307_n 0.00103949f $X=5.63 $Y=2.565 $X2=6.23
+ $Y2=2.565
cc_587 N_CK_M1021_g N_ECK_c_1308_n 6.73508e-19 $X=5.585 $Y=1.05 $X2=6.23
+ $Y2=2.45
cc_588 N_CK_c_722_n N_ECK_c_1308_n 0.00825539f $X=5.63 $Y=2.36 $X2=6.23 $Y2=2.45
cc_589 N_CK_M1021_g N_ECK_c_1309_n 7.99941e-19 $X=5.585 $Y=1.05 $X2=6.23
+ $Y2=1.455
cc_590 N_CK_c_722_n ECK 0.0012208f $X=5.63 $Y=2.36 $X2=6.23 $Y2=2.565
cc_591 N_CK_c_727_n ECK 0.0172304f $X=5.63 $Y=2.565 $X2=6.23 $Y2=2.565
cc_592 N_A_43_110#_c_899_n N_A_687_110#_M1009_g 0.00883234f $X=3.662 $Y=2.03
+ $X2=4.205 $Y2=1.05
cc_593 N_A_43_110#_c_900_n N_A_687_110#_M1009_g 0.0248201f $X=3.75 $Y=1.625
+ $X2=4.205 $Y2=1.05
cc_594 N_A_43_110#_c_905_n N_A_687_110#_M1008_g 0.0170958f $X=3.75 $Y=2.83
+ $X2=4.205 $Y2=4.56
cc_595 N_A_43_110#_c_906_n N_A_687_110#_M1008_g 0.0245862f $X=3.75 $Y=2.98
+ $X2=4.205 $Y2=4.56
cc_596 N_A_43_110#_c_898_n N_A_687_110#_c_1076_n 0.0213149f $X=3.66 $Y=2.195
+ $X2=4.145 $Y2=2.195
cc_597 N_A_43_110#_c_913_n N_A_687_110#_c_1076_n 0.00104076f $X=3.66 $Y=2.195
+ $X2=4.145 $Y2=2.195
cc_598 N_A_43_110#_c_920_n N_A_687_110#_c_1076_n 9.12123e-19 $X=3.66 $Y=2.195
+ $X2=4.145 $Y2=2.195
cc_599 N_A_43_110#_c_900_n N_A_687_110#_c_1078_n 0.00804393f $X=3.75 $Y=1.625
+ $X2=3.56 $Y2=0.8
cc_600 N_A_43_110#_c_904_n N_A_687_110#_c_1078_n 0.00485394f $X=3.75 $Y=1.775
+ $X2=3.56 $Y2=0.8
cc_601 N_A_43_110#_c_905_n N_A_687_110#_c_1081_n 0.00486816f $X=3.75 $Y=2.83
+ $X2=3.56 $Y2=2.935
cc_602 N_A_43_110#_c_906_n N_A_687_110#_c_1081_n 0.00708078f $X=3.75 $Y=2.98
+ $X2=3.56 $Y2=2.935
cc_603 N_A_43_110#_c_899_n N_A_687_110#_c_1082_n 0.00816842f $X=3.662 $Y=2.03
+ $X2=4.06 $Y2=1.825
cc_604 N_A_43_110#_c_904_n N_A_687_110#_c_1082_n 0.011031f $X=3.75 $Y=1.775
+ $X2=4.06 $Y2=1.825
cc_605 N_A_43_110#_c_913_n N_A_687_110#_c_1082_n 0.00924735f $X=3.66 $Y=2.195
+ $X2=4.06 $Y2=1.825
cc_606 N_A_43_110#_c_920_n N_A_687_110#_c_1082_n 0.0037949f $X=3.66 $Y=2.195
+ $X2=4.06 $Y2=1.825
cc_607 N_A_43_110#_c_898_n N_A_687_110#_c_1084_n 0.00303508f $X=3.66 $Y=2.195
+ $X2=3.645 $Y2=1.825
cc_608 N_A_43_110#_c_913_n N_A_687_110#_c_1084_n 0.00899348f $X=3.66 $Y=2.195
+ $X2=3.645 $Y2=1.825
cc_609 N_A_43_110#_c_916_n N_A_687_110#_c_1084_n 0.0011692f $X=3.515 $Y=2.195
+ $X2=3.645 $Y2=1.825
cc_610 N_A_43_110#_c_920_n N_A_687_110#_c_1084_n 0.00331526f $X=3.66 $Y=2.195
+ $X2=3.645 $Y2=1.825
cc_611 N_A_43_110#_c_905_n N_A_687_110#_c_1085_n 0.0122834f $X=3.75 $Y=2.83
+ $X2=4.06 $Y2=2.74
cc_612 N_A_43_110#_c_906_n N_A_687_110#_c_1085_n 0.00248624f $X=3.75 $Y=2.98
+ $X2=4.06 $Y2=2.74
cc_613 N_A_43_110#_c_913_n N_A_687_110#_c_1085_n 0.00388233f $X=3.66 $Y=2.195
+ $X2=4.06 $Y2=2.74
cc_614 N_A_43_110#_c_898_n N_A_687_110#_c_1086_n 0.00271474f $X=3.66 $Y=2.195
+ $X2=3.645 $Y2=2.74
cc_615 N_A_43_110#_c_913_n N_A_687_110#_c_1086_n 0.00388844f $X=3.66 $Y=2.195
+ $X2=3.645 $Y2=2.74
cc_616 N_A_43_110#_c_898_n N_A_687_110#_c_1087_n 0.00116148f $X=3.66 $Y=2.195
+ $X2=4.145 $Y2=2.195
cc_617 N_A_43_110#_c_899_n N_A_687_110#_c_1087_n 0.0022611f $X=3.662 $Y=2.03
+ $X2=4.145 $Y2=2.195
cc_618 N_A_43_110#_c_905_n N_A_687_110#_c_1087_n 0.00474984f $X=3.75 $Y=2.83
+ $X2=4.145 $Y2=2.195
cc_619 N_A_43_110#_c_913_n N_A_687_110#_c_1087_n 0.00887114f $X=3.66 $Y=2.195
+ $X2=4.145 $Y2=2.195
cc_620 N_A_43_110#_c_920_n N_A_687_110#_c_1087_n 0.0035858f $X=3.66 $Y=2.195
+ $X2=4.145 $Y2=2.195
cc_621 N_A_43_110#_c_906_n N_A_687_110#_c_1089_n 0.0083553f $X=3.75 $Y=2.98
+ $X2=4.805 $Y2=2.935
cc_622 N_A_43_110#_c_906_n N_A_687_110#_c_1090_n 0.00392333f $X=3.75 $Y=2.98
+ $X2=3.705 $Y2=2.935
cc_623 N_A_687_110#_M1016_g N_A_963_612#_c_1218_n 0.0140282f $X=5.155 $Y=4.56
+ $X2=5.205 $Y2=3.605
cc_624 N_A_687_110#_c_1089_n N_A_963_612#_c_1218_n 0.00520961f $X=4.805 $Y=2.935
+ $X2=5.205 $Y2=3.605
cc_625 N_A_687_110#_c_1088_n N_A_963_612#_c_1235_n 0.00369517f $X=4.95 $Y=2.65
+ $X2=5.025 $Y2=3.605
cc_626 N_A_687_110#_c_1089_n N_A_963_612#_c_1235_n 0.00431991f $X=4.805 $Y=2.935
+ $X2=5.025 $Y2=3.605
cc_627 N_A_687_110#_M1018_g N_A_963_612#_c_1194_n 0.0139576f $X=5.155 $Y=1.05
+ $X2=5.29 $Y2=3.52
cc_628 N_A_687_110#_M1016_g N_A_963_612#_c_1194_n 0.0219414f $X=5.155 $Y=4.56
+ $X2=5.29 $Y2=3.52
cc_629 N_A_687_110#_c_1077_n N_A_963_612#_c_1194_n 0.00663709f $X=5.155 $Y=2.65
+ $X2=5.29 $Y2=3.52
cc_630 N_A_687_110#_c_1088_n N_A_963_612#_c_1194_n 0.0344462f $X=4.95 $Y=2.65
+ $X2=5.29 $Y2=3.52
cc_631 N_A_687_110#_c_1089_n N_A_963_612#_c_1194_n 0.0078142f $X=4.805 $Y=2.935
+ $X2=5.29 $Y2=3.52
cc_632 N_A_687_110#_M1018_g N_A_963_612#_c_1195_n 0.00765999f $X=5.155 $Y=1.05
+ $X2=5.37 $Y2=0.8
cc_633 N_A_687_110#_M1018_g N_A_963_612#_c_1200_n 0.00698836f $X=5.155 $Y=1.05
+ $X2=5.33 $Y2=1.91
cc_634 N_A_687_110#_M1018_g N_A_856_110#_c_1269_n 0.00193244f $X=5.155 $Y=1.05
+ $X2=4.42 $Y2=0.8
cc_635 N_A_687_110#_M1008_g N_A_856_110#_c_1275_n 0.0120377f $X=4.205 $Y=4.56
+ $X2=4.42 $Y2=3.305
cc_636 N_A_687_110#_M1016_g N_A_856_110#_c_1275_n 0.00233754f $X=5.155 $Y=4.56
+ $X2=4.42 $Y2=3.305
cc_637 N_A_687_110#_c_1089_n N_A_856_110#_c_1275_n 0.0367582f $X=4.805 $Y=2.935
+ $X2=4.42 $Y2=3.305
cc_638 N_A_687_110#_M1016_g N_A_856_110#_c_1277_n 0.00474969f $X=5.155 $Y=4.56
+ $X2=4.42 $Y2=3.43
cc_639 N_A_687_110#_M1009_g N_A_856_110#_c_1273_n 0.00595737f $X=4.205 $Y=1.05
+ $X2=4.452 $Y2=1.57
cc_640 N_A_687_110#_M1018_g N_A_856_110#_c_1273_n 0.0206234f $X=5.155 $Y=1.05
+ $X2=4.452 $Y2=1.57
cc_641 N_A_687_110#_M1009_g N_A_856_110#_c_1274_n 0.0349327f $X=4.205 $Y=1.05
+ $X2=4.452 $Y2=3.135
cc_642 N_A_687_110#_M1016_g N_A_856_110#_c_1274_n 0.00464383f $X=5.155 $Y=4.56
+ $X2=4.452 $Y2=3.135
cc_643 N_A_687_110#_c_1077_n N_A_856_110#_c_1274_n 0.00266931f $X=5.155 $Y=2.65
+ $X2=4.452 $Y2=3.135
cc_644 N_A_687_110#_c_1082_n N_A_856_110#_c_1274_n 0.0135849f $X=4.06 $Y=1.825
+ $X2=4.452 $Y2=3.135
cc_645 N_A_687_110#_c_1085_n N_A_856_110#_c_1274_n 0.0135737f $X=4.06 $Y=2.74
+ $X2=4.452 $Y2=3.135
cc_646 N_A_687_110#_c_1087_n N_A_856_110#_c_1274_n 0.0520698f $X=4.145 $Y=2.195
+ $X2=4.452 $Y2=3.135
cc_647 N_A_687_110#_c_1088_n N_A_856_110#_c_1274_n 0.0224071f $X=4.95 $Y=2.65
+ $X2=4.452 $Y2=3.135
cc_648 N_A_687_110#_c_1089_n N_A_856_110#_c_1274_n 0.0184728f $X=4.805 $Y=2.935
+ $X2=4.452 $Y2=3.135
cc_649 N_A_963_612#_c_1205_n N_A_856_110#_c_1277_n 0.101221f $X=4.94 $Y=3.77
+ $X2=4.42 $Y2=3.43
cc_650 N_A_963_612#_c_1235_n N_A_856_110#_c_1277_n 0.0079413f $X=5.025 $Y=3.605
+ $X2=4.42 $Y2=3.43
cc_651 N_A_963_612#_c_1194_n N_A_856_110#_c_1274_n 0.0199414f $X=5.29 $Y=3.52
+ $X2=4.452 $Y2=3.135
cc_652 N_A_963_612#_c_1200_n N_A_856_110#_c_1274_n 0.00493879f $X=5.33 $Y=1.91
+ $X2=4.452 $Y2=3.135
cc_653 N_A_963_612#_c_1218_n A_1046_612# 0.00613297f $X=5.205 $Y=3.605 $X2=5.23
+ $Y2=3.06
cc_654 N_A_963_612#_c_1194_n A_1046_612# 0.00377193f $X=5.29 $Y=3.52 $X2=5.23
+ $Y2=3.06
cc_655 N_A_963_612#_M1013_g N_ECK_c_1304_n 0.0057847f $X=6.015 $Y=1.05 $X2=6.23
+ $Y2=0.8
cc_656 N_A_963_612#_c_1191_n N_ECK_c_1304_n 0.00168f $X=6.05 $Y=2.075 $X2=6.23
+ $Y2=0.8
cc_657 N_A_963_612#_c_1198_n N_ECK_c_1304_n 0.00510008f $X=6.11 $Y=1.91 $X2=6.23
+ $Y2=0.8
cc_658 N_A_963_612#_c_1191_n N_ECK_c_1307_n 0.00125776f $X=6.05 $Y=2.075
+ $X2=6.23 $Y2=2.565
cc_659 N_A_963_612#_c_1192_n N_ECK_c_1307_n 0.0115869f $X=6.032 $Y=2.785
+ $X2=6.23 $Y2=2.565
cc_660 N_A_963_612#_c_1193_n N_ECK_c_1307_n 0.00755607f $X=6.032 $Y=2.935
+ $X2=6.23 $Y2=2.565
cc_661 N_A_963_612#_c_1198_n N_ECK_c_1307_n 0.00273485f $X=6.11 $Y=1.91 $X2=6.23
+ $Y2=2.565
cc_662 N_A_963_612#_M1013_g N_ECK_c_1308_n 0.00406656f $X=6.015 $Y=1.05 $X2=6.23
+ $Y2=2.45
cc_663 N_A_963_612#_c_1191_n N_ECK_c_1308_n 0.00704613f $X=6.05 $Y=2.075
+ $X2=6.23 $Y2=2.45
cc_664 N_A_963_612#_c_1192_n N_ECK_c_1308_n 0.00892438f $X=6.032 $Y=2.785
+ $X2=6.23 $Y2=2.45
cc_665 N_A_963_612#_c_1198_n N_ECK_c_1308_n 0.0151477f $X=6.11 $Y=1.91 $X2=6.23
+ $Y2=2.45
cc_666 N_A_963_612#_M1013_g N_ECK_c_1309_n 0.00669813f $X=6.015 $Y=1.05 $X2=6.23
+ $Y2=1.455
cc_667 N_A_963_612#_c_1191_n N_ECK_c_1309_n 0.00154864f $X=6.05 $Y=2.075
+ $X2=6.23 $Y2=1.455
cc_668 N_A_963_612#_c_1198_n N_ECK_c_1309_n 0.00238892f $X=6.11 $Y=1.91 $X2=6.23
+ $Y2=1.455
cc_669 N_A_963_612#_c_1191_n ECK 4.58687e-19 $X=6.05 $Y=2.075 $X2=6.23 $Y2=2.565
cc_670 N_A_963_612#_c_1192_n ECK 0.00592444f $X=6.032 $Y=2.785 $X2=6.23
+ $Y2=2.565
cc_671 N_A_963_612#_c_1198_n ECK 0.00181779f $X=6.11 $Y=1.91 $X2=6.23 $Y2=2.565
