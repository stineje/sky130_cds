* File: sky130_osu_sc_12T_ms__dffnr_l.pxi.spice
* Created: Fri Feb 12 20:30:18 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%GND N_GND_M1021_s N_GND_M1018_s N_GND_M1005_d
+ N_GND_M1007_s N_GND_M1027_d N_GND_M1023_d N_GND_M1012_s N_GND_M1013_d
+ N_GND_M1016_d N_GND_M1021_b N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_12_p
+ N_GND_c_41_p N_GND_c_42_p N_GND_c_43_p N_GND_c_44_p N_GND_c_45_p N_GND_c_46_p
+ N_GND_c_47_p N_GND_c_48_p N_GND_c_49_p N_GND_c_19_p N_GND_c_16_p N_GND_c_175_p
+ N_GND_c_176_p GND N_GND_c_5_p PM_SKY130_OSU_SC_12T_MS__DFFNR_L%GND
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%VDD N_VDD_M1004_s N_VDD_M1002_d N_VDD_M1028_s
+ N_VDD_M1022_d N_VDD_M1009_d N_VDD_M1030_d N_VDD_M1011_d N_VDD_M1004_b
+ N_VDD_c_250_p N_VDD_c_251_p N_VDD_c_270_p N_VDD_c_274_p N_VDD_c_276_p
+ N_VDD_c_304_p N_VDD_c_291_p N_VDD_c_324_p N_VDD_c_262_p N_VDD_c_263_p
+ N_VDD_c_334_p N_VDD_c_335_p VDD N_VDD_c_252_p N_VDD_c_360_p
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%RN N_RN_M1021_g N_RN_c_383_n N_RN_M1004_g
+ N_RN_c_385_n N_RN_c_386_n RN PM_SKY130_OSU_SC_12T_MS__DFFNR_L%RN
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_110_115# N_A_110_115#_M1021_d
+ N_A_110_115#_M1004_d N_A_110_115#_c_416_n N_A_110_115#_M1018_g
+ N_A_110_115#_M1015_g N_A_110_115#_c_421_n N_A_110_115#_M1030_g
+ N_A_110_115#_c_424_n N_A_110_115#_M1013_g N_A_110_115#_c_428_n
+ N_A_110_115#_c_432_n N_A_110_115#_c_433_n N_A_110_115#_c_434_n
+ N_A_110_115#_c_436_n N_A_110_115#_c_437_n N_A_110_115#_c_536_p
+ N_A_110_115#_c_438_n N_A_110_115#_c_458_n N_A_110_115#_c_565_p
+ N_A_110_115#_c_462_n N_A_110_115#_c_463_n N_A_110_115#_c_464_n
+ N_A_110_115#_c_466_n N_A_110_115#_c_468_n
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_110_115#
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_342_442# N_A_342_442#_M1031_d
+ N_A_342_442#_M1024_d N_A_342_442#_M1002_g N_A_342_442#_M1005_g
+ N_A_342_442#_c_618_n N_A_342_442#_c_633_n N_A_342_442#_c_619_n
+ N_A_342_442#_c_621_n N_A_342_442#_c_623_n N_A_342_442#_c_636_n
+ N_A_342_442#_c_624_n N_A_342_442#_c_625_n N_A_342_442#_c_626_n
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_342_442#
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%D N_D_M1007_g N_D_M1028_g D N_D_c_703_n
+ N_D_c_704_n PM_SKY130_OSU_SC_12T_MS__DFFNR_L%D
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_618_424# N_A_618_424#_M1010_d
+ N_A_618_424#_M1029_d N_A_618_424#_M1024_g N_A_618_424#_M1026_g
+ N_A_618_424#_M1019_g N_A_618_424#_M1000_g N_A_618_424#_c_739_n
+ N_A_618_424#_c_740_n N_A_618_424#_c_741_n N_A_618_424#_c_742_n
+ N_A_618_424#_c_743_n N_A_618_424#_c_744_n N_A_618_424#_c_745_n
+ N_A_618_424#_c_776_n N_A_618_424#_c_746_n N_A_618_424#_c_779_n
+ N_A_618_424#_c_871_p N_A_618_424#_c_749_n N_A_618_424#_c_753_n
+ N_A_618_424#_c_754_n N_A_618_424#_c_755_n N_A_618_424#_c_756_n
+ N_A_618_424#_c_757_n N_A_618_424#_c_758_n N_A_618_424#_c_759_n
+ N_A_618_424#_c_760_n N_A_618_424#_c_761_n N_A_618_424#_c_762_n
+ N_A_618_424#_c_763_n N_A_618_424#_c_766_n N_A_618_424#_c_769_n
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_618_424#
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_217_605# N_A_217_605#_M1018_d
+ N_A_217_605#_M1015_s N_A_217_605#_M1027_g N_A_217_605#_M1022_g
+ N_A_217_605#_M1025_g N_A_217_605#_M1014_g N_A_217_605#_c_1005_n
+ N_A_217_605#_c_1006_n N_A_217_605#_c_1007_n N_A_217_605#_c_1009_n
+ N_A_217_605#_c_1010_n N_A_217_605#_c_1011_n N_A_217_605#_c_1012_n
+ N_A_217_605#_c_1013_n N_A_217_605#_c_1014_n N_A_217_605#_c_1015_n
+ N_A_217_605#_c_1061_n N_A_217_605#_c_1016_n N_A_217_605#_c_1018_n
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_217_605#
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%CK N_CK_c_1135_n N_CK_M1031_g N_CK_c_1138_n
+ N_CK_c_1139_n N_CK_c_1140_n N_CK_M1017_g N_CK_c_1142_n N_CK_M1003_g
+ N_CK_c_1144_n N_CK_M1020_g N_CK_c_1148_n N_CK_M1010_g N_CK_c_1153_n
+ N_CK_M1029_g N_CK_c_1154_n N_CK_c_1155_n N_CK_c_1156_n N_CK_c_1157_n
+ N_CK_c_1158_n N_CK_c_1159_n N_CK_c_1160_n N_CK_c_1246_n N_CK_c_1161_n CK
+ N_CK_c_1163_n N_CK_c_1164_n PM_SKY130_OSU_SC_12T_MS__DFFNR_L%CK
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_1160_89# N_A_1160_89#_M1012_d
+ N_A_1160_89#_M1006_s N_A_1160_89#_M1023_g N_A_1160_89#_M1009_g
+ N_A_1160_89#_M1016_g N_A_1160_89#_M1011_g N_A_1160_89#_c_1345_n
+ N_A_1160_89#_c_1349_n N_A_1160_89#_c_1350_n N_A_1160_89#_c_1351_n
+ N_A_1160_89#_c_1352_n N_A_1160_89#_c_1353_n N_A_1160_89#_c_1354_n
+ N_A_1160_89#_c_1385_n N_A_1160_89#_c_1388_n N_A_1160_89#_c_1389_n
+ N_A_1160_89#_c_1355_n N_A_1160_89#_c_1358_n N_A_1160_89#_c_1359_n
+ N_A_1160_89#_c_1361_n N_A_1160_89#_c_1363_n N_A_1160_89#_c_1364_n
+ N_A_1160_89#_c_1365_n N_A_1160_89#_c_1366_n N_A_1160_89#_c_1367_n
+ N_A_1160_89#_c_1368_n N_A_1160_89#_c_1369_n N_A_1160_89#_c_1370_n
+ N_A_1160_89#_c_1371_n N_A_1160_89#_c_1372_n N_A_1160_89#_c_1373_n
+ N_A_1160_89#_c_1374_n PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_1160_89#
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_998_115# N_A_998_115#_M1019_d
+ N_A_998_115#_M1003_d N_A_998_115#_M1012_g N_A_998_115#_M1006_g
+ N_A_998_115#_c_1599_n N_A_998_115#_c_1639_n N_A_998_115#_c_1572_n
+ N_A_998_115#_c_1554_n N_A_998_115#_c_1557_n N_A_998_115#_c_1558_n
+ N_A_998_115#_c_1559_n N_A_998_115#_c_1561_n N_A_998_115#_c_1562_n
+ N_A_998_115#_c_1563_n N_A_998_115#_c_1564_n N_A_998_115#_c_1565_n
+ N_A_998_115#_c_1567_n PM_SKY130_OSU_SC_12T_MS__DFFNR_L%A_998_115#
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%QN N_QN_M1016_s N_QN_M1011_s N_QN_M1008_g
+ N_QN_M1001_g N_QN_c_1700_n N_QN_c_1704_n N_QN_c_1706_n N_QN_c_1707_n
+ N_QN_c_1708_n N_QN_c_1709_n N_QN_c_1710_n N_QN_c_1711_n QN
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%QN
x_PM_SKY130_OSU_SC_12T_MS__DFFNR_L%Q N_Q_M1008_d N_Q_M1001_d N_Q_c_1791_n
+ N_Q_c_1795_n N_Q_c_1793_n N_Q_c_1794_n Q N_Q_c_1802_n
+ PM_SKY130_OSU_SC_12T_MS__DFFNR_L%Q
cc_1 N_GND_M1021_b N_RN_M1021_g 0.0616724f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_RN_M1021_g 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_RN_M1021_g 0.00606474f $X=1.125 $Y=0.152 $X2=0.475 $Y2=0.835
cc_4 N_GND_c_4_p N_RN_M1021_g 0.00359543f $X=1.21 $Y=0.74 $X2=0.475 $Y2=0.835
cc_5 N_GND_c_5_p N_RN_M1021_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.475 $Y2=0.835
cc_6 N_GND_M1021_b N_RN_c_383_n 0.0376794f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.99
cc_7 N_GND_M1021_b N_RN_M1004_g 0.0288885f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.235
cc_8 N_GND_M1021_b N_RN_c_385_n 0.020332f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.825
cc_9 N_GND_M1021_b N_RN_c_386_n 0.0149094f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_10 N_GND_M1021_b N_A_110_115#_c_416_n 0.0181101f $X=-0.05 $Y=0 $X2=0.475
+ $Y2=3.235
cc_11 N_GND_c_4_p N_A_110_115#_c_416_n 0.00502587f $X=1.21 $Y=0.74 $X2=0.475
+ $Y2=3.235
cc_12 N_GND_c_12_p N_A_110_115#_c_416_n 0.00606474f $X=1.985 $Y=0.152 $X2=0.475
+ $Y2=3.235
cc_13 N_GND_c_5_p N_A_110_115#_c_416_n 0.00468827f $X=9.175 $Y=0.19 $X2=0.475
+ $Y2=3.235
cc_14 N_GND_M1021_b N_A_110_115#_M1015_g 0.060904f $X=-0.05 $Y=0 $X2=0.53
+ $Y2=1.825
cc_15 N_GND_M1021_b N_A_110_115#_c_421_n 0.0603547f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_16 N_GND_c_16_p N_A_110_115#_c_421_n 0.00335985f $X=7.9 $Y=0.74 $X2=0 $Y2=0
cc_17 N_GND_M1021_b N_A_110_115#_M1030_g 0.0560323f $X=-0.05 $Y=0 $X2=0.32
+ $Y2=2.85
cc_18 N_GND_M1021_b N_A_110_115#_c_424_n 0.0181101f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_19 N_GND_c_19_p N_A_110_115#_c_424_n 0.00606474f $X=7.815 $Y=0.152 $X2=0
+ $Y2=0
cc_20 N_GND_c_16_p N_A_110_115#_c_424_n 0.00502587f $X=7.9 $Y=0.74 $X2=0 $Y2=0
cc_21 N_GND_c_5_p N_A_110_115#_c_424_n 0.00468827f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_22 N_GND_M1021_b N_A_110_115#_c_428_n 0.00155788f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_23 N_GND_c_3_p N_A_110_115#_c_428_n 0.0075272f $X=1.125 $Y=0.152 $X2=0 $Y2=0
cc_24 N_GND_c_4_p N_A_110_115#_c_428_n 0.0140971f $X=1.21 $Y=0.74 $X2=0 $Y2=0
cc_25 N_GND_c_5_p N_A_110_115#_c_428_n 0.00474817f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_26 N_GND_M1021_b N_A_110_115#_c_432_n 0.0021895f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_27 N_GND_M1021_b N_A_110_115#_c_433_n 0.0188948f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_28 N_GND_M1021_b N_A_110_115#_c_434_n 0.00886322f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_29 N_GND_c_4_p N_A_110_115#_c_434_n 4.91534e-19 $X=1.21 $Y=0.74 $X2=0 $Y2=0
cc_30 N_GND_M1021_b N_A_110_115#_c_436_n 0.0159872f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_31 N_GND_M1021_b N_A_110_115#_c_437_n 0.0162344f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_32 N_GND_M1018_s N_A_110_115#_c_438_n 5.79494e-19 $X=1.085 $Y=0.575 $X2=0
+ $Y2=0
cc_33 N_GND_M1005_d N_A_110_115#_c_438_n 0.00254601f $X=1.93 $Y=0.575 $X2=0
+ $Y2=0
cc_34 N_GND_M1007_s N_A_110_115#_c_438_n 0.00263312f $X=2.465 $Y=0.575 $X2=0
+ $Y2=0
cc_35 N_GND_M1027_d N_A_110_115#_c_438_n 0.00722605f $X=4.2 $Y=0.575 $X2=0 $Y2=0
cc_36 N_GND_M1023_d N_A_110_115#_c_438_n 0.00362717f $X=5.95 $Y=0.575 $X2=0
+ $Y2=0
cc_37 N_GND_M1012_s N_A_110_115#_c_438_n 0.00254601f $X=6.915 $Y=0.575 $X2=0
+ $Y2=0
cc_38 N_GND_M1013_d N_A_110_115#_c_438_n 0.00227813f $X=7.76 $Y=0.575 $X2=0
+ $Y2=0
cc_39 N_GND_M1021_b N_A_110_115#_c_438_n 0.0161221f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_40 N_GND_c_12_p N_A_110_115#_c_438_n 0.00424466f $X=1.985 $Y=0.152 $X2=0
+ $Y2=0
cc_41 N_GND_c_41_p N_A_110_115#_c_438_n 0.0070662f $X=2.07 $Y=0.74 $X2=0 $Y2=0
cc_42 N_GND_c_42_p N_A_110_115#_c_438_n 0.00599718f $X=2.505 $Y=0.152 $X2=0
+ $Y2=0
cc_43 N_GND_c_43_p N_A_110_115#_c_438_n 0.012085f $X=2.59 $Y=0.755 $X2=0 $Y2=0
cc_44 N_GND_c_44_p N_A_110_115#_c_438_n 0.0196453f $X=4.255 $Y=0.152 $X2=0 $Y2=0
cc_45 N_GND_c_45_p N_A_110_115#_c_438_n 0.00720909f $X=4.34 $Y=0.74 $X2=0 $Y2=0
cc_46 N_GND_c_46_p N_A_110_115#_c_438_n 0.0196423f $X=6.005 $Y=0.152 $X2=0 $Y2=0
cc_47 N_GND_c_47_p N_A_110_115#_c_438_n 0.0141132f $X=6.09 $Y=0.755 $X2=0 $Y2=0
cc_48 N_GND_c_48_p N_A_110_115#_c_438_n 0.00580139f $X=6.955 $Y=0.152 $X2=0
+ $Y2=0
cc_49 N_GND_c_49_p N_A_110_115#_c_438_n 0.00632479f $X=7.04 $Y=0.74 $X2=0 $Y2=0
cc_50 N_GND_c_19_p N_A_110_115#_c_438_n 0.00815276f $X=7.815 $Y=0.152 $X2=0
+ $Y2=0
cc_51 N_GND_c_16_p N_A_110_115#_c_438_n 0.00655132f $X=7.9 $Y=0.74 $X2=0 $Y2=0
cc_52 N_GND_M1018_s N_A_110_115#_c_458_n 0.0017057f $X=1.085 $Y=0.575 $X2=0
+ $Y2=0
cc_53 N_GND_M1021_b N_A_110_115#_c_458_n 0.00113133f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_54 N_GND_c_4_p N_A_110_115#_c_458_n 0.00660647f $X=1.21 $Y=0.74 $X2=0 $Y2=0
cc_55 N_GND_c_12_p N_A_110_115#_c_458_n 0.00391005f $X=1.985 $Y=0.152 $X2=0
+ $Y2=0
cc_56 N_GND_M1021_b N_A_110_115#_c_462_n 0.00487424f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_57 N_GND_M1021_b N_A_110_115#_c_463_n 0.00285541f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_58 N_GND_M1021_b N_A_110_115#_c_464_n 0.0015072f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_59 N_GND_c_4_p N_A_110_115#_c_464_n 0.00797325f $X=1.21 $Y=0.74 $X2=0 $Y2=0
cc_60 N_GND_M1021_b N_A_110_115#_c_466_n 0.0450929f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_61 N_GND_c_4_p N_A_110_115#_c_466_n 0.00336f $X=1.21 $Y=0.74 $X2=0 $Y2=0
cc_62 N_GND_M1021_b N_A_110_115#_c_468_n 0.00428422f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_63 N_GND_c_16_p N_A_110_115#_c_468_n 0.00849521f $X=7.9 $Y=0.74 $X2=0 $Y2=0
cc_64 N_GND_M1021_b N_A_342_442#_M1005_g 0.087851f $X=-0.05 $Y=0 $X2=0.53
+ $Y2=1.825
cc_65 N_GND_c_12_p N_A_342_442#_M1005_g 0.00606474f $X=1.985 $Y=0.152 $X2=0.53
+ $Y2=1.825
cc_66 N_GND_c_41_p N_A_342_442#_M1005_g 0.00502587f $X=2.07 $Y=0.74 $X2=0.53
+ $Y2=1.825
cc_67 N_GND_c_5_p N_A_342_442#_M1005_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.53
+ $Y2=1.825
cc_68 N_GND_M1021_b N_A_342_442#_c_618_n 0.0182652f $X=-0.05 $Y=0 $X2=0.32
+ $Y2=2.85
cc_69 N_GND_M1021_b N_A_342_442#_c_619_n 0.0217838f $X=-0.05 $Y=0 $X2=0.53
+ $Y2=1.825
cc_70 N_GND_c_43_p N_A_342_442#_c_619_n 0.00673409f $X=2.59 $Y=0.755 $X2=0.53
+ $Y2=1.825
cc_71 N_GND_M1021_b N_A_342_442#_c_621_n 0.00653128f $X=-0.05 $Y=0 $X2=0.32
+ $Y2=2.85
cc_72 N_GND_c_41_p N_A_342_442#_c_621_n 0.00470355f $X=2.07 $Y=0.74 $X2=0.32
+ $Y2=2.85
cc_73 N_GND_M1021_b N_A_342_442#_c_623_n 0.00198494f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_74 N_GND_M1021_b N_A_342_442#_c_624_n 0.0066411f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_75 N_GND_M1021_b N_A_342_442#_c_625_n 0.0245154f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_76 N_GND_M1021_b N_A_342_442#_c_626_n 0.00311983f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_77 N_GND_c_44_p N_A_342_442#_c_626_n 0.0147897f $X=4.255 $Y=0.152 $X2=0 $Y2=0
cc_78 N_GND_c_5_p N_A_342_442#_c_626_n 0.0098977f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_79 N_GND_M1021_b N_D_M1007_g 0.0418787f $X=-0.05 $Y=0 $X2=0.475 $Y2=0.835
cc_80 N_GND_c_43_p N_D_M1007_g 0.00509529f $X=2.59 $Y=0.755 $X2=0.475 $Y2=0.835
cc_81 N_GND_c_44_p N_D_M1007_g 0.00606474f $X=4.255 $Y=0.152 $X2=0.475 $Y2=0.835
cc_82 N_GND_c_5_p N_D_M1007_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.475 $Y2=0.835
cc_83 N_GND_M1021_b N_D_M1028_g 0.0359102f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.235
cc_84 N_GND_M1021_b D 0.00973922f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.99
cc_85 N_GND_M1021_b N_D_c_703_n 0.00311208f $X=-0.05 $Y=0 $X2=0.53 $Y2=1.825
cc_86 N_GND_M1021_b N_D_c_704_n 0.0324288f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_87 N_GND_M1021_b N_A_618_424#_c_739_n 0.00609317f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_88 N_GND_M1021_b N_A_618_424#_c_740_n 0.00920685f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_89 N_GND_M1021_b N_A_618_424#_c_741_n 0.0254608f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_90 N_GND_M1021_b N_A_618_424#_c_742_n 0.008127f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_91 N_GND_M1021_b N_A_618_424#_c_743_n 0.0267352f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_92 N_GND_M1021_b N_A_618_424#_c_744_n 0.00482713f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_93 N_GND_M1021_b N_A_618_424#_c_745_n 5.00459e-19 $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_94 N_GND_M1021_b N_A_618_424#_c_746_n 0.0195179f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_95 N_GND_c_47_p N_A_618_424#_c_746_n 0.00147792f $X=6.09 $Y=0.755 $X2=0 $Y2=0
cc_96 N_GND_c_49_p N_A_618_424#_c_746_n 0.00354837f $X=7.04 $Y=0.74 $X2=0 $Y2=0
cc_97 N_GND_M1021_b N_A_618_424#_c_749_n 0.00401094f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_98 N_GND_c_48_p N_A_618_424#_c_749_n 0.0121407f $X=6.955 $Y=0.152 $X2=0 $Y2=0
cc_99 N_GND_c_49_p N_A_618_424#_c_749_n 0.01517f $X=7.04 $Y=0.74 $X2=0 $Y2=0
cc_100 N_GND_c_5_p N_A_618_424#_c_749_n 0.0108718f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_101 N_GND_M1021_b N_A_618_424#_c_753_n 0.00889426f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_102 N_GND_M1021_b N_A_618_424#_c_754_n 0.0338168f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_103 N_GND_M1021_b N_A_618_424#_c_755_n 0.00714094f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_104 N_GND_M1021_b N_A_618_424#_c_756_n 0.019097f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_105 N_GND_M1021_b N_A_618_424#_c_757_n 0.0025628f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_106 N_GND_M1021_b N_A_618_424#_c_758_n 0.00276905f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_107 N_GND_M1021_b N_A_618_424#_c_759_n 0.00119864f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_108 N_GND_M1021_b N_A_618_424#_c_760_n 0.00296941f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_109 N_GND_M1021_b N_A_618_424#_c_761_n 0.0101616f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_110 N_GND_M1021_b N_A_618_424#_c_762_n 0.0244095f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_111 N_GND_M1021_b N_A_618_424#_c_763_n 0.0173906f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_112 N_GND_c_44_p N_A_618_424#_c_763_n 0.00606474f $X=4.255 $Y=0.152 $X2=0
+ $Y2=0
cc_113 N_GND_c_5_p N_A_618_424#_c_763_n 0.00468827f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_114 N_GND_M1021_b N_A_618_424#_c_766_n 0.0174883f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_115 N_GND_c_46_p N_A_618_424#_c_766_n 0.00606474f $X=6.005 $Y=0.152 $X2=0
+ $Y2=0
cc_116 N_GND_c_5_p N_A_618_424#_c_766_n 0.00468827f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_117 N_GND_M1021_b N_A_618_424#_c_769_n 0.0220032f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_118 N_GND_M1021_b N_A_217_605#_M1027_g 0.0171926f $X=-0.05 $Y=0 $X2=0.32
+ $Y2=1.825
cc_119 N_GND_c_44_p N_A_217_605#_M1027_g 0.00606474f $X=4.255 $Y=0.152 $X2=0.32
+ $Y2=1.825
cc_120 N_GND_c_45_p N_A_217_605#_M1027_g 0.00308284f $X=4.34 $Y=0.74 $X2=0.32
+ $Y2=1.825
cc_121 N_GND_c_5_p N_A_217_605#_M1027_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.32
+ $Y2=1.825
cc_122 N_GND_M1021_b N_A_217_605#_M1025_g 0.0170177f $X=-0.05 $Y=0 $X2=0.325
+ $Y2=2.85
cc_123 N_GND_c_45_p N_A_217_605#_M1025_g 0.00308284f $X=4.34 $Y=0.74 $X2=0.325
+ $Y2=2.85
cc_124 N_GND_c_46_p N_A_217_605#_M1025_g 0.00606474f $X=6.005 $Y=0.152 $X2=0.325
+ $Y2=2.85
cc_125 N_GND_c_5_p N_A_217_605#_M1025_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.325
+ $Y2=2.85
cc_126 N_GND_M1021_b N_A_217_605#_c_1005_n 0.0105855f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_127 N_GND_M1021_b N_A_217_605#_c_1006_n 0.0105265f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_128 N_GND_M1021_b N_A_217_605#_c_1007_n 0.0240311f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_129 N_GND_c_45_p N_A_217_605#_c_1007_n 9.93645e-19 $X=4.34 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_GND_M1021_b N_A_217_605#_c_1009_n 0.0232417f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_131 N_GND_M1021_b N_A_217_605#_c_1010_n 0.011276f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_132 N_GND_M1021_b N_A_217_605#_c_1011_n 0.0127277f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_133 N_GND_M1021_b N_A_217_605#_c_1012_n 0.00259716f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_134 N_GND_M1021_b N_A_217_605#_c_1013_n 0.00871176f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_135 N_GND_M1021_b N_A_217_605#_c_1014_n 0.0335787f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_136 N_GND_M1021_b N_A_217_605#_c_1015_n 0.00340906f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_137 N_GND_M1021_b N_A_217_605#_c_1016_n 0.00210386f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_138 N_GND_c_45_p N_A_217_605#_c_1016_n 0.00441035f $X=4.34 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_GND_M1021_b N_A_217_605#_c_1018_n 0.017579f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_140 N_GND_c_12_p N_A_217_605#_c_1018_n 0.00734006f $X=1.985 $Y=0.152 $X2=0
+ $Y2=0
cc_141 N_GND_c_5_p N_A_217_605#_c_1018_n 0.00475776f $X=9.175 $Y=0.19 $X2=0
+ $Y2=0
cc_142 N_GND_M1021_b N_CK_c_1135_n 0.0173059f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.655
cc_143 N_GND_c_44_p N_CK_c_1135_n 0.00606474f $X=4.255 $Y=0.152 $X2=0.475
+ $Y2=1.655
cc_144 N_GND_c_5_p N_CK_c_1135_n 0.00468827f $X=9.175 $Y=0.19 $X2=0.475
+ $Y2=1.655
cc_145 N_GND_M1021_b N_CK_c_1138_n 0.0203057f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.99
cc_146 N_GND_M1021_b N_CK_c_1139_n 0.0187566f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.235
cc_147 N_GND_M1021_b N_CK_c_1140_n 0.00755029f $X=-0.05 $Y=0 $X2=0.475 $Y2=3.235
cc_148 N_GND_M1021_b N_CK_M1017_g 0.032457f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.99
cc_149 N_GND_M1021_b N_CK_c_1142_n 0.0559794f $X=-0.05 $Y=0 $X2=0.53 $Y2=1.825
cc_150 N_GND_M1021_b N_CK_M1003_g 0.0319667f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_151 N_GND_M1021_b N_CK_c_1144_n 0.0187483f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_152 N_GND_M1021_b N_CK_M1020_g 0.0322593f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_153 N_GND_c_46_p N_CK_M1020_g 0.00606474f $X=6.005 $Y=0.152 $X2=0 $Y2=0
cc_154 N_GND_c_5_p N_CK_M1020_g 0.00468827f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_155 N_GND_M1021_b N_CK_c_1148_n 0.0185814f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_156 N_GND_c_47_p N_CK_c_1148_n 0.00313598f $X=6.09 $Y=0.755 $X2=0 $Y2=0
cc_157 N_GND_c_48_p N_CK_c_1148_n 0.00577402f $X=6.955 $Y=0.152 $X2=0 $Y2=0
cc_158 N_GND_c_49_p N_CK_c_1148_n 0.00384149f $X=7.04 $Y=0.74 $X2=0 $Y2=0
cc_159 N_GND_c_5_p N_CK_c_1148_n 0.00468827f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_160 N_GND_M1021_b N_CK_c_1153_n 0.0293856f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_161 N_GND_M1021_b N_CK_c_1154_n 0.0441689f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_162 N_GND_M1021_b N_CK_c_1155_n 0.0141736f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_163 N_GND_M1021_b N_CK_c_1156_n 0.00426512f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_164 N_GND_M1021_b N_CK_c_1157_n 0.00426512f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_165 N_GND_M1021_b N_CK_c_1158_n 0.0144521f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_166 N_GND_M1021_b N_CK_c_1159_n 0.00169461f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_167 N_GND_M1021_b N_CK_c_1160_n 0.00465235f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_168 N_GND_M1021_b N_CK_c_1161_n 0.00323244f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_169 N_GND_M1021_b CK 0.00178225f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_170 N_GND_M1021_b N_CK_c_1163_n 0.0333891f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_171 N_GND_M1021_b N_CK_c_1164_n 0.00141731f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_172 N_GND_M1021_b N_A_1160_89#_M1009_g 0.00746385f $X=-0.05 $Y=0 $X2=0.53
+ $Y2=1.825
cc_173 N_GND_M1021_b N_A_1160_89#_M1016_g 0.0259924f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_174 N_GND_c_16_p N_A_1160_89#_M1016_g 0.00359543f $X=7.9 $Y=0.74 $X2=0 $Y2=0
cc_175 N_GND_c_175_p N_A_1160_89#_M1016_g 0.00606474f $X=8.765 $Y=0.152 $X2=0
+ $Y2=0
cc_176 N_GND_c_176_p N_A_1160_89#_M1016_g 0.00308284f $X=8.85 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_GND_c_5_p N_A_1160_89#_M1016_g 0.00468827f $X=9.175 $Y=0.19 $X2=0 $Y2=0
cc_178 N_GND_M1021_b N_A_1160_89#_c_1345_n 0.0161097f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_179 N_GND_c_46_p N_A_1160_89#_c_1345_n 0.00606474f $X=6.005 $Y=0.152 $X2=0
+ $Y2=0
cc_180 N_GND_c_47_p N_A_1160_89#_c_1345_n 0.00315235f $X=6.09 $Y=0.755 $X2=0
+ $Y2=0
cc_181 N_GND_c_5_p N_A_1160_89#_c_1345_n 0.00468827f $X=9.175 $Y=0.19 $X2=0
+ $Y2=0
cc_182 N_GND_M1021_b N_A_1160_89#_c_1349_n 0.00990896f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_183 N_GND_M1021_b N_A_1160_89#_c_1350_n 0.0116478f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_184 N_GND_M1021_b N_A_1160_89#_c_1351_n 0.00918377f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_185 N_GND_M1021_b N_A_1160_89#_c_1352_n 0.0136411f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_186 N_GND_M1021_b N_A_1160_89#_c_1353_n 0.0341464f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_187 N_GND_M1021_b N_A_1160_89#_c_1354_n 0.00495925f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_188 N_GND_M1021_b N_A_1160_89#_c_1355_n 0.011707f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_189 N_GND_c_19_p N_A_1160_89#_c_1355_n 0.0075556f $X=7.815 $Y=0.152 $X2=0
+ $Y2=0
cc_190 N_GND_c_5_p N_A_1160_89#_c_1355_n 0.00475776f $X=9.175 $Y=0.19 $X2=0
+ $Y2=0
cc_191 N_GND_M1021_b N_A_1160_89#_c_1358_n 0.00350278f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_192 N_GND_M1021_b N_A_1160_89#_c_1359_n 0.00183023f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_193 N_GND_c_47_p N_A_1160_89#_c_1359_n 4.59543e-19 $X=6.09 $Y=0.755 $X2=0
+ $Y2=0
cc_194 N_GND_M1021_b N_A_1160_89#_c_1361_n 0.0272158f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_195 N_GND_c_47_p N_A_1160_89#_c_1361_n 0.00110843f $X=6.09 $Y=0.755 $X2=0
+ $Y2=0
cc_196 N_GND_M1021_b N_A_1160_89#_c_1363_n 0.00139765f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_197 N_GND_M1021_b N_A_1160_89#_c_1364_n 0.00795534f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_198 N_GND_M1021_b N_A_1160_89#_c_1365_n 0.00111103f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_199 N_GND_M1021_b N_A_1160_89#_c_1366_n 0.00690501f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_200 N_GND_M1021_b N_A_1160_89#_c_1367_n 0.00198809f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_201 N_GND_M1021_b N_A_1160_89#_c_1368_n 0.00201111f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_202 N_GND_M1021_b N_A_1160_89#_c_1369_n 0.00280684f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_203 N_GND_M1021_b N_A_1160_89#_c_1370_n 0.0181474f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_204 N_GND_M1021_b N_A_1160_89#_c_1371_n 0.038213f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_205 N_GND_M1021_b N_A_1160_89#_c_1372_n 0.0119185f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_206 N_GND_M1021_b N_A_1160_89#_c_1373_n 0.0294757f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_207 N_GND_M1021_b N_A_1160_89#_c_1374_n 0.0171478f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_208 N_GND_M1021_b N_A_998_115#_M1012_g 0.0279847f $X=-0.05 $Y=0 $X2=0.32
+ $Y2=1.825
cc_209 N_GND_c_49_p N_A_998_115#_M1012_g 0.00502587f $X=7.04 $Y=0.74 $X2=0.32
+ $Y2=1.825
cc_210 N_GND_c_19_p N_A_998_115#_M1012_g 0.00606474f $X=7.815 $Y=0.152 $X2=0.32
+ $Y2=1.825
cc_211 N_GND_c_5_p N_A_998_115#_M1012_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.32
+ $Y2=1.825
cc_212 N_GND_M1021_b N_A_998_115#_M1006_g 0.0469083f $X=-0.05 $Y=0 $X2=0.53
+ $Y2=1.825
cc_213 N_GND_M1021_b N_A_998_115#_c_1554_n 0.00312748f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_214 N_GND_c_46_p N_A_998_115#_c_1554_n 0.0150341f $X=6.005 $Y=0.152 $X2=0
+ $Y2=0
cc_215 N_GND_c_5_p N_A_998_115#_c_1554_n 0.00994746f $X=9.175 $Y=0.19 $X2=0
+ $Y2=0
cc_216 N_GND_M1021_b N_A_998_115#_c_1557_n 0.00241727f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_217 N_GND_M1021_b N_A_998_115#_c_1558_n 0.00125111f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_218 N_GND_M1021_b N_A_998_115#_c_1559_n 0.0148243f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_219 N_GND_c_47_p N_A_998_115#_c_1559_n 7.83815e-19 $X=6.09 $Y=0.755 $X2=0
+ $Y2=0
cc_220 N_GND_M1021_b N_A_998_115#_c_1561_n 0.00209768f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_221 N_GND_M1021_b N_A_998_115#_c_1562_n 0.0113462f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_222 N_GND_M1021_b N_A_998_115#_c_1563_n 0.00904057f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_223 N_GND_M1021_b N_A_998_115#_c_1564_n 5.61996e-19 $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_224 N_GND_M1021_b N_A_998_115#_c_1565_n 0.00676232f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_225 N_GND_c_49_p N_A_998_115#_c_1565_n 0.00491851f $X=7.04 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_GND_M1021_b N_A_998_115#_c_1567_n 0.043899f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_227 N_GND_c_49_p N_A_998_115#_c_1567_n 0.00154898f $X=7.04 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_GND_M1021_b N_QN_M1008_g 0.0651437f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.825
cc_229 N_GND_c_176_p N_QN_M1008_g 0.00308284f $X=8.85 $Y=0.74 $X2=0.32 $Y2=1.825
cc_230 N_GND_c_5_p N_QN_M1008_g 0.00468827f $X=9.175 $Y=0.19 $X2=0.32 $Y2=1.825
cc_231 N_GND_M1021_b N_QN_M1001_g 0.0186095f $X=-0.05 $Y=0 $X2=0.53 $Y2=1.825
cc_232 N_GND_M1021_b N_QN_c_1700_n 0.00776412f $X=-0.05 $Y=0 $X2=0.325 $Y2=2.85
cc_233 N_GND_c_16_p N_QN_c_1700_n 0.0140971f $X=7.9 $Y=0.74 $X2=0.325 $Y2=2.85
cc_234 N_GND_c_175_p N_QN_c_1700_n 0.00736239f $X=8.765 $Y=0.152 $X2=0.325
+ $Y2=2.85
cc_235 N_GND_c_5_p N_QN_c_1700_n 0.00476261f $X=9.175 $Y=0.19 $X2=0.325 $Y2=2.85
cc_236 N_GND_M1021_b N_QN_c_1704_n 0.0134367f $X=-0.05 $Y=0 $X2=0.53 $Y2=1.825
cc_237 N_GND_c_176_p N_QN_c_1704_n 0.00779875f $X=8.85 $Y=0.74 $X2=0.53
+ $Y2=1.825
cc_238 N_GND_M1021_b N_QN_c_1706_n 0.00232247f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_239 N_GND_M1021_b N_QN_c_1707_n 0.0138306f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_240 N_GND_M1021_b N_QN_c_1708_n 0.00434805f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_241 N_GND_M1021_b N_QN_c_1709_n 0.00362324f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_242 N_GND_M1021_b N_QN_c_1710_n 0.0291868f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_243 N_GND_M1021_b N_QN_c_1711_n 0.00138285f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_244 N_GND_M1021_b QN 0.00270537f $X=-0.05 $Y=0 $X2=0 $Y2=0
cc_245 N_GND_M1021_b N_Q_c_1791_n 0.0098062f $X=-0.05 $Y=0 $X2=0.32 $Y2=1.825
cc_246 N_GND_c_5_p N_Q_c_1791_n 0.00467398f $X=9.175 $Y=0.19 $X2=0.32 $Y2=1.825
cc_247 N_GND_M1021_b N_Q_c_1793_n 0.0625704f $X=-0.05 $Y=0 $X2=0.32 $Y2=2.85
cc_248 N_GND_M1021_b N_Q_c_1794_n 0.0189963f $X=-0.05 $Y=0 $X2=0.53 $Y2=1.825
cc_249 N_VDD_M1004_b N_RN_M1004_g 0.0266406f $X=-0.05 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_250 N_VDD_c_250_p N_RN_M1004_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_251 N_VDD_c_251_p N_RN_M1004_g 0.00606474f $X=1.915 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_252 N_VDD_c_252_p N_RN_M1004_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.475
+ $Y2=3.235
cc_253 N_VDD_M1004_s N_RN_c_386_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32
+ $Y2=2.85
cc_254 N_VDD_M1004_b N_RN_c_386_n 0.00618364f $X=-0.05 $Y=2.425 $X2=0.32
+ $Y2=2.85
cc_255 N_VDD_c_250_p N_RN_c_386_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_256 N_VDD_M1004_s RN 0.016276f $X=0.135 $Y=2.605 $X2=0.325 $Y2=2.85
cc_257 N_VDD_c_250_p RN 0.00522047f $X=0.26 $Y=3.635 $X2=0.325 $Y2=2.85
cc_258 N_VDD_M1004_b N_A_110_115#_M1015_g 0.0463013f $X=-0.05 $Y=2.425 $X2=0.53
+ $Y2=1.825
cc_259 N_VDD_c_251_p N_A_110_115#_M1015_g 0.00606474f $X=1.915 $Y=4.287 $X2=0.53
+ $Y2=1.825
cc_260 N_VDD_c_252_p N_A_110_115#_M1015_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_261 N_VDD_M1004_b N_A_110_115#_M1030_g 0.0450939f $X=-0.05 $Y=2.425 $X2=0.32
+ $Y2=2.85
cc_262 N_VDD_c_262_p N_A_110_115#_M1030_g 0.00606474f $X=7.745 $Y=4.287 $X2=0.32
+ $Y2=2.85
cc_263 N_VDD_c_263_p N_A_110_115#_M1030_g 0.00713292f $X=7.83 $Y=3.275 $X2=0.32
+ $Y2=2.85
cc_264 N_VDD_c_252_p N_A_110_115#_M1030_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.32
+ $Y2=2.85
cc_265 N_VDD_M1004_b N_A_110_115#_c_432_n 0.00549797f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_266 N_VDD_c_251_p N_A_110_115#_c_432_n 0.00757793f $X=1.915 $Y=4.287 $X2=0
+ $Y2=0
cc_267 N_VDD_c_252_p N_A_110_115#_c_432_n 0.00476261f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_268 N_VDD_M1004_b N_A_342_442#_M1002_g 0.0430317f $X=-0.05 $Y=2.425 $X2=0.32
+ $Y2=1.825
cc_269 N_VDD_c_251_p N_A_342_442#_M1002_g 0.00606474f $X=1.915 $Y=4.287 $X2=0.32
+ $Y2=1.825
cc_270 N_VDD_c_270_p N_A_342_442#_M1002_g 0.00713292f $X=2 $Y=3.275 $X2=0.32
+ $Y2=1.825
cc_271 N_VDD_c_252_p N_A_342_442#_M1002_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.32
+ $Y2=1.825
cc_272 N_VDD_M1028_s N_A_342_442#_c_633_n 0.0125004f $X=2.465 $Y=2.605 $X2=0.325
+ $Y2=2.85
cc_273 N_VDD_M1004_b N_A_342_442#_c_633_n 0.0199377f $X=-0.05 $Y=2.425 $X2=0.325
+ $Y2=2.85
cc_274 N_VDD_c_274_p N_A_342_442#_c_633_n 0.00952036f $X=2.59 $Y=3.295 $X2=0.325
+ $Y2=2.85
cc_275 N_VDD_M1004_b N_A_342_442#_c_636_n 0.00313975f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_276 N_VDD_c_276_p N_A_342_442#_c_636_n 0.0151129f $X=4.255 $Y=4.287 $X2=0
+ $Y2=0
cc_277 N_VDD_c_252_p N_A_342_442#_c_636_n 0.00958198f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_278 N_VDD_M1004_b N_A_342_442#_c_624_n 0.0146567f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_279 N_VDD_c_270_p N_A_342_442#_c_624_n 0.00826787f $X=2 $Y=3.275 $X2=0 $Y2=0
cc_280 N_VDD_M1004_b N_A_342_442#_c_625_n 0.015181f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_281 N_VDD_c_270_p N_A_342_442#_c_625_n 9.61776e-19 $X=2 $Y=3.275 $X2=0 $Y2=0
cc_282 N_VDD_M1004_b N_D_M1028_g 0.0219788f $X=-0.05 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_283 N_VDD_c_270_p N_D_M1028_g 0.00284049f $X=2 $Y=3.275 $X2=0.475 $Y2=3.235
cc_284 N_VDD_c_274_p N_D_M1028_g 0.00636672f $X=2.59 $Y=3.295 $X2=0.475
+ $Y2=3.235
cc_285 N_VDD_c_276_p N_D_M1028_g 0.00606474f $X=4.255 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_286 N_VDD_c_252_p N_D_M1028_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.475
+ $Y2=3.235
cc_287 N_VDD_M1004_b N_A_618_424#_M1024_g 0.020128f $X=-0.05 $Y=2.425 $X2=0.32
+ $Y2=1.825
cc_288 N_VDD_c_276_p N_A_618_424#_M1024_g 0.00606474f $X=4.255 $Y=4.287 $X2=0.32
+ $Y2=1.825
cc_289 N_VDD_c_252_p N_A_618_424#_M1024_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.32
+ $Y2=1.825
cc_290 N_VDD_M1004_b N_A_618_424#_M1000_g 0.0201163f $X=-0.05 $Y=2.425 $X2=0.53
+ $Y2=1.825
cc_291 N_VDD_c_291_p N_A_618_424#_M1000_g 0.00606474f $X=6.005 $Y=4.287 $X2=0.53
+ $Y2=1.825
cc_292 N_VDD_c_252_p N_A_618_424#_M1000_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_293 N_VDD_M1004_b N_A_618_424#_c_776_n 0.00156053f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_294 N_VDD_c_262_p N_A_618_424#_c_776_n 0.00736239f $X=7.745 $Y=4.287 $X2=0
+ $Y2=0
cc_295 N_VDD_c_252_p N_A_618_424#_c_776_n 0.00476261f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_296 N_VDD_M1004_b N_A_618_424#_c_779_n 0.0164285f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_297 N_VDD_M1004_b N_A_618_424#_c_758_n 6.42499e-19 $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_298 N_VDD_M1004_b N_A_618_424#_c_759_n 0.0022456f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_299 N_VDD_M1004_b N_A_618_424#_c_761_n 0.00489351f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_300 N_VDD_M1004_b N_A_618_424#_c_762_n 0.00487135f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_301 N_VDD_M1004_b N_A_618_424#_c_769_n 0.00485139f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_302 N_VDD_M1004_b N_A_217_605#_M1022_g 0.0192219f $X=-0.05 $Y=2.425 $X2=0.53
+ $Y2=1.825
cc_303 N_VDD_c_276_p N_A_217_605#_M1022_g 0.00606474f $X=4.255 $Y=4.287 $X2=0.53
+ $Y2=1.825
cc_304 N_VDD_c_304_p N_A_217_605#_M1022_g 0.00337744f $X=4.34 $Y=3.295 $X2=0.53
+ $Y2=1.825
cc_305 N_VDD_c_252_p N_A_217_605#_M1022_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_306 N_VDD_M1004_b N_A_217_605#_M1014_g 0.0181098f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_307 N_VDD_c_304_p N_A_217_605#_M1014_g 0.00337744f $X=4.34 $Y=3.295 $X2=0
+ $Y2=0
cc_308 N_VDD_c_291_p N_A_217_605#_M1014_g 0.00606474f $X=6.005 $Y=4.287 $X2=0
+ $Y2=0
cc_309 N_VDD_c_252_p N_A_217_605#_M1014_g 0.00468827f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_310 N_VDD_c_304_p N_A_217_605#_c_1009_n 8.24975e-19 $X=4.34 $Y=3.295 $X2=0
+ $Y2=0
cc_311 N_VDD_M1004_b N_A_217_605#_c_1010_n 0.0163203f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_312 N_VDD_c_251_p N_A_217_605#_c_1010_n 0.00745733f $X=1.915 $Y=4.287 $X2=0
+ $Y2=0
cc_313 N_VDD_c_252_p N_A_217_605#_c_1010_n 0.00476261f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_314 N_VDD_M1004_b N_A_217_605#_c_1013_n 0.00424346f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_315 N_VDD_c_304_p N_A_217_605#_c_1013_n 0.004428f $X=4.34 $Y=3.295 $X2=0
+ $Y2=0
cc_316 N_VDD_M1004_b N_CK_M1017_g 0.0215131f $X=-0.05 $Y=2.425 $X2=0.32 $Y2=1.99
cc_317 N_VDD_c_276_p N_CK_M1017_g 0.00606474f $X=4.255 $Y=4.287 $X2=0.32
+ $Y2=1.99
cc_318 N_VDD_c_252_p N_CK_M1017_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.32 $Y2=1.99
cc_319 N_VDD_M1004_b N_CK_M1003_g 0.0214821f $X=-0.05 $Y=2.425 $X2=0.32 $Y2=2.85
cc_320 N_VDD_c_291_p N_CK_M1003_g 0.00606474f $X=6.005 $Y=4.287 $X2=0.32
+ $Y2=2.85
cc_321 N_VDD_c_252_p N_CK_M1003_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.32 $Y2=2.85
cc_322 N_VDD_M1004_b N_CK_c_1153_n 0.00880158f $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_323 N_VDD_M1004_b N_CK_M1029_g 0.0242017f $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_324 N_VDD_c_324_p N_CK_M1029_g 0.00409291f $X=6.09 $Y=3.21 $X2=0 $Y2=0
cc_325 N_VDD_c_262_p N_CK_M1029_g 0.00606474f $X=7.745 $Y=4.287 $X2=0 $Y2=0
cc_326 N_VDD_c_252_p N_CK_M1029_g 0.00468827f $X=9.175 $Y=4.25 $X2=0 $Y2=0
cc_327 N_VDD_M1004_b N_CK_c_1159_n 2.23352e-19 $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_328 N_VDD_M1004_b N_A_1160_89#_M1009_g 0.0178558f $X=-0.05 $Y=2.425 $X2=0.53
+ $Y2=1.825
cc_329 N_VDD_c_291_p N_A_1160_89#_M1009_g 0.00606474f $X=6.005 $Y=4.287 $X2=0.53
+ $Y2=1.825
cc_330 N_VDD_c_324_p N_A_1160_89#_M1009_g 0.00409291f $X=6.09 $Y=3.21 $X2=0.53
+ $Y2=1.825
cc_331 N_VDD_c_252_p N_A_1160_89#_M1009_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_332 N_VDD_M1004_b N_A_1160_89#_M1011_g 0.0412931f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_333 N_VDD_c_263_p N_A_1160_89#_M1011_g 0.00453298f $X=7.83 $Y=3.275 $X2=0
+ $Y2=0
cc_334 N_VDD_c_334_p N_A_1160_89#_M1011_g 0.00606474f $X=8.765 $Y=4.287 $X2=0
+ $Y2=0
cc_335 N_VDD_c_335_p N_A_1160_89#_M1011_g 0.00602599f $X=8.85 $Y=3.265 $X2=0
+ $Y2=0
cc_336 N_VDD_c_252_p N_A_1160_89#_M1011_g 0.00468827f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_337 N_VDD_M1004_b N_A_1160_89#_c_1354_n 0.00913729f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_338 N_VDD_M1004_b N_A_1160_89#_c_1385_n 0.00156053f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_339 N_VDD_c_262_p N_A_1160_89#_c_1385_n 0.00736239f $X=7.745 $Y=4.287 $X2=0
+ $Y2=0
cc_340 N_VDD_c_252_p N_A_1160_89#_c_1385_n 0.00476261f $X=9.175 $Y=4.25 $X2=0
+ $Y2=0
cc_341 N_VDD_M1004_b N_A_1160_89#_c_1388_n 0.00251697f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_342 N_VDD_M1004_b N_A_1160_89#_c_1389_n 0.00359218f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_343 N_VDD_M1004_b N_A_1160_89#_c_1358_n 0.0041567f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_344 N_VDD_M1004_b N_A_1160_89#_c_1364_n 0.0103988f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_345 N_VDD_c_324_p N_A_1160_89#_c_1364_n 0.00425473f $X=6.09 $Y=3.21 $X2=0
+ $Y2=0
cc_346 N_VDD_M1004_b N_A_1160_89#_c_1365_n 0.00604093f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_347 N_VDD_c_324_p N_A_1160_89#_c_1365_n 0.003295f $X=6.09 $Y=3.21 $X2=0 $Y2=0
cc_348 N_VDD_M1004_b N_A_1160_89#_c_1368_n 0.00238208f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_349 N_VDD_c_324_p N_A_1160_89#_c_1368_n 4.62798e-19 $X=6.09 $Y=3.21 $X2=0
+ $Y2=0
cc_350 N_VDD_M1004_b N_A_998_115#_M1006_g 0.0487718f $X=-0.05 $Y=2.425 $X2=0.53
+ $Y2=1.825
cc_351 N_VDD_c_262_p N_A_998_115#_M1006_g 0.00606474f $X=7.745 $Y=4.287 $X2=0.53
+ $Y2=1.825
cc_352 N_VDD_c_252_p N_A_998_115#_M1006_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_353 N_VDD_M1004_b N_A_998_115#_c_1572_n 0.00313975f $X=-0.05 $Y=2.425
+ $X2=0.53 $Y2=1.825
cc_354 N_VDD_c_291_p N_A_998_115#_c_1572_n 0.0149205f $X=6.005 $Y=4.287 $X2=0.53
+ $Y2=1.825
cc_355 N_VDD_c_252_p N_A_998_115#_c_1572_n 0.00958198f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_356 N_VDD_M1004_b N_A_998_115#_c_1562_n 0.00168314f $X=-0.05 $Y=2.425 $X2=0
+ $Y2=0
cc_357 N_VDD_M1004_b N_QN_M1001_g 0.051339f $X=-0.05 $Y=2.425 $X2=0.53 $Y2=1.825
cc_358 N_VDD_c_335_p N_QN_M1001_g 0.00601131f $X=8.85 $Y=3.265 $X2=0.53
+ $Y2=1.825
cc_359 N_VDD_c_252_p N_QN_M1001_g 0.00468827f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_360 N_VDD_c_360_p N_QN_M1001_g 0.00606474f $X=9.175 $Y=4.22 $X2=0.53
+ $Y2=1.825
cc_361 N_VDD_c_335_p N_QN_c_1707_n 0.00856258f $X=8.85 $Y=3.265 $X2=0 $Y2=0
cc_362 N_VDD_c_335_p N_QN_c_1710_n 2.00737e-19 $X=8.85 $Y=3.265 $X2=0 $Y2=0
cc_363 N_VDD_M1004_b N_QN_c_1711_n 0.0181975f $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_364 N_VDD_c_263_p N_QN_c_1711_n 0.0313352f $X=7.83 $Y=3.275 $X2=0 $Y2=0
cc_365 N_VDD_c_334_p N_QN_c_1711_n 0.00736239f $X=8.765 $Y=4.287 $X2=0 $Y2=0
cc_366 N_VDD_c_335_p N_QN_c_1711_n 0.0159141f $X=8.85 $Y=3.265 $X2=0 $Y2=0
cc_367 N_VDD_c_252_p N_QN_c_1711_n 0.00476261f $X=9.175 $Y=4.25 $X2=0 $Y2=0
cc_368 N_VDD_M1004_b QN 0.0110801f $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_369 N_VDD_M1004_b N_Q_c_1795_n 0.00508086f $X=-0.05 $Y=2.425 $X2=0.53
+ $Y2=1.825
cc_370 N_VDD_c_335_p N_Q_c_1795_n 0.00454099f $X=8.85 $Y=3.265 $X2=0.53
+ $Y2=1.825
cc_371 N_VDD_c_252_p N_Q_c_1795_n 0.00476261f $X=9.175 $Y=4.25 $X2=0.53
+ $Y2=1.825
cc_372 N_VDD_c_360_p N_Q_c_1795_n 0.00736239f $X=9.175 $Y=4.22 $X2=0.53
+ $Y2=1.825
cc_373 N_VDD_M1004_b N_Q_c_1793_n 0.0127419f $X=-0.05 $Y=2.425 $X2=0.32 $Y2=2.85
cc_374 N_VDD_M1004_b Q 0.0106945f $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_375 N_VDD_c_335_p Q 0.00675808f $X=8.85 $Y=3.265 $X2=0 $Y2=0
cc_376 N_VDD_M1004_b N_Q_c_1802_n 0.0190821f $X=-0.05 $Y=2.425 $X2=0 $Y2=0
cc_377 N_VDD_c_335_p N_Q_c_1802_n 0.00905719f $X=8.85 $Y=3.265 $X2=0 $Y2=0
cc_378 RN N_A_110_115#_M1004_d 0.00410657f $X=0.325 $Y=2.85 $X2=1.085 $Y2=0.575
cc_379 N_RN_c_383_n N_A_110_115#_M1015_g 0.00315143f $X=0.475 $Y=1.99 $X2=0
+ $Y2=0
cc_380 N_RN_M1004_g N_A_110_115#_c_432_n 0.00968001f $X=0.475 $Y=3.235 $X2=0
+ $Y2=0
cc_381 N_RN_c_386_n N_A_110_115#_c_432_n 0.0281933f $X=0.32 $Y=2.85 $X2=0 $Y2=0
cc_382 RN N_A_110_115#_c_432_n 0.0097626f $X=0.325 $Y=2.85 $X2=0 $Y2=0
cc_383 N_RN_M1021_g N_A_110_115#_c_433_n 0.0107733f $X=0.475 $Y=0.835 $X2=0
+ $Y2=0
cc_384 N_RN_c_383_n N_A_110_115#_c_433_n 0.00370757f $X=0.475 $Y=1.99 $X2=0
+ $Y2=0
cc_385 N_RN_M1004_g N_A_110_115#_c_433_n 0.00363549f $X=0.475 $Y=3.235 $X2=0
+ $Y2=0
cc_386 N_RN_c_385_n N_A_110_115#_c_433_n 0.0248372f $X=0.32 $Y=1.825 $X2=0 $Y2=0
cc_387 N_RN_c_386_n N_A_110_115#_c_433_n 0.0072511f $X=0.32 $Y=2.85 $X2=0 $Y2=0
cc_388 N_RN_M1021_g N_A_110_115#_c_436_n 0.0067448f $X=0.475 $Y=0.835 $X2=0
+ $Y2=0
cc_389 N_RN_c_383_n N_A_110_115#_c_436_n 0.00166615f $X=0.475 $Y=1.99 $X2=0
+ $Y2=0
cc_390 N_RN_c_385_n N_A_110_115#_c_436_n 3.95917e-19 $X=0.32 $Y=1.825 $X2=0
+ $Y2=0
cc_391 N_RN_c_383_n N_A_110_115#_c_437_n 0.00191737f $X=0.475 $Y=1.99 $X2=0
+ $Y2=0
cc_392 N_RN_M1004_g N_A_110_115#_c_437_n 0.00385986f $X=0.475 $Y=3.235 $X2=0
+ $Y2=0
cc_393 N_RN_c_385_n N_A_110_115#_c_437_n 7.08415e-19 $X=0.32 $Y=1.825 $X2=0
+ $Y2=0
cc_394 N_RN_c_386_n N_A_110_115#_c_437_n 0.0113366f $X=0.32 $Y=2.85 $X2=0 $Y2=0
cc_395 N_RN_M1021_g N_A_110_115#_c_466_n 0.00524963f $X=0.475 $Y=0.835 $X2=0
+ $Y2=0
cc_396 N_RN_M1004_g N_A_217_605#_c_1010_n 0.0035258f $X=0.475 $Y=3.235 $X2=0
+ $Y2=0
cc_397 RN N_A_217_605#_c_1010_n 8.83853e-19 $X=0.325 $Y=2.85 $X2=0 $Y2=0
cc_398 N_A_110_115#_c_438_n N_A_342_442#_M1031_d 0.0032387f $X=7.805 $Y=1
+ $X2=0.135 $Y2=0.575
cc_399 N_A_110_115#_c_416_n N_A_342_442#_M1005_g 0.0597799f $X=1.425 $Y=1.045
+ $X2=0 $Y2=0
cc_400 N_A_110_115#_c_438_n N_A_342_442#_M1005_g 0.00770937f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_401 N_A_110_115#_c_438_n N_A_342_442#_c_619_n 0.0257941f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_402 N_A_110_115#_c_438_n N_A_342_442#_c_621_n 0.00300956f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_403 N_A_110_115#_c_438_n N_A_342_442#_c_623_n 0.0151351f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_404 N_A_110_115#_M1015_g N_A_342_442#_c_624_n 9.08764e-19 $X=1.425 $Y=3.445
+ $X2=0 $Y2=0
cc_405 N_A_110_115#_M1015_g N_A_342_442#_c_625_n 0.106726f $X=1.425 $Y=3.445
+ $X2=0 $Y2=0
cc_406 N_A_110_115#_c_438_n N_A_342_442#_c_626_n 0.0133869f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_407 N_A_110_115#_c_438_n N_D_M1007_g 0.00683925f $X=7.805 $Y=1 $X2=1.93
+ $Y2=0.575
cc_408 N_A_110_115#_c_438_n N_A_618_424#_M1010_d 0.00357716f $X=7.805 $Y=1
+ $X2=0.135 $Y2=0.575
cc_409 N_A_110_115#_c_438_n N_A_618_424#_c_740_n 0.00493929f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_410 N_A_110_115#_c_438_n N_A_618_424#_c_741_n 8.06574e-19 $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_411 N_A_110_115#_c_438_n N_A_618_424#_c_742_n 0.00493657f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_412 N_A_110_115#_c_438_n N_A_618_424#_c_743_n 8.06574e-19 $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_413 N_A_110_115#_c_438_n N_A_618_424#_c_746_n 0.0167515f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_414 N_A_110_115#_c_438_n N_A_618_424#_c_749_n 0.0144841f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_415 N_A_110_115#_c_438_n N_A_618_424#_c_763_n 0.0064255f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_416 N_A_110_115#_c_438_n N_A_618_424#_c_766_n 0.00633231f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_417 N_A_110_115#_c_438_n N_A_217_605#_M1018_d 0.00142852f $X=7.805 $Y=1
+ $X2=0.135 $Y2=0.575
cc_418 N_A_110_115#_c_438_n N_A_217_605#_M1027_g 0.00607163f $X=7.805 $Y=1
+ $X2=8.71 $Y2=0.575
cc_419 N_A_110_115#_c_438_n N_A_217_605#_M1025_g 0.00632589f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_420 N_A_110_115#_c_438_n N_A_217_605#_c_1007_n 2.42482e-19 $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_421 N_A_110_115#_M1015_g N_A_217_605#_c_1010_n 0.0409873f $X=1.425 $Y=3.445
+ $X2=0 $Y2=0
cc_422 N_A_110_115#_c_432_n N_A_217_605#_c_1010_n 0.0652498f $X=0.69 $Y=2.95
+ $X2=0 $Y2=0
cc_423 N_A_110_115#_c_433_n N_A_217_605#_c_1010_n 0.0210459f $X=0.87 $Y=2.175
+ $X2=0 $Y2=0
cc_424 N_A_110_115#_c_437_n N_A_217_605#_c_1010_n 0.0134441f $X=0.87 $Y=2.26
+ $X2=0 $Y2=0
cc_425 N_A_110_115#_M1015_g N_A_217_605#_c_1011_n 0.0188678f $X=1.425 $Y=3.445
+ $X2=0 $Y2=0
cc_426 N_A_110_115#_c_462_n N_A_217_605#_c_1011_n 0.00181457f $X=1.22 $Y=1.37
+ $X2=0 $Y2=0
cc_427 N_A_110_115#_c_464_n N_A_217_605#_c_1011_n 0.00235169f $X=1.22 $Y=1.21
+ $X2=0 $Y2=0
cc_428 N_A_110_115#_c_466_n N_A_217_605#_c_1011_n 6.98912e-19 $X=1.425 $Y=1.21
+ $X2=0 $Y2=0
cc_429 N_A_110_115#_c_433_n N_A_217_605#_c_1012_n 0.0142099f $X=0.87 $Y=2.175
+ $X2=0 $Y2=0
cc_430 N_A_110_115#_c_434_n N_A_217_605#_c_1012_n 2.13728e-19 $X=1.135 $Y=1.21
+ $X2=0 $Y2=0
cc_431 N_A_110_115#_c_462_n N_A_217_605#_c_1012_n 0.00574122f $X=1.22 $Y=1.37
+ $X2=0 $Y2=0
cc_432 N_A_110_115#_c_464_n N_A_217_605#_c_1012_n 0.00732624f $X=1.22 $Y=1.21
+ $X2=0 $Y2=0
cc_433 N_A_110_115#_c_466_n N_A_217_605#_c_1012_n 0.00117358f $X=1.425 $Y=1.21
+ $X2=0 $Y2=0
cc_434 N_A_110_115#_c_438_n N_A_217_605#_c_1014_n 0.184203f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_435 N_A_110_115#_M1015_g N_A_217_605#_c_1015_n 0.00152013f $X=1.425 $Y=3.445
+ $X2=0 $Y2=0
cc_436 N_A_110_115#_c_536_p N_A_217_605#_c_1015_n 3.8078e-19 $X=1.22 $Y=1.255
+ $X2=0 $Y2=0
cc_437 N_A_110_115#_c_438_n N_A_217_605#_c_1015_n 0.0254104f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_438 N_A_110_115#_c_462_n N_A_217_605#_c_1015_n 0.0252399f $X=1.22 $Y=1.37
+ $X2=0 $Y2=0
cc_439 N_A_110_115#_c_464_n N_A_217_605#_c_1015_n 9.3821e-19 $X=1.22 $Y=1.21
+ $X2=0 $Y2=0
cc_440 N_A_110_115#_c_466_n N_A_217_605#_c_1015_n 0.0015251f $X=1.425 $Y=1.21
+ $X2=0 $Y2=0
cc_441 N_A_110_115#_c_438_n N_A_217_605#_c_1061_n 0.0259207f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_442 N_A_110_115#_c_438_n N_A_217_605#_c_1016_n 0.00476535f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_443 N_A_110_115#_c_416_n N_A_217_605#_c_1018_n 0.00886891f $X=1.425 $Y=1.045
+ $X2=0 $Y2=0
cc_444 N_A_110_115#_c_433_n N_A_217_605#_c_1018_n 0.00730421f $X=0.87 $Y=2.175
+ $X2=0 $Y2=0
cc_445 N_A_110_115#_c_436_n N_A_217_605#_c_1018_n 0.00143173f $X=0.955 $Y=1.21
+ $X2=0 $Y2=0
cc_446 N_A_110_115#_c_536_p N_A_217_605#_c_1018_n 0.00177859f $X=1.22 $Y=1.255
+ $X2=0 $Y2=0
cc_447 N_A_110_115#_c_438_n N_A_217_605#_c_1018_n 0.0195703f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_448 N_A_110_115#_c_462_n N_A_217_605#_c_1018_n 0.00122345f $X=1.22 $Y=1.37
+ $X2=0 $Y2=0
cc_449 N_A_110_115#_c_464_n N_A_217_605#_c_1018_n 0.0197974f $X=1.22 $Y=1.21
+ $X2=0 $Y2=0
cc_450 N_A_110_115#_c_438_n N_CK_c_1135_n 0.00599689f $X=7.805 $Y=1 $X2=0.135
+ $Y2=0.575
cc_451 N_A_110_115#_c_438_n N_CK_M1020_g 0.00631256f $X=7.805 $Y=1 $X2=0 $Y2=0
cc_452 N_A_110_115#_c_438_n N_CK_c_1148_n 0.00702161f $X=7.805 $Y=1 $X2=0 $Y2=0
cc_453 N_A_110_115#_c_438_n N_CK_c_1158_n 0.00157179f $X=7.805 $Y=1 $X2=0 $Y2=0
cc_454 N_A_110_115#_c_438_n N_A_1160_89#_M1012_d 0.00142852f $X=7.805 $Y=1
+ $X2=0.135 $Y2=0.575
cc_455 N_A_110_115#_c_421_n N_A_1160_89#_M1016_g 0.00187137f $X=7.615 $Y=1.52
+ $X2=0 $Y2=0
cc_456 N_A_110_115#_c_438_n N_A_1160_89#_c_1345_n 0.00599085f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_457 N_A_110_115#_c_438_n N_A_1160_89#_c_1349_n 5.89421e-19 $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_458 N_A_110_115#_c_421_n N_A_1160_89#_c_1352_n 0.00416492f $X=7.615 $Y=1.52
+ $X2=0 $Y2=0
cc_459 N_A_110_115#_c_468_n N_A_1160_89#_c_1352_n 4.20096e-19 $X=7.89 $Y=1.21
+ $X2=0 $Y2=0
cc_460 N_A_110_115#_M1030_g N_A_1160_89#_c_1388_n 0.00633587f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_461 N_A_110_115#_c_421_n N_A_1160_89#_c_1355_n 0.00411162f $X=7.615 $Y=1.52
+ $X2=0 $Y2=0
cc_462 N_A_110_115#_M1030_g N_A_1160_89#_c_1355_n 0.00587172f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_463 N_A_110_115#_c_424_n N_A_1160_89#_c_1355_n 0.00633298f $X=7.685 $Y=1.045
+ $X2=0 $Y2=0
cc_464 N_A_110_115#_c_438_n N_A_1160_89#_c_1355_n 0.0249056f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_465 N_A_110_115#_c_565_p N_A_1160_89#_c_1355_n 0.00235259f $X=7.89 $Y=1.255
+ $X2=0 $Y2=0
cc_466 N_A_110_115#_c_463_n N_A_1160_89#_c_1355_n 0.00272511f $X=7.89 $Y=1.37
+ $X2=0 $Y2=0
cc_467 N_A_110_115#_c_468_n N_A_1160_89#_c_1355_n 0.0183071f $X=7.89 $Y=1.21
+ $X2=0 $Y2=0
cc_468 N_A_110_115#_M1030_g N_A_1160_89#_c_1358_n 0.0483827f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_469 N_A_110_115#_M1030_g N_A_1160_89#_c_1363_n 0.00122231f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_470 N_A_110_115#_c_421_n N_A_1160_89#_c_1370_n 0.00465519f $X=7.615 $Y=1.52
+ $X2=0 $Y2=0
cc_471 N_A_110_115#_M1030_g N_A_1160_89#_c_1370_n 0.0118805f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_472 N_A_110_115#_c_438_n N_A_1160_89#_c_1370_n 0.00335122f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_473 N_A_110_115#_c_463_n N_A_1160_89#_c_1370_n 0.00122291f $X=7.89 $Y=1.37
+ $X2=0 $Y2=0
cc_474 N_A_110_115#_c_468_n N_A_1160_89#_c_1370_n 0.0151944f $X=7.89 $Y=1.21
+ $X2=0 $Y2=0
cc_475 N_A_110_115#_c_421_n N_A_1160_89#_c_1371_n 0.00234211f $X=7.615 $Y=1.52
+ $X2=0 $Y2=0
cc_476 N_A_110_115#_M1030_g N_A_1160_89#_c_1371_n 0.0111655f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_477 N_A_110_115#_c_463_n N_A_1160_89#_c_1371_n 0.028449f $X=7.89 $Y=1.37
+ $X2=0 $Y2=0
cc_478 N_A_110_115#_c_468_n N_A_1160_89#_c_1371_n 0.00196064f $X=7.89 $Y=1.21
+ $X2=0 $Y2=0
cc_479 N_A_110_115#_M1030_g N_A_1160_89#_c_1373_n 0.00507506f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_480 N_A_110_115#_c_463_n N_A_1160_89#_c_1374_n 6.06666e-19 $X=7.89 $Y=1.37
+ $X2=0 $Y2=0
cc_481 N_A_110_115#_c_468_n N_A_1160_89#_c_1374_n 2.80323e-19 $X=7.89 $Y=1.21
+ $X2=0 $Y2=0
cc_482 N_A_110_115#_c_438_n N_A_998_115#_M1019_d 0.0032738f $X=7.805 $Y=1
+ $X2=0.135 $Y2=0.575
cc_483 N_A_110_115#_c_424_n N_A_998_115#_M1012_g 0.0122299f $X=7.685 $Y=1.045
+ $X2=8.71 $Y2=0.575
cc_484 N_A_110_115#_c_438_n N_A_998_115#_M1012_g 0.0119892f $X=7.805 $Y=1
+ $X2=8.71 $Y2=0.575
cc_485 N_A_110_115#_M1030_g N_A_998_115#_M1006_g 0.0812648f $X=7.615 $Y=3.445
+ $X2=0 $Y2=0
cc_486 N_A_110_115#_c_438_n N_A_998_115#_c_1554_n 0.0230872f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_487 N_A_110_115#_c_438_n N_A_998_115#_c_1557_n 0.0328521f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_488 N_A_110_115#_c_438_n N_A_998_115#_c_1558_n 0.0259499f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_489 N_A_110_115#_c_438_n N_A_998_115#_c_1559_n 0.122091f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_490 N_A_110_115#_c_438_n N_A_998_115#_c_1561_n 0.0224792f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_491 N_A_110_115#_c_438_n N_A_998_115#_c_1562_n 0.00554379f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_492 N_A_110_115#_c_438_n N_A_998_115#_c_1563_n 0.00648735f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_493 N_A_110_115#_c_438_n N_A_998_115#_c_1564_n 0.0260564f $X=7.805 $Y=1 $X2=0
+ $Y2=0
cc_494 N_A_110_115#_c_463_n N_A_998_115#_c_1564_n 0.011315f $X=7.89 $Y=1.37
+ $X2=0 $Y2=0
cc_495 N_A_110_115#_c_438_n N_A_998_115#_c_1565_n 0.00160369f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_496 N_A_110_115#_c_421_n N_A_998_115#_c_1567_n 0.0934947f $X=7.615 $Y=1.52
+ $X2=0 $Y2=0
cc_497 N_A_110_115#_c_438_n N_A_998_115#_c_1567_n 0.00151039f $X=7.805 $Y=1
+ $X2=0 $Y2=0
cc_498 N_A_110_115#_c_421_n N_QN_c_1700_n 0.00222227f $X=7.615 $Y=1.52 $X2=0
+ $Y2=0
cc_499 N_A_110_115#_c_424_n N_QN_c_1700_n 0.00298655f $X=7.685 $Y=1.045 $X2=0
+ $Y2=0
cc_500 N_A_110_115#_c_438_n N_QN_c_1700_n 0.00875851f $X=7.805 $Y=1 $X2=0 $Y2=0
cc_501 N_A_110_115#_c_565_p N_QN_c_1700_n 7.96604e-19 $X=7.89 $Y=1.255 $X2=0
+ $Y2=0
cc_502 N_A_110_115#_c_463_n N_QN_c_1700_n 2.00168e-19 $X=7.89 $Y=1.37 $X2=0
+ $Y2=0
cc_503 N_A_110_115#_c_468_n N_QN_c_1700_n 0.00781846f $X=7.89 $Y=1.21 $X2=0
+ $Y2=0
cc_504 N_A_110_115#_c_421_n N_QN_c_1706_n 6.86262e-19 $X=7.615 $Y=1.52 $X2=0
+ $Y2=0
cc_505 N_A_110_115#_c_463_n N_QN_c_1706_n 0.00464864f $X=7.89 $Y=1.37 $X2=0
+ $Y2=0
cc_506 N_A_110_115#_c_468_n N_QN_c_1706_n 0.00565014f $X=7.89 $Y=1.21 $X2=0
+ $Y2=0
cc_507 N_A_110_115#_M1030_g N_QN_c_1708_n 0.00423893f $X=7.615 $Y=3.445 $X2=0
+ $Y2=0
cc_508 N_A_110_115#_M1030_g N_QN_c_1711_n 0.0144714f $X=7.615 $Y=3.445 $X2=0
+ $Y2=0
cc_509 N_A_110_115#_M1030_g QN 0.00472165f $X=7.615 $Y=3.445 $X2=0 $Y2=0
cc_510 N_A_110_115#_c_438_n A_576_115# 0.00381028f $X=7.805 $Y=1 $X2=0.135
+ $Y2=0.575
cc_511 N_A_110_115#_c_438_n A_768_115# 0.00473401f $X=7.805 $Y=1 $X2=0.135
+ $Y2=0.575
cc_512 N_A_110_115#_c_438_n A_926_115# 0.00429254f $X=7.805 $Y=1 $X2=0.135
+ $Y2=0.575
cc_513 N_A_110_115#_c_438_n A_1118_115# 0.00465218f $X=7.805 $Y=1 $X2=0.135
+ $Y2=0.575
cc_514 N_A_342_442#_c_618_n N_D_M1007_g 0.0137346f $X=2.11 $Y=2.21 $X2=1.93
+ $Y2=0.575
cc_515 N_A_342_442#_c_619_n N_D_M1007_g 0.0122665f $X=3.28 $Y=1.285 $X2=1.93
+ $Y2=0.575
cc_516 N_A_342_442#_c_621_n N_D_M1007_g 0.00158134f $X=2.2 $Y=1.285 $X2=1.93
+ $Y2=0.575
cc_517 N_A_342_442#_c_633_n N_D_M1028_g 0.0211478f $X=3.295 $Y=2.705 $X2=6.915
+ $Y2=0.575
cc_518 N_A_342_442#_c_624_n N_D_M1028_g 0.00767395f $X=1.94 $Y=2.375 $X2=6.915
+ $Y2=0.575
cc_519 N_A_342_442#_c_625_n N_D_M1028_g 0.00395324f $X=1.94 $Y=2.375 $X2=6.915
+ $Y2=0.575
cc_520 N_A_342_442#_c_618_n D 0.0055149f $X=2.11 $Y=2.21 $X2=0 $Y2=0
cc_521 N_A_342_442#_c_619_n D 0.00200799f $X=3.28 $Y=1.285 $X2=0 $Y2=0
cc_522 N_A_342_442#_c_618_n N_D_c_703_n 0.00613892f $X=2.11 $Y=2.21 $X2=0 $Y2=0
cc_523 N_A_342_442#_c_619_n N_D_c_703_n 0.0086486f $X=3.28 $Y=1.285 $X2=0 $Y2=0
cc_524 N_A_342_442#_c_619_n N_D_c_704_n 0.00207628f $X=3.28 $Y=1.285 $X2=0 $Y2=0
cc_525 N_A_342_442#_c_633_n N_A_618_424#_M1024_g 0.0153421f $X=3.295 $Y=2.705
+ $X2=8.71 $Y2=0.575
cc_526 N_A_342_442#_c_633_n N_A_618_424#_c_739_n 0.00883015f $X=3.295 $Y=2.705
+ $X2=0 $Y2=0
cc_527 N_A_342_442#_c_619_n N_A_618_424#_c_739_n 0.0019742f $X=3.28 $Y=1.285
+ $X2=0 $Y2=0
cc_528 N_A_342_442#_c_619_n N_A_618_424#_c_740_n 0.012316f $X=3.28 $Y=1.285
+ $X2=0 $Y2=0
cc_529 N_A_342_442#_c_626_n N_A_618_424#_c_740_n 5.6626e-19 $X=3.365 $Y=0.755
+ $X2=0 $Y2=0
cc_530 N_A_342_442#_c_619_n N_A_618_424#_c_741_n 9.45214e-19 $X=3.28 $Y=1.285
+ $X2=0 $Y2=0
cc_531 N_A_342_442#_c_626_n N_A_618_424#_c_741_n 0.00165184f $X=3.365 $Y=0.755
+ $X2=0 $Y2=0
cc_532 N_A_342_442#_c_633_n N_A_618_424#_c_754_n 0.00601583f $X=3.295 $Y=2.705
+ $X2=0 $Y2=0
cc_533 N_A_342_442#_c_633_n N_A_618_424#_c_755_n 0.00409373f $X=3.295 $Y=2.705
+ $X2=0 $Y2=0
cc_534 N_A_342_442#_c_633_n N_A_618_424#_c_758_n 0.0101098f $X=3.295 $Y=2.705
+ $X2=0 $Y2=0
cc_535 N_A_342_442#_c_619_n N_A_618_424#_c_758_n 0.00224443f $X=3.28 $Y=1.285
+ $X2=0 $Y2=0
cc_536 N_A_342_442#_c_633_n N_A_618_424#_c_762_n 0.00150627f $X=3.295 $Y=2.705
+ $X2=0 $Y2=0
cc_537 N_A_342_442#_c_623_n N_A_618_424#_c_763_n 0.00464203f $X=3.365 $Y=1.2
+ $X2=0 $Y2=0
cc_538 N_A_342_442#_c_626_n N_A_618_424#_c_763_n 0.00243799f $X=3.365 $Y=0.755
+ $X2=0 $Y2=0
cc_539 N_A_342_442#_c_624_n N_A_217_605#_c_1010_n 0.0100421f $X=1.94 $Y=2.375
+ $X2=0 $Y2=0
cc_540 N_A_342_442#_M1005_g N_A_217_605#_c_1011_n 0.00176497f $X=1.855 $Y=0.755
+ $X2=0 $Y2=0
cc_541 N_A_342_442#_c_618_n N_A_217_605#_c_1011_n 0.00954176f $X=2.11 $Y=2.21
+ $X2=0 $Y2=0
cc_542 N_A_342_442#_c_625_n N_A_217_605#_c_1011_n 6.21732e-19 $X=1.94 $Y=2.375
+ $X2=0 $Y2=0
cc_543 N_A_342_442#_M1005_g N_A_217_605#_c_1014_n 0.0112415f $X=1.855 $Y=0.755
+ $X2=0 $Y2=0
cc_544 N_A_342_442#_c_619_n N_A_217_605#_c_1014_n 0.0476148f $X=3.28 $Y=1.285
+ $X2=0 $Y2=0
cc_545 N_A_342_442#_c_621_n N_A_217_605#_c_1014_n 0.0198865f $X=2.2 $Y=1.285
+ $X2=0 $Y2=0
cc_546 N_A_342_442#_c_626_n N_A_217_605#_c_1014_n 8.84066e-19 $X=3.365 $Y=0.755
+ $X2=0 $Y2=0
cc_547 N_A_342_442#_M1005_g N_A_217_605#_c_1015_n 0.00236248f $X=1.855 $Y=0.755
+ $X2=0 $Y2=0
cc_548 N_A_342_442#_c_618_n N_A_217_605#_c_1015_n 6.00227e-19 $X=2.11 $Y=2.21
+ $X2=0 $Y2=0
cc_549 N_A_342_442#_c_621_n N_A_217_605#_c_1015_n 0.00125688f $X=2.2 $Y=1.285
+ $X2=0 $Y2=0
cc_550 N_A_342_442#_M1005_g N_A_217_605#_c_1018_n 0.0102637f $X=1.855 $Y=0.755
+ $X2=0 $Y2=0
cc_551 N_A_342_442#_c_618_n N_A_217_605#_c_1018_n 0.012524f $X=2.11 $Y=2.21
+ $X2=0 $Y2=0
cc_552 N_A_342_442#_c_621_n N_A_217_605#_c_1018_n 0.011766f $X=2.2 $Y=1.285
+ $X2=0 $Y2=0
cc_553 N_A_342_442#_c_619_n N_CK_c_1135_n 0.0022787f $X=3.28 $Y=1.285 $X2=0.135
+ $Y2=0.575
cc_554 N_A_342_442#_c_623_n N_CK_c_1135_n 0.00492892f $X=3.365 $Y=1.2 $X2=0.135
+ $Y2=0.575
cc_555 N_A_342_442#_c_626_n N_CK_c_1135_n 0.00116801f $X=3.365 $Y=0.755
+ $X2=0.135 $Y2=0.575
cc_556 N_A_342_442#_c_619_n N_CK_c_1138_n 0.00326059f $X=3.28 $Y=1.285 $X2=4.2
+ $Y2=0.575
cc_557 N_A_342_442#_c_619_n N_CK_c_1155_n 0.00984832f $X=3.28 $Y=1.285 $X2=0
+ $Y2=0
cc_558 N_A_342_442#_c_633_n A_576_521# 0.00732587f $X=3.295 $Y=2.705 $X2=0.135
+ $Y2=0.575
cc_559 D N_A_618_424#_c_740_n 0.00551577f $X=2.865 $Y=1.74 $X2=0 $Y2=0
cc_560 N_D_c_703_n N_A_618_424#_c_740_n 0.00478177f $X=2.865 $Y=1.74 $X2=0 $Y2=0
cc_561 N_D_c_704_n N_A_618_424#_c_740_n 2.89615e-19 $X=2.865 $Y=1.74 $X2=0 $Y2=0
cc_562 N_D_M1028_g N_A_618_424#_c_755_n 0.00515433f $X=2.805 $Y=3.235 $X2=0
+ $Y2=0
cc_563 D N_A_618_424#_c_755_n 0.00375733f $X=2.865 $Y=1.74 $X2=0 $Y2=0
cc_564 N_D_M1028_g N_A_618_424#_c_758_n 0.00494364f $X=2.805 $Y=3.235 $X2=0
+ $Y2=0
cc_565 N_D_M1028_g N_A_618_424#_c_762_n 0.11474f $X=2.805 $Y=3.235 $X2=0 $Y2=0
cc_566 N_D_M1007_g N_A_217_605#_c_1014_n 0.0030176f $X=2.805 $Y=0.835 $X2=0
+ $Y2=0
cc_567 D N_A_217_605#_c_1014_n 0.0353362f $X=2.865 $Y=1.74 $X2=0 $Y2=0
cc_568 N_D_c_703_n N_A_217_605#_c_1014_n 0.00111625f $X=2.865 $Y=1.74 $X2=0
+ $Y2=0
cc_569 N_D_c_704_n N_A_217_605#_c_1014_n 7.9412e-19 $X=2.865 $Y=1.74 $X2=0 $Y2=0
cc_570 N_D_M1007_g N_CK_c_1135_n 0.0567053f $X=2.805 $Y=0.835 $X2=0.135
+ $Y2=0.575
cc_571 N_D_M1007_g N_CK_c_1138_n 0.00932846f $X=2.805 $Y=0.835 $X2=4.2 $Y2=0.575
cc_572 D N_CK_c_1138_n 0.00342011f $X=2.865 $Y=1.74 $X2=4.2 $Y2=0.575
cc_573 N_D_c_703_n N_CK_c_1138_n 0.00164409f $X=2.865 $Y=1.74 $X2=4.2 $Y2=0.575
cc_574 N_D_c_704_n N_CK_c_1138_n 0.0210215f $X=2.865 $Y=1.74 $X2=4.2 $Y2=0.575
cc_575 D N_CK_c_1140_n 4.62757e-19 $X=2.865 $Y=1.74 $X2=6.915 $Y2=0.575
cc_576 N_A_618_424#_c_740_n N_A_217_605#_M1027_g 0.00109079f $X=3.705 $Y=1.37
+ $X2=8.71 $Y2=0.575
cc_577 N_A_618_424#_c_763_n N_A_217_605#_M1027_g 0.0338208f $X=3.705 $Y=1.205
+ $X2=8.71 $Y2=0.575
cc_578 N_A_618_424#_c_742_n N_A_217_605#_M1025_g 3.67139e-19 $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_579 N_A_618_424#_c_766_n N_A_217_605#_M1025_g 0.0333732f $X=4.975 $Y=1.205
+ $X2=0 $Y2=0
cc_580 N_A_618_424#_c_741_n N_A_217_605#_c_1005_n 0.0338208f $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_581 N_A_618_424#_c_754_n N_A_217_605#_c_1006_n 0.00679967f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_582 N_A_618_424#_c_743_n N_A_217_605#_c_1007_n 0.0333732f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_583 N_A_618_424#_c_754_n N_A_217_605#_c_1009_n 0.00772879f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_584 N_A_618_424#_c_739_n N_A_217_605#_c_1013_n 0.00401809f $X=3.62 $Y=2.11
+ $X2=0 $Y2=0
cc_585 N_A_618_424#_c_740_n N_A_217_605#_c_1013_n 0.0203851f $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_586 N_A_618_424#_c_741_n N_A_217_605#_c_1013_n 7.30049e-19 $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_587 N_A_618_424#_c_754_n N_A_217_605#_c_1013_n 0.0206884f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_588 N_A_618_424#_c_739_n N_A_217_605#_c_1014_n 0.00443421f $X=3.62 $Y=2.11
+ $X2=0 $Y2=0
cc_589 N_A_618_424#_c_740_n N_A_217_605#_c_1014_n 0.0149971f $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_590 N_A_618_424#_c_741_n N_A_217_605#_c_1014_n 0.00383172f $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_591 N_A_618_424#_c_755_n N_A_217_605#_c_1014_n 0.0126164f $X=3.37 $Y=2.11
+ $X2=0 $Y2=0
cc_592 N_A_618_424#_c_758_n N_A_217_605#_c_1014_n 7.12046e-19 $X=3.225 $Y=2.11
+ $X2=0 $Y2=0
cc_593 N_A_618_424#_c_740_n N_A_217_605#_c_1061_n 0.00143592f $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_594 N_A_618_424#_c_741_n N_A_217_605#_c_1061_n 3.3031e-19 $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_595 N_A_618_424#_c_754_n N_A_217_605#_c_1061_n 0.0129652f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_596 N_A_618_424#_c_740_n N_A_217_605#_c_1016_n 0.00742068f $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_597 N_A_618_424#_c_741_n N_A_217_605#_c_1016_n 7.18106e-19 $X=3.705 $Y=1.37
+ $X2=0 $Y2=0
cc_598 N_A_618_424#_c_754_n N_A_217_605#_c_1016_n 0.00102309f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_599 N_A_618_424#_c_763_n N_CK_c_1135_n 0.0171207f $X=3.705 $Y=1.205 $X2=0.135
+ $Y2=0.575
cc_600 N_A_618_424#_c_740_n N_CK_c_1138_n 0.00613747f $X=3.705 $Y=1.37 $X2=4.2
+ $Y2=0.575
cc_601 N_A_618_424#_c_740_n N_CK_c_1139_n 0.00630484f $X=3.705 $Y=1.37 $X2=5.95
+ $Y2=0.575
cc_602 N_A_618_424#_c_741_n N_CK_c_1139_n 0.0183603f $X=3.705 $Y=1.37 $X2=5.95
+ $Y2=0.575
cc_603 N_A_618_424#_c_754_n N_CK_c_1139_n 0.00613485f $X=5.31 $Y=2.11 $X2=5.95
+ $Y2=0.575
cc_604 N_A_618_424#_c_739_n N_CK_c_1140_n 0.00878348f $X=3.62 $Y=2.11 $X2=6.915
+ $Y2=0.575
cc_605 N_A_618_424#_c_755_n N_CK_c_1140_n 0.00137501f $X=3.37 $Y=2.11 $X2=6.915
+ $Y2=0.575
cc_606 N_A_618_424#_c_758_n N_CK_c_1140_n 0.00109468f $X=3.225 $Y=2.11 $X2=6.915
+ $Y2=0.575
cc_607 N_A_618_424#_c_762_n N_CK_c_1140_n 0.00904036f $X=3.225 $Y=2.285
+ $X2=6.915 $Y2=0.575
cc_608 N_A_618_424#_M1024_g N_CK_M1017_g 0.0316011f $X=3.165 $Y=3.235 $X2=0
+ $Y2=0
cc_609 N_A_618_424#_c_739_n N_CK_M1017_g 0.0081071f $X=3.62 $Y=2.11 $X2=0 $Y2=0
cc_610 N_A_618_424#_c_740_n N_CK_M1017_g 0.00478024f $X=3.705 $Y=1.37 $X2=0
+ $Y2=0
cc_611 N_A_618_424#_c_754_n N_CK_M1017_g 0.00938974f $X=5.31 $Y=2.11 $X2=0 $Y2=0
cc_612 N_A_618_424#_c_755_n N_CK_M1017_g 4.2e-19 $X=3.37 $Y=2.11 $X2=0 $Y2=0
cc_613 N_A_618_424#_c_758_n N_CK_M1017_g 0.00184124f $X=3.225 $Y=2.11 $X2=0
+ $Y2=0
cc_614 N_A_618_424#_c_762_n N_CK_M1017_g 0.0128384f $X=3.225 $Y=2.285 $X2=0
+ $Y2=0
cc_615 N_A_618_424#_c_754_n N_CK_c_1142_n 0.00607908f $X=5.31 $Y=2.11 $X2=0
+ $Y2=0
cc_616 N_A_618_424#_M1000_g N_CK_M1003_g 0.0316011f $X=5.515 $Y=3.235 $X2=0
+ $Y2=0
cc_617 N_A_618_424#_c_742_n N_CK_M1003_g 0.00399495f $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_618 N_A_618_424#_c_745_n N_CK_M1003_g 0.00654233f $X=5.06 $Y=2.11 $X2=0 $Y2=0
cc_619 N_A_618_424#_c_754_n N_CK_M1003_g 0.00497421f $X=5.31 $Y=2.11 $X2=0 $Y2=0
cc_620 N_A_618_424#_c_757_n N_CK_M1003_g 4.2e-19 $X=5.6 $Y=2.11 $X2=0 $Y2=0
cc_621 N_A_618_424#_c_759_n N_CK_M1003_g 0.00128351f $X=5.455 $Y=2.11 $X2=0
+ $Y2=0
cc_622 N_A_618_424#_c_769_n N_CK_M1003_g 0.0118393f $X=5.455 $Y=2.285 $X2=0
+ $Y2=0
cc_623 N_A_618_424#_c_742_n N_CK_c_1144_n 0.00635358f $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_624 N_A_618_424#_c_744_n N_CK_c_1144_n 0.00842176f $X=5.37 $Y=2.11 $X2=0
+ $Y2=0
cc_625 N_A_618_424#_c_754_n N_CK_c_1144_n 0.00519056f $X=5.31 $Y=2.11 $X2=0
+ $Y2=0
cc_626 N_A_618_424#_c_757_n N_CK_c_1144_n 0.00150125f $X=5.6 $Y=2.11 $X2=0 $Y2=0
cc_627 N_A_618_424#_c_742_n N_CK_M1020_g 4.67639e-19 $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_628 N_A_618_424#_c_743_n N_CK_M1020_g 0.012357f $X=4.975 $Y=1.37 $X2=0 $Y2=0
cc_629 N_A_618_424#_c_766_n N_CK_M1020_g 0.017109f $X=4.975 $Y=1.205 $X2=0 $Y2=0
cc_630 N_A_618_424#_c_746_n N_CK_c_1148_n 0.00770147f $X=6.69 $Y=1.76 $X2=0
+ $Y2=0
cc_631 N_A_618_424#_c_749_n N_CK_c_1148_n 0.00275877f $X=6.69 $Y=0.755 $X2=0
+ $Y2=0
cc_632 N_A_618_424#_c_871_p N_CK_c_1153_n 0.00377332f $X=6.605 $Y=2.705 $X2=0
+ $Y2=0
cc_633 N_A_618_424#_c_756_n N_CK_c_1153_n 0.00215772f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_634 N_A_618_424#_c_760_n N_CK_c_1153_n 5.55731e-19 $X=6.87 $Y=2.11 $X2=0
+ $Y2=0
cc_635 N_A_618_424#_c_761_n N_CK_c_1153_n 0.00297273f $X=6.87 $Y=2.11 $X2=0
+ $Y2=0
cc_636 N_A_618_424#_c_761_n N_CK_M1029_g 0.00350595f $X=6.87 $Y=2.11 $X2=0 $Y2=0
cc_637 N_A_618_424#_c_753_n N_CK_c_1154_n 0.00185331f $X=6.87 $Y=1.845 $X2=0
+ $Y2=0
cc_638 N_A_618_424#_c_756_n N_CK_c_1154_n 0.00173153f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_639 N_A_618_424#_c_760_n N_CK_c_1154_n 4.95116e-19 $X=6.87 $Y=2.11 $X2=0
+ $Y2=0
cc_640 N_A_618_424#_c_761_n N_CK_c_1154_n 0.0014377f $X=6.87 $Y=2.11 $X2=0 $Y2=0
cc_641 N_A_618_424#_c_741_n N_CK_c_1155_n 0.0216263f $X=3.705 $Y=1.37 $X2=0
+ $Y2=0
cc_642 N_A_618_424#_c_758_n N_CK_c_1155_n 2.45465e-19 $X=3.225 $Y=2.11 $X2=0
+ $Y2=0
cc_643 N_A_618_424#_c_740_n N_CK_c_1156_n 0.00568091f $X=3.705 $Y=1.37 $X2=0
+ $Y2=0
cc_644 N_A_618_424#_c_742_n N_CK_c_1157_n 0.00436024f $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_645 N_A_618_424#_c_743_n N_CK_c_1157_n 0.0183603f $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_646 N_A_618_424#_c_746_n N_CK_c_1158_n 0.0105063f $X=6.69 $Y=1.76 $X2=0 $Y2=0
cc_647 N_A_618_424#_c_749_n N_CK_c_1158_n 0.00193837f $X=6.69 $Y=0.755 $X2=0
+ $Y2=0
cc_648 N_A_618_424#_c_871_p N_CK_c_1159_n 0.00671583f $X=6.605 $Y=2.705 $X2=0
+ $Y2=0
cc_649 N_A_618_424#_c_756_n N_CK_c_1159_n 0.0115099f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_650 N_A_618_424#_c_760_n N_CK_c_1159_n 8.71161e-19 $X=6.87 $Y=2.11 $X2=0
+ $Y2=0
cc_651 N_A_618_424#_c_761_n N_CK_c_1159_n 0.0161379f $X=6.87 $Y=2.11 $X2=0 $Y2=0
cc_652 N_A_618_424#_c_756_n N_CK_c_1160_n 0.0456907f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_653 N_A_618_424#_c_742_n N_CK_c_1246_n 0.00243046f $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_654 N_A_618_424#_c_757_n N_CK_c_1246_n 0.0296144f $X=5.6 $Y=2.11 $X2=0 $Y2=0
cc_655 N_A_618_424#_c_759_n N_CK_c_1246_n 4.75808e-19 $X=5.455 $Y=2.11 $X2=0
+ $Y2=0
cc_656 N_A_618_424#_c_746_n N_CK_c_1161_n 0.00505303f $X=6.69 $Y=1.76 $X2=0
+ $Y2=0
cc_657 N_A_618_424#_c_753_n N_CK_c_1161_n 0.00953369f $X=6.87 $Y=1.845 $X2=0
+ $Y2=0
cc_658 N_A_618_424#_c_756_n N_CK_c_1161_n 0.00699207f $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_659 N_A_618_424#_c_760_n N_CK_c_1161_n 7.68977e-19 $X=6.87 $Y=2.11 $X2=0
+ $Y2=0
cc_660 N_A_618_424#_c_761_n N_CK_c_1161_n 0.00575856f $X=6.87 $Y=2.11 $X2=0
+ $Y2=0
cc_661 N_A_618_424#_c_746_n CK 0.00414445f $X=6.69 $Y=1.76 $X2=0 $Y2=0
cc_662 N_A_618_424#_c_753_n CK 0.00280277f $X=6.87 $Y=1.845 $X2=0 $Y2=0
cc_663 N_A_618_424#_c_756_n CK 0.0257388f $X=6.725 $Y=2.11 $X2=0 $Y2=0
cc_664 N_A_618_424#_c_742_n N_CK_c_1163_n 0.003871f $X=4.975 $Y=1.37 $X2=0 $Y2=0
cc_665 N_A_618_424#_c_743_n N_CK_c_1163_n 9.99307e-19 $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_666 N_A_618_424#_c_756_n N_CK_c_1163_n 3.23651e-19 $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_667 N_A_618_424#_c_759_n N_CK_c_1163_n 0.0010914f $X=5.455 $Y=2.11 $X2=0
+ $Y2=0
cc_668 N_A_618_424#_c_769_n N_CK_c_1163_n 0.0165037f $X=5.455 $Y=2.285 $X2=0
+ $Y2=0
cc_669 N_A_618_424#_c_742_n N_CK_c_1164_n 0.0107188f $X=4.975 $Y=1.37 $X2=0
+ $Y2=0
cc_670 N_A_618_424#_c_744_n N_CK_c_1164_n 0.00447505f $X=5.37 $Y=2.11 $X2=0
+ $Y2=0
cc_671 N_A_618_424#_c_756_n N_CK_c_1164_n 2.90862e-19 $X=6.725 $Y=2.11 $X2=0
+ $Y2=0
cc_672 N_A_618_424#_c_757_n N_CK_c_1164_n 0.0019318f $X=5.6 $Y=2.11 $X2=0 $Y2=0
cc_673 N_A_618_424#_c_759_n N_CK_c_1164_n 0.00985566f $X=5.455 $Y=2.11 $X2=0
+ $Y2=0
cc_674 N_A_618_424#_c_769_n N_CK_c_1164_n 7.90579e-19 $X=5.455 $Y=2.285 $X2=0
+ $Y2=0
cc_675 N_A_618_424#_M1000_g N_A_1160_89#_M1009_g 0.0565466f $X=5.515 $Y=3.235
+ $X2=0 $Y2=0
cc_676 N_A_618_424#_c_756_n N_A_1160_89#_c_1350_n 0.00145834f $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_677 N_A_618_424#_c_757_n N_A_1160_89#_c_1350_n 6.89974e-19 $X=5.6 $Y=2.11
+ $X2=0 $Y2=0
cc_678 N_A_618_424#_c_759_n N_A_1160_89#_c_1350_n 0.00103465f $X=5.455 $Y=2.11
+ $X2=0 $Y2=0
cc_679 N_A_618_424#_c_756_n N_A_1160_89#_c_1351_n 0.00136902f $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_680 N_A_618_424#_c_757_n N_A_1160_89#_c_1351_n 4.36292e-19 $X=5.6 $Y=2.11
+ $X2=0 $Y2=0
cc_681 N_A_618_424#_c_759_n N_A_1160_89#_c_1351_n 0.0011802f $X=5.455 $Y=2.11
+ $X2=0 $Y2=0
cc_682 N_A_618_424#_c_769_n N_A_1160_89#_c_1351_n 0.0565466f $X=5.455 $Y=2.285
+ $X2=0 $Y2=0
cc_683 N_A_618_424#_c_776_n N_A_1160_89#_c_1385_n 0.0313767f $X=6.52 $Y=2.955
+ $X2=0 $Y2=0
cc_684 N_A_618_424#_c_776_n N_A_1160_89#_c_1389_n 0.00815518f $X=6.52 $Y=2.955
+ $X2=0 $Y2=0
cc_685 N_A_618_424#_c_746_n N_A_1160_89#_c_1355_n 0.0101818f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_686 N_A_618_424#_c_779_n N_A_1160_89#_c_1358_n 0.00734016f $X=6.785 $Y=2.705
+ $X2=0 $Y2=0
cc_687 N_A_618_424#_c_753_n N_A_1160_89#_c_1358_n 0.00206046f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_688 N_A_618_424#_c_761_n N_A_1160_89#_c_1358_n 0.0155125f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_689 N_A_618_424#_c_746_n N_A_1160_89#_c_1359_n 9.27607e-19 $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_690 N_A_618_424#_c_756_n N_A_1160_89#_c_1359_n 0.00382734f $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_691 N_A_618_424#_c_757_n N_A_1160_89#_c_1359_n 0.00126344f $X=5.6 $Y=2.11
+ $X2=0 $Y2=0
cc_692 N_A_618_424#_c_756_n N_A_1160_89#_c_1361_n 8.07535e-19 $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_693 N_A_618_424#_c_746_n N_A_1160_89#_c_1363_n 0.00167736f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_694 N_A_618_424#_c_753_n N_A_1160_89#_c_1363_n 0.00161719f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_695 N_A_618_424#_c_779_n N_A_1160_89#_c_1364_n 0.00931805f $X=6.785 $Y=2.705
+ $X2=0 $Y2=0
cc_696 N_A_618_424#_c_871_p N_A_1160_89#_c_1364_n 0.00729659f $X=6.605 $Y=2.705
+ $X2=0 $Y2=0
cc_697 N_A_618_424#_c_756_n N_A_1160_89#_c_1364_n 0.0518575f $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_698 N_A_618_424#_c_760_n N_A_1160_89#_c_1364_n 0.025445f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_699 N_A_618_424#_c_761_n N_A_1160_89#_c_1364_n 0.0212559f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_700 N_A_618_424#_c_756_n N_A_1160_89#_c_1365_n 0.0253083f $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_701 N_A_618_424#_c_759_n N_A_1160_89#_c_1365_n 0.0025579f $X=5.455 $Y=2.11
+ $X2=0 $Y2=0
cc_702 N_A_618_424#_c_769_n N_A_1160_89#_c_1365_n 0.00405956f $X=5.455 $Y=2.285
+ $X2=0 $Y2=0
cc_703 N_A_618_424#_c_760_n N_A_1160_89#_c_1366_n 0.0246666f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_704 N_A_618_424#_c_761_n N_A_1160_89#_c_1366_n 0.00761196f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_705 N_A_618_424#_c_746_n N_A_1160_89#_c_1367_n 0.00339939f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_706 N_A_618_424#_c_753_n N_A_1160_89#_c_1367_n 0.00544921f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_707 N_A_618_424#_c_756_n N_A_1160_89#_c_1368_n 0.0100909f $X=6.725 $Y=2.11
+ $X2=0 $Y2=0
cc_708 N_A_618_424#_c_757_n N_A_1160_89#_c_1368_n 8.19742e-19 $X=5.6 $Y=2.11
+ $X2=0 $Y2=0
cc_709 N_A_618_424#_c_759_n N_A_1160_89#_c_1368_n 0.0150485f $X=5.455 $Y=2.11
+ $X2=0 $Y2=0
cc_710 N_A_618_424#_c_769_n N_A_1160_89#_c_1368_n 0.00225243f $X=5.455 $Y=2.285
+ $X2=0 $Y2=0
cc_711 N_A_618_424#_c_746_n N_A_998_115#_M1012_g 0.00404242f $X=6.69 $Y=1.76
+ $X2=8.71 $Y2=0.575
cc_712 N_A_618_424#_c_776_n N_A_998_115#_M1006_g 0.00440688f $X=6.52 $Y=2.955
+ $X2=0 $Y2=0
cc_713 N_A_618_424#_c_746_n N_A_998_115#_M1006_g 0.00190027f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_714 N_A_618_424#_c_779_n N_A_998_115#_M1006_g 0.00370122f $X=6.785 $Y=2.705
+ $X2=0 $Y2=0
cc_715 N_A_618_424#_c_753_n N_A_998_115#_M1006_g 0.00175055f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_716 N_A_618_424#_c_760_n N_A_998_115#_M1006_g 7.50221e-19 $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_717 N_A_618_424#_c_761_n N_A_998_115#_M1006_g 0.00735884f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_718 N_A_618_424#_c_744_n N_A_998_115#_c_1599_n 0.00843004f $X=5.37 $Y=2.11
+ $X2=0 $Y2=0
cc_719 N_A_618_424#_c_745_n N_A_998_115#_c_1599_n 0.00323798f $X=5.06 $Y=2.11
+ $X2=0 $Y2=0
cc_720 N_A_618_424#_c_754_n N_A_998_115#_c_1599_n 0.012754f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_721 N_A_618_424#_c_757_n N_A_998_115#_c_1599_n 0.00146098f $X=5.6 $Y=2.11
+ $X2=0 $Y2=0
cc_722 N_A_618_424#_c_759_n N_A_998_115#_c_1599_n 0.00103871f $X=5.455 $Y=2.11
+ $X2=0 $Y2=0
cc_723 N_A_618_424#_c_769_n N_A_998_115#_c_1599_n 0.00150627f $X=5.455 $Y=2.285
+ $X2=0 $Y2=0
cc_724 N_A_618_424#_c_742_n N_A_998_115#_c_1554_n 9.01642e-19 $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_725 N_A_618_424#_c_743_n N_A_998_115#_c_1554_n 0.00191034f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_726 N_A_618_424#_c_766_n N_A_998_115#_c_1554_n 0.00389012f $X=4.975 $Y=1.205
+ $X2=0 $Y2=0
cc_727 N_A_618_424#_c_742_n N_A_998_115#_c_1557_n 0.0123759f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_728 N_A_618_424#_c_743_n N_A_998_115#_c_1557_n 0.0042095f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_729 N_A_618_424#_c_744_n N_A_998_115#_c_1557_n 0.00195757f $X=5.37 $Y=2.11
+ $X2=0 $Y2=0
cc_730 N_A_618_424#_c_742_n N_A_998_115#_c_1558_n 6.325e-19 $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_731 N_A_618_424#_c_743_n N_A_998_115#_c_1558_n 3.88864e-19 $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_732 N_A_618_424#_c_754_n N_A_998_115#_c_1558_n 0.0128239f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_733 N_A_618_424#_c_746_n N_A_998_115#_c_1559_n 0.016053f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_734 N_A_618_424#_c_753_n N_A_998_115#_c_1559_n 0.00391402f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_735 N_A_618_424#_c_760_n N_A_998_115#_c_1559_n 0.0080672f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_736 N_A_618_424#_c_742_n N_A_998_115#_c_1561_n 0.00114522f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_737 N_A_618_424#_c_743_n N_A_998_115#_c_1561_n 4.42421e-19 $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_738 N_A_618_424#_c_744_n N_A_998_115#_c_1561_n 6.62932e-19 $X=5.37 $Y=2.11
+ $X2=0 $Y2=0
cc_739 N_A_618_424#_c_754_n N_A_998_115#_c_1561_n 0.00662656f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_740 N_A_618_424#_c_742_n N_A_998_115#_c_1562_n 0.0571231f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_741 N_A_618_424#_c_743_n N_A_998_115#_c_1562_n 0.00215979f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_742 N_A_618_424#_c_745_n N_A_998_115#_c_1562_n 0.0116326f $X=5.06 $Y=2.11
+ $X2=0 $Y2=0
cc_743 N_A_618_424#_c_754_n N_A_998_115#_c_1562_n 0.020361f $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_744 N_A_618_424#_c_757_n N_A_998_115#_c_1562_n 6.61118e-19 $X=5.6 $Y=2.11
+ $X2=0 $Y2=0
cc_745 N_A_618_424#_c_759_n N_A_998_115#_c_1562_n 0.00613815f $X=5.455 $Y=2.11
+ $X2=0 $Y2=0
cc_746 N_A_618_424#_c_742_n N_A_998_115#_c_1563_n 0.0169532f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_747 N_A_618_424#_c_743_n N_A_998_115#_c_1563_n 0.00154744f $X=4.975 $Y=1.37
+ $X2=0 $Y2=0
cc_748 N_A_618_424#_c_744_n N_A_998_115#_c_1563_n 0.00114215f $X=5.37 $Y=2.11
+ $X2=0 $Y2=0
cc_749 N_A_618_424#_c_754_n N_A_998_115#_c_1563_n 2.84338e-19 $X=5.31 $Y=2.11
+ $X2=0 $Y2=0
cc_750 N_A_618_424#_c_766_n N_A_998_115#_c_1563_n 0.00321467f $X=4.975 $Y=1.205
+ $X2=0 $Y2=0
cc_751 N_A_618_424#_c_746_n N_A_998_115#_c_1564_n 0.00181561f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_752 N_A_618_424#_c_753_n N_A_998_115#_c_1564_n 0.00133282f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_753 N_A_618_424#_c_760_n N_A_998_115#_c_1564_n 0.00527522f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_754 N_A_618_424#_c_746_n N_A_998_115#_c_1565_n 0.0201321f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_755 N_A_618_424#_c_760_n N_A_998_115#_c_1565_n 0.00103848f $X=6.87 $Y=2.11
+ $X2=0 $Y2=0
cc_756 N_A_618_424#_c_746_n N_A_998_115#_c_1567_n 0.00258415f $X=6.69 $Y=1.76
+ $X2=0 $Y2=0
cc_757 N_A_618_424#_c_753_n N_A_998_115#_c_1567_n 0.00141635f $X=6.87 $Y=1.845
+ $X2=0 $Y2=0
cc_758 N_A_217_605#_c_1014_n N_CK_c_1138_n 0.00253253f $X=4.06 $Y=1.37 $X2=4.2
+ $Y2=0.575
cc_759 N_A_217_605#_c_1014_n N_CK_c_1139_n 0.00296105f $X=4.06 $Y=1.37 $X2=5.95
+ $Y2=0.575
cc_760 N_A_217_605#_c_1006_n N_CK_M1017_g 0.114035f $X=4.2 $Y=2.285 $X2=0 $Y2=0
cc_761 N_A_217_605#_c_1013_n N_CK_M1017_g 0.00486364f $X=4.295 $Y=2.285 $X2=0
+ $Y2=0
cc_762 N_A_217_605#_c_1005_n N_CK_c_1142_n 0.0342351f $X=4.2 $Y=1.37 $X2=0 $Y2=0
cc_763 N_A_217_605#_c_1006_n N_CK_c_1142_n 0.0307748f $X=4.2 $Y=2.285 $X2=0
+ $Y2=0
cc_764 N_A_217_605#_c_1013_n N_CK_c_1142_n 0.0113171f $X=4.295 $Y=2.285 $X2=0
+ $Y2=0
cc_765 N_A_217_605#_c_1014_n N_CK_c_1142_n 0.00486036f $X=4.06 $Y=1.37 $X2=0
+ $Y2=0
cc_766 N_A_217_605#_c_1061_n N_CK_c_1142_n 4.12801e-19 $X=4.205 $Y=1.37 $X2=0
+ $Y2=0
cc_767 N_A_217_605#_c_1016_n N_CK_c_1142_n 8.69982e-19 $X=4.205 $Y=1.37 $X2=0
+ $Y2=0
cc_768 N_A_217_605#_c_1009_n N_CK_M1003_g 0.110621f $X=4.48 $Y=2.285 $X2=0 $Y2=0
cc_769 N_A_217_605#_M1022_g N_A_998_115#_c_1639_n 9.13132e-19 $X=4.125 $Y=3.235
+ $X2=0 $Y2=0
cc_770 N_A_217_605#_M1014_g N_A_998_115#_c_1639_n 0.0096885f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_771 N_A_217_605#_c_1007_n N_A_998_115#_c_1558_n 0.00229064f $X=4.48 $Y=1.37
+ $X2=0 $Y2=0
cc_772 N_A_217_605#_c_1061_n N_A_998_115#_c_1558_n 0.0241863f $X=4.205 $Y=1.37
+ $X2=0 $Y2=0
cc_773 N_A_217_605#_c_1016_n N_A_998_115#_c_1558_n 0.0012094f $X=4.205 $Y=1.37
+ $X2=0 $Y2=0
cc_774 N_A_217_605#_M1022_g N_A_998_115#_c_1562_n 9.36754e-19 $X=4.125 $Y=3.235
+ $X2=0 $Y2=0
cc_775 N_A_217_605#_M1025_g N_A_998_115#_c_1562_n 0.00190555f $X=4.555 $Y=0.835
+ $X2=0 $Y2=0
cc_776 N_A_217_605#_M1014_g N_A_998_115#_c_1562_n 0.00479454f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_777 N_A_217_605#_c_1007_n N_A_998_115#_c_1562_n 0.0061959f $X=4.48 $Y=1.37
+ $X2=0 $Y2=0
cc_778 N_A_217_605#_c_1009_n N_A_998_115#_c_1562_n 0.00738718f $X=4.48 $Y=2.285
+ $X2=0 $Y2=0
cc_779 N_A_217_605#_c_1013_n N_A_998_115#_c_1562_n 0.0702347f $X=4.295 $Y=2.285
+ $X2=0 $Y2=0
cc_780 N_A_217_605#_c_1061_n N_A_998_115#_c_1562_n 4.18442e-19 $X=4.205 $Y=1.37
+ $X2=0 $Y2=0
cc_781 N_A_217_605#_c_1016_n N_A_998_115#_c_1562_n 0.0157315f $X=4.205 $Y=1.37
+ $X2=0 $Y2=0
cc_782 N_CK_c_1153_n N_A_1160_89#_M1009_g 0.0422237f $X=6.305 $Y=2.45 $X2=0
+ $Y2=0
cc_783 N_CK_c_1159_n N_A_1160_89#_M1009_g 5.64099e-19 $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_784 N_CK_M1020_g N_A_1160_89#_c_1345_n 0.0575597f $X=5.515 $Y=0.835 $X2=0
+ $Y2=0
cc_785 N_CK_c_1148_n N_A_1160_89#_c_1345_n 0.0170151f $X=6.305 $Y=1.205 $X2=0
+ $Y2=0
cc_786 N_CK_c_1154_n N_A_1160_89#_c_1349_n 0.0101199f $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_787 N_CK_c_1158_n N_A_1160_89#_c_1349_n 0.00850844f $X=6.385 $Y=1.28 $X2=0
+ $Y2=0
cc_788 N_CK_c_1154_n N_A_1160_89#_c_1350_n 0.00666671f $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_789 N_CK_c_1161_n N_A_1160_89#_c_1350_n 4.90616e-19 $X=6.305 $Y=1.74 $X2=0
+ $Y2=0
cc_790 N_CK_c_1153_n N_A_1160_89#_c_1351_n 0.00547635f $X=6.305 $Y=2.45 $X2=0
+ $Y2=0
cc_791 N_CK_c_1159_n N_A_1160_89#_c_1351_n 3.94643e-19 $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_792 N_CK_c_1154_n N_A_1160_89#_c_1359_n 7.5283e-19 $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_793 N_CK_c_1160_n N_A_1160_89#_c_1359_n 0.0121286f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_794 N_CK_c_1246_n N_A_1160_89#_c_1359_n 8.23182e-19 $X=5.6 $Y=1.74 $X2=0
+ $Y2=0
cc_795 N_CK_c_1161_n N_A_1160_89#_c_1359_n 0.0261745f $X=6.305 $Y=1.74 $X2=0
+ $Y2=0
cc_796 CK N_A_1160_89#_c_1359_n 9.31723e-19 $X=6.305 $Y=1.745 $X2=0 $Y2=0
cc_797 N_CK_c_1163_n N_A_1160_89#_c_1359_n 0.00126849f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_798 N_CK_c_1164_n N_A_1160_89#_c_1359_n 0.00808477f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_799 N_CK_c_1154_n N_A_1160_89#_c_1361_n 0.0213894f $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_800 N_CK_c_1160_n N_A_1160_89#_c_1361_n 0.00306708f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_801 N_CK_c_1161_n N_A_1160_89#_c_1361_n 0.0013718f $X=6.305 $Y=1.74 $X2=0
+ $Y2=0
cc_802 CK N_A_1160_89#_c_1361_n 4.68327e-19 $X=6.305 $Y=1.745 $X2=0 $Y2=0
cc_803 N_CK_c_1164_n N_A_1160_89#_c_1361_n 7.17123e-19 $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_804 N_CK_c_1153_n N_A_1160_89#_c_1364_n 0.00315539f $X=6.305 $Y=2.45 $X2=0
+ $Y2=0
cc_805 N_CK_M1029_g N_A_1160_89#_c_1364_n 0.00893989f $X=6.305 $Y=3.235 $X2=0
+ $Y2=0
cc_806 N_CK_c_1159_n N_A_1160_89#_c_1364_n 0.0119083f $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_807 N_CK_M1029_g N_A_1160_89#_c_1365_n 4.63789e-19 $X=6.305 $Y=3.235 $X2=0
+ $Y2=0
cc_808 N_CK_c_1159_n N_A_1160_89#_c_1365_n 9.171e-19 $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_809 N_CK_c_1153_n N_A_1160_89#_c_1368_n 0.00264666f $X=6.305 $Y=2.45 $X2=0
+ $Y2=0
cc_810 N_CK_c_1154_n N_A_1160_89#_c_1368_n 2.0664e-19 $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_811 N_CK_c_1159_n N_A_1160_89#_c_1368_n 0.0214867f $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_812 N_CK_c_1161_n N_A_1160_89#_c_1368_n 0.00567759f $X=6.305 $Y=1.74 $X2=0
+ $Y2=0
cc_813 N_CK_M1020_g N_A_1160_89#_c_1372_n 0.00905991f $X=5.515 $Y=0.835 $X2=0
+ $Y2=0
cc_814 N_CK_c_1163_n N_A_1160_89#_c_1372_n 0.0260042f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_815 N_CK_c_1153_n N_A_998_115#_M1006_g 0.00580112f $X=6.305 $Y=2.45 $X2=0
+ $Y2=0
cc_816 N_CK_c_1154_n N_A_998_115#_M1006_g 0.00656891f $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_817 N_CK_M1003_g N_A_998_115#_c_1599_n 0.0162544f $X=4.915 $Y=3.235 $X2=0
+ $Y2=0
cc_818 N_CK_M1020_g N_A_998_115#_c_1554_n 0.0131134f $X=5.515 $Y=0.835 $X2=0
+ $Y2=0
cc_819 N_CK_c_1142_n N_A_998_115#_c_1557_n 0.00156696f $X=4.84 $Y=1.82 $X2=0
+ $Y2=0
cc_820 N_CK_c_1144_n N_A_998_115#_c_1557_n 0.00141359f $X=5.32 $Y=1.82 $X2=0
+ $Y2=0
cc_821 N_CK_c_1157_n N_A_998_115#_c_1557_n 5.19983e-19 $X=4.915 $Y=1.82 $X2=0
+ $Y2=0
cc_822 N_CK_c_1142_n N_A_998_115#_c_1558_n 0.00120486f $X=4.84 $Y=1.82 $X2=0
+ $Y2=0
cc_823 N_CK_M1020_g N_A_998_115#_c_1559_n 0.00393577f $X=5.515 $Y=0.835 $X2=0
+ $Y2=0
cc_824 N_CK_c_1154_n N_A_998_115#_c_1559_n 0.00357331f $X=6.385 $Y=2.12 $X2=0
+ $Y2=0
cc_825 N_CK_c_1158_n N_A_998_115#_c_1559_n 0.00429194f $X=6.385 $Y=1.28 $X2=0
+ $Y2=0
cc_826 N_CK_c_1160_n N_A_998_115#_c_1559_n 0.0465449f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_827 N_CK_c_1246_n N_A_998_115#_c_1559_n 0.0139023f $X=5.6 $Y=1.74 $X2=0 $Y2=0
cc_828 N_CK_c_1161_n N_A_998_115#_c_1559_n 0.00187144f $X=6.305 $Y=1.74 $X2=0
+ $Y2=0
cc_829 CK N_A_998_115#_c_1559_n 0.0272835f $X=6.305 $Y=1.745 $X2=0 $Y2=0
cc_830 N_CK_c_1163_n N_A_998_115#_c_1559_n 5.08054e-19 $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_831 N_CK_c_1164_n N_A_998_115#_c_1559_n 0.00283556f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_832 N_CK_c_1144_n N_A_998_115#_c_1561_n 6.94944e-19 $X=5.32 $Y=1.82 $X2=0
+ $Y2=0
cc_833 N_CK_M1020_g N_A_998_115#_c_1561_n 0.00225742f $X=5.515 $Y=0.835 $X2=0
+ $Y2=0
cc_834 N_CK_c_1246_n N_A_998_115#_c_1561_n 0.0127467f $X=5.6 $Y=1.74 $X2=0 $Y2=0
cc_835 N_CK_c_1163_n N_A_998_115#_c_1561_n 0.0020361f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_836 N_CK_c_1164_n N_A_998_115#_c_1561_n 0.0012656f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_837 N_CK_c_1142_n N_A_998_115#_c_1562_n 0.0123066f $X=4.84 $Y=1.82 $X2=0
+ $Y2=0
cc_838 N_CK_M1003_g N_A_998_115#_c_1562_n 0.0111407f $X=4.915 $Y=3.235 $X2=0
+ $Y2=0
cc_839 N_CK_c_1163_n N_A_998_115#_c_1563_n 0.00206196f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_840 N_CK_c_1164_n N_A_998_115#_c_1563_n 0.00758189f $X=5.455 $Y=1.725 $X2=0
+ $Y2=0
cc_841 N_CK_c_1158_n N_A_998_115#_c_1567_n 0.00823349f $X=6.385 $Y=1.28 $X2=0
+ $Y2=0
cc_842 N_A_1160_89#_c_1355_n N_A_998_115#_M1012_g 0.00736252f $X=7.47 $Y=0.74
+ $X2=8.71 $Y2=0.575
cc_843 N_A_1160_89#_c_1388_n N_A_998_115#_M1006_g 0.0156817f $X=7.385 $Y=3.045
+ $X2=0 $Y2=0
cc_844 N_A_1160_89#_c_1358_n N_A_998_115#_M1006_g 0.0127145f $X=7.47 $Y=2.96
+ $X2=0 $Y2=0
cc_845 N_A_1160_89#_c_1363_n N_A_998_115#_M1006_g 0.00178263f $X=7.47 $Y=1.74
+ $X2=0 $Y2=0
cc_846 N_A_1160_89#_c_1364_n N_A_998_115#_M1006_g 0.00558185f $X=7.155 $Y=2.48
+ $X2=0 $Y2=0
cc_847 N_A_1160_89#_c_1366_n N_A_998_115#_M1006_g 0.00591057f $X=7.245 $Y=2.395
+ $X2=0 $Y2=0
cc_848 N_A_1160_89#_c_1367_n N_A_998_115#_M1006_g 0.0089178f $X=7.335 $Y=1.737
+ $X2=0 $Y2=0
cc_849 N_A_1160_89#_c_1349_n N_A_998_115#_c_1559_n 0.00346468f $X=5.89 $Y=1.365
+ $X2=0 $Y2=0
cc_850 N_A_1160_89#_c_1359_n N_A_998_115#_c_1559_n 0.00439053f $X=5.935 $Y=2.025
+ $X2=0 $Y2=0
cc_851 N_A_1160_89#_c_1361_n N_A_998_115#_c_1559_n 7.74479e-19 $X=5.965 $Y=1.77
+ $X2=0 $Y2=0
cc_852 N_A_1160_89#_c_1372_n N_A_998_115#_c_1559_n 0.00274919f $X=5.965 $Y=1.605
+ $X2=0 $Y2=0
cc_853 N_A_1160_89#_c_1355_n N_A_998_115#_c_1564_n 0.00286995f $X=7.47 $Y=0.74
+ $X2=0 $Y2=0
cc_854 N_A_1160_89#_c_1367_n N_A_998_115#_c_1564_n 0.00402018f $X=7.335 $Y=1.737
+ $X2=0 $Y2=0
cc_855 N_A_1160_89#_c_1355_n N_A_998_115#_c_1565_n 0.0147498f $X=7.47 $Y=0.74
+ $X2=0 $Y2=0
cc_856 N_A_1160_89#_c_1367_n N_A_998_115#_c_1567_n 4.10276e-19 $X=7.335 $Y=1.737
+ $X2=0 $Y2=0
cc_857 N_A_1160_89#_M1016_g N_QN_M1008_g 0.0210474f $X=8.635 $Y=0.755 $X2=8.71
+ $Y2=0.575
cc_858 N_A_1160_89#_c_1370_n N_QN_M1008_g 3.6337e-19 $X=8.52 $Y=1.74 $X2=8.71
+ $Y2=0.575
cc_859 N_A_1160_89#_c_1374_n N_QN_M1008_g 0.0152125f $X=8.522 $Y=1.575 $X2=8.71
+ $Y2=0.575
cc_860 N_A_1160_89#_c_1353_n N_QN_M1001_g 0.0102953f $X=8.61 $Y=2.375 $X2=0
+ $Y2=0
cc_861 N_A_1160_89#_c_1354_n N_QN_M1001_g 0.0339596f $X=8.61 $Y=2.525 $X2=0
+ $Y2=0
cc_862 N_A_1160_89#_M1016_g N_QN_c_1700_n 0.00760341f $X=8.635 $Y=0.755 $X2=0
+ $Y2=0
cc_863 N_A_1160_89#_c_1352_n N_QN_c_1700_n 0.00327645f $X=8.61 $Y=1.32 $X2=0
+ $Y2=0
cc_864 N_A_1160_89#_c_1352_n N_QN_c_1704_n 0.0108281f $X=8.61 $Y=1.32 $X2=0
+ $Y2=0
cc_865 N_A_1160_89#_c_1369_n N_QN_c_1704_n 0.0037949f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_866 N_A_1160_89#_c_1370_n N_QN_c_1704_n 0.0093039f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_867 N_A_1160_89#_c_1374_n N_QN_c_1704_n 0.00784613f $X=8.522 $Y=1.575 $X2=0
+ $Y2=0
cc_868 N_A_1160_89#_c_1369_n N_QN_c_1706_n 0.00331526f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_869 N_A_1160_89#_c_1370_n N_QN_c_1706_n 0.0101631f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_870 N_A_1160_89#_c_1371_n N_QN_c_1706_n 0.00105631f $X=8.375 $Y=1.74 $X2=0
+ $Y2=0
cc_871 N_A_1160_89#_c_1373_n N_QN_c_1706_n 0.00303508f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_872 N_A_1160_89#_c_1353_n N_QN_c_1707_n 0.0159847f $X=8.61 $Y=2.375 $X2=0
+ $Y2=0
cc_873 N_A_1160_89#_c_1354_n N_QN_c_1707_n 0.00248624f $X=8.61 $Y=2.525 $X2=0
+ $Y2=0
cc_874 N_A_1160_89#_c_1369_n N_QN_c_1707_n 0.00258299f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_875 N_A_1160_89#_c_1370_n N_QN_c_1707_n 0.0046698f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_876 N_A_1160_89#_c_1369_n N_QN_c_1708_n 0.00139444f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_877 N_A_1160_89#_c_1370_n N_QN_c_1708_n 0.00515207f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_878 N_A_1160_89#_c_1371_n N_QN_c_1708_n 4.39196e-19 $X=8.375 $Y=1.74 $X2=0
+ $Y2=0
cc_879 N_A_1160_89#_c_1373_n N_QN_c_1708_n 0.00271474f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_880 N_A_1160_89#_c_1353_n N_QN_c_1709_n 0.00226435f $X=8.61 $Y=2.375 $X2=0
+ $Y2=0
cc_881 N_A_1160_89#_c_1369_n N_QN_c_1709_n 0.00377829f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_882 N_A_1160_89#_c_1370_n N_QN_c_1709_n 0.00978463f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_883 N_A_1160_89#_c_1373_n N_QN_c_1709_n 0.0019182f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_884 N_A_1160_89#_c_1374_n N_QN_c_1709_n 0.00380475f $X=8.522 $Y=1.575 $X2=0
+ $Y2=0
cc_885 N_A_1160_89#_c_1369_n N_QN_c_1710_n 4.60229e-19 $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_886 N_A_1160_89#_c_1370_n N_QN_c_1710_n 5.0648e-19 $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_887 N_A_1160_89#_c_1373_n N_QN_c_1710_n 0.0211392f $X=8.52 $Y=1.74 $X2=0
+ $Y2=0
cc_888 N_A_1160_89#_M1011_g N_QN_c_1711_n 0.0164234f $X=8.635 $Y=3.445 $X2=0
+ $Y2=0
cc_889 N_A_1160_89#_c_1353_n N_QN_c_1711_n 0.00567875f $X=8.61 $Y=2.375 $X2=0
+ $Y2=0
cc_890 N_A_1160_89#_M1011_g QN 0.00233857f $X=8.635 $Y=3.445 $X2=0 $Y2=0
cc_891 N_A_1160_89#_c_1354_n QN 0.00508004f $X=8.61 $Y=2.525 $X2=0 $Y2=0
cc_892 N_A_1160_89#_c_1358_n QN 0.00513409f $X=7.47 $Y=2.96 $X2=0 $Y2=0
cc_893 N_A_1160_89#_c_1369_n QN 0.00881422f $X=8.52 $Y=1.74 $X2=0 $Y2=0
cc_894 N_A_1160_89#_c_1370_n QN 0.00286804f $X=8.52 $Y=1.74 $X2=0 $Y2=0
cc_895 N_A_1160_89#_c_1371_n QN 0.00487781f $X=8.375 $Y=1.74 $X2=0 $Y2=0
cc_896 N_A_1160_89#_c_1388_n A_1466_605# 0.00433061f $X=7.385 $Y=3.045 $X2=0.135
+ $Y2=0.575
cc_897 N_A_998_115#_c_1599_n A_926_521# 0.00342591f $X=5.045 $Y=2.705 $X2=0.135
+ $Y2=0.575
cc_898 N_A_998_115#_c_1639_n A_926_521# 0.00144354f $X=4.72 $Y=2.705 $X2=0.135
+ $Y2=0.575
cc_899 N_QN_M1008_g N_Q_c_1791_n 5.62519e-19 $X=9.065 $Y=0.755 $X2=8.71
+ $Y2=0.575
cc_900 N_QN_M1001_g N_Q_c_1795_n 0.00409136f $X=9.065 $Y=3.445 $X2=0 $Y2=0
cc_901 N_QN_M1008_g N_Q_c_1793_n 0.0383548f $X=9.065 $Y=0.755 $X2=0 $Y2=0
cc_902 N_QN_c_1704_n N_Q_c_1793_n 0.0111776f $X=8.92 $Y=1.37 $X2=0 $Y2=0
cc_903 N_QN_c_1707_n N_Q_c_1793_n 0.0111776f $X=8.92 $Y=2.285 $X2=0 $Y2=0
cc_904 N_QN_c_1709_n N_Q_c_1793_n 0.0438362f $X=9.005 $Y=1.915 $X2=0 $Y2=0
cc_905 N_QN_M1008_g N_Q_c_1794_n 0.00695117f $X=9.065 $Y=0.755 $X2=0 $Y2=0
cc_906 N_QN_M1001_g Q 0.0131514f $X=9.065 $Y=3.445 $X2=0 $Y2=0
cc_907 N_QN_c_1707_n Q 0.00245821f $X=8.92 $Y=2.285 $X2=0 $Y2=0
cc_908 N_QN_M1001_g N_Q_c_1802_n 0.00614447f $X=9.065 $Y=3.445 $X2=0 $Y2=0
