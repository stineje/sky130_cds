magic
tech sky130A
magscale 1 2
timestamp 1606864592
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 288 1341
<< nmos >>
rect 80 115 110 263
rect 166 115 196 263
<< pmoshvt >>
rect 80 817 110 1217
rect 166 817 196 1217
<< ndiff >>
rect 27 199 80 263
rect 27 131 35 199
rect 69 131 80 199
rect 27 115 80 131
rect 110 199 166 263
rect 110 131 121 199
rect 155 131 166 199
rect 110 115 166 131
rect 196 199 249 263
rect 196 131 207 199
rect 241 131 249 199
rect 196 115 249 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 861 35 1201
rect 69 861 80 1201
rect 27 817 80 861
rect 110 1201 166 1217
rect 110 861 121 1201
rect 155 861 166 1201
rect 110 817 166 861
rect 196 1201 249 1217
rect 196 861 207 1201
rect 241 861 249 1201
rect 196 817 249 861
<< ndiffc >>
rect 35 131 69 199
rect 121 131 155 199
rect 207 131 241 199
<< pdiffc >>
rect 35 861 69 1201
rect 121 861 155 1201
rect 207 861 241 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 80 529 110 817
rect 166 602 196 817
rect 166 572 251 602
rect 80 513 154 529
rect 80 479 110 513
rect 144 479 154 513
rect 80 463 154 479
rect 80 263 110 463
rect 221 420 251 572
rect 166 404 251 420
rect 166 370 176 404
rect 210 370 251 404
rect 166 354 251 370
rect 166 263 196 354
rect 80 89 110 115
rect 166 89 196 115
<< polycont >>
rect 110 479 144 513
rect 176 370 210 404
<< locali >>
rect 0 1311 286 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 286 1311
rect 35 1201 69 1217
rect 35 404 69 861
rect 121 1201 155 1271
rect 121 845 155 861
rect 207 1201 241 1217
rect 110 513 144 649
rect 207 609 241 861
rect 110 463 144 479
rect 176 404 210 420
rect 35 370 176 404
rect 35 199 69 370
rect 176 354 210 370
rect 35 115 69 131
rect 121 199 155 215
rect 121 61 155 131
rect 207 199 241 279
rect 207 115 241 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 110 649 144 683
rect 207 575 241 609
rect 207 279 241 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 286 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 286 1311
rect 0 1271 286 1277
rect 98 683 156 689
rect 64 649 110 683
rect 144 649 156 683
rect 98 643 156 649
rect 195 609 253 615
rect 195 575 207 609
rect 241 575 253 609
rect 195 569 253 575
rect 207 319 241 569
rect 195 313 253 319
rect 195 279 207 313
rect 241 279 253 313
rect 195 273 253 279
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 127 666 127 666 1 A
port 1 n
rlabel metal1 214 452 214 452 1 Y
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
