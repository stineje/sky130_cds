magic
tech sky130A
magscale 1 2
timestamp 1606864618
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 375 1341
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
<< nmoslvt >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 166 315
rect 110 131 121 267
rect 155 131 166 267
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 267 335 315
rect 282 131 293 267
rect 327 131 335 267
rect 282 115 335 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 166 1217
rect 110 657 121 1201
rect 155 657 166 1201
rect 110 617 166 657
rect 196 1201 252 1217
rect 196 657 207 1201
rect 241 657 252 1201
rect 196 617 252 657
rect 282 1201 335 1217
rect 282 657 293 1201
rect 327 657 335 1201
rect 282 617 335 657
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 207 131 241 267
rect 293 131 327 267
<< pdiffc >>
rect 35 793 69 1201
rect 121 657 155 1201
rect 207 657 241 1201
rect 293 657 327 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 80 592 110 617
rect 166 592 196 617
rect 252 592 282 617
rect 80 562 282 592
rect 80 494 110 562
rect 80 478 134 494
rect 80 444 90 478
rect 124 444 134 478
rect 80 428 134 444
rect 80 370 110 428
rect 80 340 282 370
rect 80 315 110 340
rect 166 315 196 340
rect 252 315 282 340
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
<< polycont >>
rect 90 444 124 478
<< locali >>
rect 0 1311 374 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 374 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 47 478 81 649
rect 121 609 155 657
rect 207 1201 241 1271
rect 207 641 241 657
rect 293 1201 327 1217
rect 293 609 327 657
rect 47 444 90 478
rect 124 444 140 478
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 279
rect 121 115 155 131
rect 207 267 241 283
rect 207 61 241 131
rect 293 267 327 279
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 47 649 81 683
rect 121 575 155 609
rect 293 575 327 609
rect 121 279 155 313
rect 293 279 327 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 374 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 374 1311
rect 0 1271 374 1277
rect 35 683 93 689
rect 35 649 47 683
rect 81 649 127 683
rect 35 643 93 649
rect 109 609 167 615
rect 281 609 339 615
rect 109 575 121 609
rect 155 575 293 609
rect 327 575 339 609
rect 109 569 167 575
rect 281 569 339 575
rect 121 319 155 569
rect 293 319 327 569
rect 109 313 167 319
rect 281 313 339 319
rect 109 279 121 313
rect 155 279 293 313
rect 327 279 339 313
rect 109 273 167 279
rect 281 273 339 279
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 152 440 152 440 1 Y
port 1 n
rlabel metal1 64 665 64 665 1 A
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
