* File: sky130_osu_sc_18T_hs__oai22_l.pex.spice
* Created: Fri Nov 12 13:52:13 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%GND 1 23 25 33 48 50
r43 48 50 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r44 35 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r45 31 44 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r46 31 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r47 25 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r48 23 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r49 23 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r50 23 35 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r51 23 25 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r52 1 33 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%VDD 1 2 21 25 29 38 49 53
r26 49 53 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r27 45 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r28 38 41 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.91 $Y=4.135
+ $X2=1.91 $Y2=5.835
r29 36 47 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.91 $Y=6.355
+ $X2=1.91 $Y2=6.507
r30 36 41 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.91 $Y=6.355
+ $X2=1.91 $Y2=5.835
r31 34 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.47 $X2=1.7
+ $Y2=6.47
r32 32 34 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r33 30 45 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r34 30 32 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r35 29 47 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=6.507
+ $X2=1.91 $Y2=6.507
r36 29 34 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=6.507
+ $X2=1.7 $Y2=6.507
r37 25 28 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r38 23 45 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r39 23 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r40 21 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r41 21 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r42 21 45 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r43 2 41 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.77
+ $Y=3.085 $X2=1.91 $Y2=5.835
r44 2 38 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=1.77
+ $Y=3.085 $X2=1.91 $Y2=4.135
r45 1 28 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r46 1 25 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%A0 3 5 8 12 15 16 19 25
r36 22 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.415 $Y=3.33
+ $X2=0.415 $Y2=3.33
r37 19 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.415 $Y=2.76
+ $X2=0.415 $Y2=3.33
r38 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=2.76 $X2=0.415 $Y2=2.76
r39 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.76
+ $X2=0.415 $Y2=2.925
r40 15 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=2.76
+ $X2=0.415 $Y2=2.595
r41 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=0.355 $Y=1.775
+ $X2=0.475 $Y2=1.775
r42 8 17 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.925
r43 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.775
r44 3 5 200.833 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.7
+ $X2=0.475 $Y2=1.075
r45 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.355 $Y=1.85
+ $X2=0.355 $Y2=1.775
r46 1 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.355 $Y=1.85
+ $X2=0.355 $Y2=2.595
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%A1 3 7 10 15 18 22
c50 22 0 1.46676e-19 $X=0.895 $Y=2.96
r51 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.895 $Y=2.96
+ $X2=0.895 $Y2=2.96
r52 18 19 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=2.96
+ $X2=0.855 $Y2=2.875
r53 15 19 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.815 $Y=2.22
+ $X2=0.815 $Y2=2.875
r54 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.815
+ $Y=2.22 $X2=0.815 $Y2=2.22
r55 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.815 $Y=2.22
+ $X2=0.815 $Y2=2.355
r56 10 11 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.815 $Y=2.22
+ $X2=0.815 $Y2=2.085
r57 7 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.085
r58 3 12 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=0.835 $Y=4.585
+ $X2=0.835 $Y2=2.355
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%B0 3 7 10 15 20 23
c51 15 0 1.46676e-19 $X=1.2 $Y=2.59
r52 17 20 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.88
+ $X2=1.325 $Y2=1.88
r53 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.59 $X2=1.2
+ $Y2=2.59
r54 13 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=2.045 $X2=1.2
+ $Y2=1.88
r55 13 15 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.2 $Y=2.045
+ $X2=1.2 $Y2=2.59
r56 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.88 $X2=1.325 $Y2=1.88
r57 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.88
+ $X2=1.325 $Y2=2.045
r58 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.88
+ $X2=1.325 $Y2=1.715
r59 7 12 1302.43 $w=1.5e-07 $l=2.54e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.045
r60 3 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=1.715
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%B1 3 6 10 11 15 18 23
r30 18 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.005 $Y=2.225
+ $X2=2.005 $Y2=2.225
r31 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=2.225 $X2=2.005 $Y2=2.225
r32 12 15 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.765 $Y=2.225
+ $X2=2.005 $Y2=2.225
r33 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.73 $Y=2.81
+ $X2=1.73 $Y2=2.96
r34 8 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.39
+ $X2=1.765 $Y2=2.225
r35 8 10 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.765 $Y=2.39
+ $X2=1.765 $Y2=2.81
r36 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.06
+ $X2=1.765 $Y2=2.225
r37 4 6 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=1.765 $Y=2.06
+ $X2=1.765 $Y2=1.075
r38 3 11 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.695 $Y=4.585
+ $X2=1.695 $Y2=2.96
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%Y 1 3 11 15 16 17 19 23 28 30 33
r48 28 33 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.665 $Y=1.735
+ $X2=1.665 $Y2=1.85
r49 27 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.665 $Y=1.595
+ $X2=1.665 $Y2=1.48
r50 27 28 0.134804 $w=1.7e-07 $l=1.4e-07 $layer=MET1_cond $X=1.665 $Y=1.595
+ $X2=1.665 $Y2=1.735
r51 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.665 $Y=1.48
+ $X2=1.665 $Y2=1.48
r52 23 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.665 $Y=1.85
+ $X2=1.665 $Y2=1.85
r53 21 23 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=1.665 $Y2=1.85
r54 17 26 13.286 $w=2.31e-07 $l=2.61954e-07 $layer=LI1_cond $X=1.55 $Y=1.245
+ $X2=1.607 $Y2=1.48
r55 17 19 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.55 $Y=1.245 $X2=1.55
+ $Y2=1.165
r56 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=3.415
+ $X2=1.665 $Y2=3.33
r57 15 16 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.58 $Y=3.415
+ $X2=1.17 $Y2=3.415
r58 11 13 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.085 $Y=3.795
+ $X2=1.085 $Y2=5.835
r59 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.085 $Y=3.5
+ $X2=1.17 $Y2=3.415
r60 9 11 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.085 $Y=3.5
+ $X2=1.085 $Y2=3.795
r61 3 13 171.429 $w=1.7e-07 $l=2.83615e-06 $layer=licon1_PDIFF $count=3 $X=0.91
+ $Y=3.085 $X2=1.085 $Y2=5.835
r62 3 11 171.429 $w=1.7e-07 $l=7.92685e-07 $layer=licon1_PDIFF $count=3 $X=0.91
+ $Y=3.085 $X2=1.085 $Y2=3.795
r63 1 19 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=1.165
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__OAI22_L%A_27_115# 1 2 3 15 17 18 23 24
r22 25 27 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.98 $Y=0.745 $X2=1.98
+ $Y2=0.825
r23 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.895 $Y=0.66
+ $X2=1.98 $Y2=0.745
r24 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=0.66
+ $X2=1.205 $Y2=0.66
r25 20 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.12 $Y=1.335
+ $X2=1.12 $Y2=0.825
r26 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.745
+ $X2=1.205 $Y2=0.66
r27 19 22 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=0.745 $X2=1.12
+ $Y2=0.825
r28 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.42
+ $X2=1.12 $Y2=1.335
r29 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.42
+ $X2=0.345 $Y2=1.42
r30 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.335
+ $X2=0.345 $Y2=1.42
r31 13 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.26 $Y=1.335
+ $X2=0.26 $Y2=0.825
r32 3 27 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r33 2 22 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r34 1 15 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

