* File: sky130_osu_sc_18T_ls__and2_2.pex.spice
* Created: Fri Nov 12 13:39:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__AND2_2%GND 1 2 27 29 37 39 47 55 57
r44 55 57 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r45 45 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.825
r46 39 45 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.305
r47 35 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r48 27 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.19 $X2=1.7
+ $Y2=0.19
r49 27 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r50 27 35 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r51 27 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r52 27 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r53 27 39 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r54 27 40 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r55 27 29 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r56 2 47 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r57 1 37 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_2%VDD 1 2 3 25 29 33 39 43 50 59 63
r36 59 63 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r37 55 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r38 50 53 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r39 48 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.98 $Y=6.355
+ $X2=1.98 $Y2=5.835
r40 46 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.47 $X2=1.7
+ $Y2=6.47
r41 44 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r42 44 46 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.7 $Y2=6.507
r43 43 48 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.98 $Y2=6.355
r44 43 46 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=6.507
+ $X2=1.7 $Y2=6.507
r45 39 42 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r46 37 57 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r47 37 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r48 34 55 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r49 34 36 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.02 $Y2=6.507
r50 33 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r51 33 36 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.02 $Y2=6.507
r52 29 32 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r53 27 55 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r54 27 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r55 25 46 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r56 25 36 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r57 25 55 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r58 3 53 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r59 3 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r60 2 42 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r61 2 39 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r62 1 32 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r63 1 29 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_2%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=3.33
+ $X2=0.275 $Y2=3.33
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.33
+ $X2=0.27 $Y2=3.33
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.765
+ $X2=0.27 $Y2=3.33
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.765 $X2=0.27 $Y2=2.765
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.765
+ $X2=0.475 $Y2=2.765
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=2.765
r38 5 7 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=0.475 $Y=2.93
+ $X2=0.475 $Y2=4.585
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=2.765
r40 1 3 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=0.475 $Y=2.6
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_2%B 3 7 10 14 22
c41 7 0 1.37149e-19 $X=0.905 $Y=4.585
r42 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.96
+ $X2=0.955 $Y2=2.96
r43 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.96
+ $X2=0.95 $Y2=2.96
r44 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.425
+ $X2=0.95 $Y2=2.96
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.425 $X2=0.95 $Y2=2.425
r46 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.59
r47 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.425
+ $X2=0.922 $Y2=2.26
r48 7 12 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.59
r49 3 11 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.835 $Y=1.075
+ $X2=0.835 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_2%A_27_115# 1 3 11 13 15 17 18 22 24 26 27
+ 31 35 37 38 43 49 51 52 53
r87 52 53 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.545
+ $X2=0.65 $Y2=3.715
r88 47 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=0.61 $Y2=1.935
r89 47 49 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.935
+ $X2=1.43 $Y2=1.935
r90 43 45 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.69 $Y=3.795
+ $X2=0.69 $Y2=5.835
r91 43 53 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.795 $X2=0.69
+ $Y2=3.715
r92 39 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=2.02 $X2=0.61
+ $Y2=1.935
r93 39 52 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=2.02
+ $X2=0.61 $Y2=3.545
r94 37 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.61 $Y2=1.935
r95 37 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.935
+ $X2=0.345 $Y2=1.935
r96 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.345 $Y2=1.935
r97 33 35 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r98 31 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.935 $X2=1.43 $Y2=1.935
r99 29 31 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.935 $X2=1.43
+ $Y2=1.935
r100 28 29 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.935
+ $X2=1.37 $Y2=1.935
r101 24 26 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.765 $Y=2.96
+ $X2=1.765 $Y2=4.585
r102 20 31 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.43 $Y2=1.935
r103 20 22 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r104 19 27 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.885
+ $X2=1.352 $Y2=2.885
r105 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.765 $Y2=2.96
r106 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.885
+ $X2=1.445 $Y2=2.885
r107 17 27 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.81
+ $X2=1.352 $Y2=2.885
r108 16 29 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=1.935
r109 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=2.1
+ $X2=1.37 $Y2=2.81
r110 13 27 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.352 $Y2=2.885
r111 13 15 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.335 $Y=2.96
+ $X2=1.335 $Y2=4.585
r112 9 28 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.935
r113 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r114 3 45 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r115 3 43 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.795
r116 1 35 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AND2_2%Y 1 3 10 16 26 29 32
c42 16 0 1.37149e-19 $X=1.55 $Y=2.59
r43 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.59
r44 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.475
+ $X2=1.55 $Y2=2.22
r45 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=1.48
r46 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.595
+ $X2=1.55 $Y2=2.22
r47 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r48 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=2.59
r49 16 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.55 $Y=2.59
+ $X2=1.55 $Y2=3.455
r50 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r51 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r52 3 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r53 3 19 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r54 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

