* File: sky130_osu_sc_15T_ms__dffs_1.spice
* Created: Fri Nov 12 14:42:48 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__dffs_1.pex.spice"
.subckt sky130_osu_sc_15T_ms__dffs_1  GND VDD SN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* VDD	VDD
* GND	GND
MM1016 A_110_115# N_SN_M1016_g N_A_27_115#_M1016_s N_GND_M1016_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.5 A=0.078 P=1.34 MULT=1
MM1002 N_GND_M1002_d N_A_152_89#_M1002_g A_110_115# N_GND_M1016_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.0546 PD=1.57 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1003 A_386_115# N_D_M1003_g N_GND_M1003_s N_GND_M1016_b NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1024 N_A_152_89#_M1024_d N_A_428_89#_M1024_g A_386_115# N_GND_M1016_b NSHORT
+ L=0.15 W=0.74 AD=0.1665 AS=0.0777 PD=1.19 PS=0.95 NRD=13.776 NRS=8.1 M=1
+ R=4.93333 SA=75000.6 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1021 A_578_115# N_CK_M1021_g N_A_152_89#_M1024_d N_GND_M1016_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1665 PD=0.95 PS=1.19 NRD=8.1 NRS=13.776 M=1 R=4.93333
+ SA=75001.1 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1023 N_GND_M1023_d N_A_27_115#_M1023_g A_578_115# N_GND_M1016_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.0777 PD=1.02 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.5 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1017 A_736_115# N_A_27_115#_M1017_g N_GND_M1023_d N_GND_M1016_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1036 PD=0.95 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1011 N_A_808_115#_M1011_d N_CK_M1011_g A_736_115# N_GND_M1016_b NSHORT L=0.15
+ W=0.74 AD=0.1665 AS=0.0777 PD=1.19 PS=0.95 NRD=13.776 NRS=8.1 M=1 R=4.93333
+ SA=75002.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1005 A_928_115# N_A_428_89#_M1005_g N_A_808_115#_M1011_d N_GND_M1016_b NSHORT
+ L=0.15 W=0.74 AD=0.0777 AS=0.1665 PD=0.95 PS=1.19 NRD=8.1 NRS=13.776 M=1
+ R=4.93333 SA=75002.9 SB=75001 A=0.111 P=1.78 MULT=1
MM1008 N_GND_M1008_d N_A_970_89#_M1008_g A_928_115# N_GND_M1016_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.0777 PD=1.02 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75003.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_428_89#_M1006_d N_CK_M1006_g N_GND_M1008_d N_GND_M1016_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 A_1276_115# N_A_808_115#_M1007_g N_A_970_89#_M1007_s N_GND_M1016_b NSHORT
+ L=0.15 W=0.52 AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.5 A=0.078 P=1.34 MULT=1
MM1026 N_GND_M1026_d N_SN_M1026_g A_1276_115# N_GND_M1016_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0546 PD=1.57 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75000.5
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_GND_M1010_d N_A_970_89#_M1010_g N_QN_M1010_s N_GND_M1016_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1028 N_Q_M1028_d N_QN_M1028_g N_GND_M1010_d N_GND_M1016_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_115#_M1012_d N_SN_M1012_g N_VDD_M1012_s N_VDD_M1012_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_VDD_M1027_d N_A_152_89#_M1027_g N_A_27_115#_M1012_d N_VDD_M1012_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1013 A_386_565# N_D_M1013_g N_VDD_M1013_s N_VDD_M1012_b PSHORT L=0.15 W=2
+ AD=0.21 AS=0.53 PD=2.21 PS=4.53 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75003.7 A=0.3 P=4.3 MULT=1
MM1000 N_A_152_89#_M1000_d N_CK_M1000_g A_386_565# N_VDD_M1012_b PSHORT L=0.15
+ W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75000.5 SB=75003.3 A=0.3 P=4.3 MULT=1
MM1025 A_578_565# N_A_428_89#_M1025_g N_A_152_89#_M1000_d N_VDD_M1012_b PSHORT
+ L=0.15 W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75001.1 SB=75002.7 A=0.3 P=4.3 MULT=1
MM1029 N_VDD_M1029_d N_A_27_115#_M1029_g A_578_565# N_VDD_M1012_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001.5
+ SB=75002.4 A=0.3 P=4.3 MULT=1
MM1022 A_736_565# N_A_27_115#_M1022_g N_VDD_M1029_d N_VDD_M1012_b PSHORT L=0.15
+ W=2 AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75001.9
+ SB=75001.9 A=0.3 P=4.3 MULT=1
MM1020 N_A_808_115#_M1020_d N_A_428_89#_M1020_g A_736_565# N_VDD_M1012_b PSHORT
+ L=0.15 W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75002.3 SB=75001.6 A=0.3 P=4.3 MULT=1
MM1014 A_928_565# N_CK_M1014_g N_A_808_115#_M1020_d N_VDD_M1012_b PSHORT L=0.15
+ W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75002.9 SB=75001 A=0.3 P=4.3 MULT=1
MM1018 N_VDD_M1018_d N_A_970_89#_M1018_g A_928_565# N_VDD_M1012_b PSHORT L=0.15
+ W=2 AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75003.3
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1015 N_A_428_89#_M1015_d N_CK_M1015_g N_VDD_M1018_d N_VDD_M1012_b PSHORT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75003.7 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1001 N_A_970_89#_M1001_d N_A_808_115#_M1001_g N_VDD_M1001_s N_VDD_M1012_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_SN_M1004_g N_A_970_89#_M1001_d N_VDD_M1012_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1019 N_VDD_M1019_d N_A_970_89#_M1019_g N_QN_M1019_s N_VDD_M1012_b PSHORT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1009 N_Q_M1009_d N_QN_M1009_g N_VDD_M1019_d N_VDD_M1012_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX30_noxref N_GND_M1016_b N_VDD_M1012_b NWDIODE A=25.8272 P=23.41
pX31_noxref noxref_23 SN SN PROBETYPE=1
pX32_noxref noxref_24 D D PROBETYPE=1
pX33_noxref noxref_25 CK CK PROBETYPE=1
pX34_noxref noxref_26 QN QN PROBETYPE=1
pX35_noxref noxref_27 Q Q PROBETYPE=1
c_1473 A_736_565# 0 1.57671e-19 $X=3.68 $Y=2.825
*
.include "sky130_osu_sc_15T_ms__dffs_1.pxi.spice"
*
.ends
*
*
