magic
tech sky130A
magscale 1 2
timestamp 1612371333
<< nwell >>
rect -9 529 837 1119
<< nmoslvt >>
rect 80 115 110 243
rect 178 115 208 243
rect 250 115 280 243
rect 442 115 472 283
rect 540 115 570 283
rect 626 115 656 283
rect 712 115 742 283
<< pmos >>
rect 80 565 110 965
rect 178 565 208 965
rect 264 565 294 965
rect 362 565 392 965
rect 552 565 582 965
rect 638 565 668 965
rect 710 565 740 965
<< ndiff >>
rect 27 224 80 243
rect 27 131 35 224
rect 69 131 80 224
rect 27 115 80 131
rect 110 224 178 243
rect 110 131 133 224
rect 167 131 178 224
rect 110 115 178 131
rect 208 115 250 243
rect 280 224 333 243
rect 280 131 291 224
rect 325 131 333 224
rect 280 115 333 131
rect 389 233 442 283
rect 389 131 397 233
rect 431 131 442 233
rect 389 115 442 131
rect 472 233 540 283
rect 472 131 495 233
rect 529 131 540 233
rect 472 115 540 131
rect 570 233 626 283
rect 570 131 581 233
rect 615 131 626 233
rect 570 115 626 131
rect 656 247 712 283
rect 656 179 667 247
rect 701 179 712 247
rect 656 115 712 179
rect 742 233 795 283
rect 742 131 753 233
rect 787 131 795 233
rect 742 115 795 131
<< pdiff >>
rect 27 949 80 965
rect 27 609 35 949
rect 69 609 80 949
rect 27 565 80 609
rect 110 949 178 965
rect 110 609 133 949
rect 167 609 178 949
rect 110 565 178 609
rect 208 949 264 965
rect 208 677 219 949
rect 253 677 264 949
rect 208 565 264 677
rect 294 949 362 965
rect 294 677 305 949
rect 339 677 362 949
rect 294 565 362 677
rect 392 949 445 965
rect 392 609 403 949
rect 437 609 445 949
rect 392 565 445 609
rect 499 949 552 965
rect 499 609 507 949
rect 541 609 552 949
rect 499 565 552 609
rect 582 949 638 965
rect 582 609 593 949
rect 627 609 638 949
rect 582 565 638 609
rect 668 565 710 965
rect 740 949 796 965
rect 740 609 751 949
rect 785 609 796 949
rect 740 565 796 609
<< ndiffc >>
rect 35 131 69 224
rect 133 131 167 224
rect 291 131 325 224
rect 397 131 431 233
rect 495 131 529 233
rect 581 131 615 233
rect 667 179 701 247
rect 753 131 787 233
<< pdiffc >>
rect 35 609 69 949
rect 133 609 167 949
rect 219 677 253 949
rect 305 677 339 949
rect 403 609 437 949
rect 507 609 541 949
rect 593 609 627 949
rect 751 609 785 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
rect 571 1049 595 1083
rect 629 1049 653 1083
rect 707 1049 731 1083
rect 765 1049 789 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
rect 595 1049 629 1083
rect 731 1049 765 1083
<< poly >>
rect 80 965 110 991
rect 178 965 208 991
rect 264 965 294 991
rect 362 965 392 991
rect 552 965 582 991
rect 638 965 668 991
rect 710 965 740 991
rect 80 351 110 565
rect 178 425 208 565
rect 264 499 294 565
rect 154 409 208 425
rect 154 375 164 409
rect 198 375 208 409
rect 154 359 208 375
rect 43 335 110 351
rect 43 301 53 335
rect 87 301 110 335
rect 43 285 110 301
rect 80 243 110 285
rect 178 243 208 359
rect 250 483 304 499
rect 250 449 260 483
rect 294 449 304 483
rect 250 433 304 449
rect 362 497 392 565
rect 552 497 582 565
rect 362 467 582 497
rect 250 243 280 433
rect 362 372 392 467
rect 638 425 668 565
rect 710 499 740 565
rect 710 483 764 499
rect 710 449 720 483
rect 754 449 764 483
rect 710 433 764 449
rect 338 356 392 372
rect 614 409 668 425
rect 614 375 624 409
rect 658 375 668 409
rect 614 359 668 375
rect 338 322 348 356
rect 382 328 392 356
rect 382 322 570 328
rect 338 298 570 322
rect 338 293 377 298
rect 442 283 472 298
rect 540 283 570 298
rect 626 283 656 359
rect 712 283 742 433
rect 80 89 110 115
rect 178 89 208 115
rect 250 89 280 115
rect 442 89 472 115
rect 540 89 570 115
rect 626 89 656 115
rect 712 89 742 115
<< polycont >>
rect 164 375 198 409
rect 53 301 87 335
rect 260 449 294 483
rect 720 449 754 483
rect 624 375 658 409
rect 348 322 382 356
<< locali >>
rect 0 1089 836 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 595 1089
rect 629 1049 731 1089
rect 765 1049 836 1089
rect 35 949 69 965
rect 35 575 69 597
rect 133 949 167 1049
rect 133 593 167 609
rect 219 949 253 965
rect 219 567 253 677
rect 305 949 339 1049
rect 305 661 339 677
rect 403 949 437 965
rect 219 533 362 567
rect 260 483 294 499
rect 260 433 294 449
rect 148 375 164 409
rect 198 375 214 409
rect 328 372 362 533
rect 403 557 437 609
rect 507 949 541 965
rect 403 523 418 557
rect 328 356 382 372
rect 328 340 348 356
rect 37 301 53 335
rect 87 301 110 335
rect 291 322 348 340
rect 291 306 382 322
rect 35 224 69 226
rect 35 115 69 131
rect 133 224 167 249
rect 133 61 167 131
rect 291 224 325 306
rect 418 267 452 523
rect 507 555 541 609
rect 593 949 627 1049
rect 593 593 627 609
rect 751 949 785 965
rect 751 555 785 609
rect 507 521 785 555
rect 507 335 541 521
rect 704 449 720 483
rect 754 449 770 483
rect 608 375 624 409
rect 658 375 674 409
rect 541 301 667 335
rect 291 115 325 131
rect 397 233 452 267
rect 495 233 529 249
rect 397 115 431 131
rect 495 61 529 131
rect 581 233 615 249
rect 667 247 701 301
rect 667 163 701 179
rect 753 233 787 249
rect 581 129 615 131
rect 753 129 787 131
rect 581 95 787 129
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 836 61
rect 0 0 836 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 595 1083 629 1089
rect 595 1055 629 1083
rect 731 1083 765 1089
rect 731 1055 765 1083
rect 35 609 69 631
rect 35 597 69 609
rect 260 449 294 483
rect 164 375 198 409
rect 418 523 452 557
rect 110 301 144 335
rect 35 226 69 260
rect 720 449 754 483
rect 624 375 658 409
rect 507 301 541 335
rect 667 301 701 335
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
<< metal1 >>
rect 0 1089 836 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 595 1089
rect 629 1055 731 1089
rect 765 1055 836 1089
rect 0 1049 836 1055
rect 23 631 81 637
rect 23 597 35 631
rect 69 597 81 631
rect 23 591 81 597
rect 35 266 69 591
rect 406 557 464 563
rect 406 523 418 557
rect 452 523 486 557
rect 406 517 464 523
rect 248 483 306 489
rect 708 483 766 489
rect 248 449 260 483
rect 294 449 720 483
rect 754 449 766 483
rect 248 448 766 449
rect 248 443 306 448
rect 708 443 766 448
rect 152 410 210 415
rect 612 410 670 415
rect 152 409 670 410
rect 152 375 164 409
rect 198 375 624 409
rect 658 375 670 409
rect 152 369 210 375
rect 612 369 670 375
rect 98 335 156 341
rect 495 335 553 341
rect 655 335 713 341
rect 98 301 110 335
rect 144 301 507 335
rect 541 301 553 335
rect 633 301 667 335
rect 701 301 713 335
rect 98 295 156 301
rect 495 295 553 301
rect 655 295 713 301
rect 23 260 81 266
rect 23 226 35 260
rect 69 226 81 260
rect 23 220 81 226
rect 0 55 836 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 836 55
rect 0 0 836 21
<< labels >>
rlabel metal1 50 425 50 425 1 S
port 1 n
rlabel viali 737 466 737 466 1 A
port 2 n
rlabel viali 642 392 642 392 1 B
port 3 n
rlabel viali 435 540 435 540 1 CO
port 4 n
rlabel viali 684 318 684 318 1 CON
port 5 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
