* File: sky130_osu_sc_12T_ls__buf_l.spice
* Created: Fri Nov 12 15:35:38 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__buf_l.pex.spice"
.subckt sky130_osu_sc_12T_ls__buf_l  GND VDD A Y
* 
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NSHORT L=0.15
+ W=0.36 AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4 SA=75000.2
+ SB=75000.6 A=0.054 P=1.02 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1002_d N_GND_M1002_b NSHORT L=0.15
+ W=0.36 AD=0.0954 AS=0.0504 PD=1.25 PS=0.64 NRD=0 NRS=0 M=1 R=2.4 SA=75000.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_VDD_M1001_d N_VDD_M1001_b PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=2.50965 P=6.35
pX5_noxref noxref_6 A A PROBETYPE=1
pX6_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__buf_l.pxi.spice"
*
.ends
*
*
