* File: sky130_osu_sc_18T_ls__dffs_1.spice
* Created: Fri Nov 12 14:16:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_ls__dffs_1.pex.spice"
.subckt sky130_osu_sc_18T_ls__dffs_1  GND VDD SN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* VDD	VDD
* GND	GND
MM1015 A_110_115# N_SN_M1015_g N_A_27_115#_M1015_s N_GND_M1015_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1002 N_GND_M1002_d N_A_152_89#_M1002_g A_110_115# N_GND_M1015_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 A_386_115# N_D_M1003_g N_GND_M1003_s N_GND_M1015_b NSHORT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1024 N_A_152_89#_M1024_d N_A_428_89#_M1024_g A_386_115# N_GND_M1015_b NSHORT
+ L=0.15 W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1
+ R=6.66667 SA=75000.5 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1020 A_578_115# N_CK_M1020_g N_A_152_89#_M1024_d N_GND_M1015_b NSHORT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.1 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1022 N_GND_M1022_d N_A_27_115#_M1022_g A_578_115# N_GND_M1015_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.5
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1016 A_736_115# N_A_27_115#_M1016_g N_GND_M1022_d N_GND_M1015_b NSHORT L=0.15
+ W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1012 N_A_808_115#_M1012_d N_CK_M1012_g A_736_115# N_GND_M1015_b NSHORT L=0.15
+ W=1 AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1 R=6.66667
+ SA=75002.3 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1004 A_928_115# N_A_428_89#_M1004_g N_A_808_115#_M1012_d N_GND_M1015_b NSHORT
+ L=0.15 W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1
+ R=6.66667 SA=75002.9 SB=75001 A=0.15 P=2.3 MULT=1
MM1008 N_GND_M1008_d N_A_970_89#_M1008_g A_928_115# N_GND_M1015_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75003.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_428_89#_M1005_d N_CK_M1005_g N_GND_M1008_d N_GND_M1015_b NSHORT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 A_1276_115# N_A_808_115#_M1006_g N_A_970_89#_M1006_s N_GND_M1015_b NSHORT
+ L=0.15 W=0.74 AD=0.0777 AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1026 N_GND_M1026_d N_SN_M1026_g A_1276_115# N_GND_M1015_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_GND_M1010_d N_A_970_89#_M1010_g N_QN_M1010_s N_GND_M1015_b NSHORT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1027 N_Q_M1027_d N_QN_M1027_g N_GND_M1010_d N_GND_M1015_b NSHORT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1023 N_A_27_115#_M1023_d N_SN_M1023_g N_VDD_M1023_s N_VDD_M1023_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1009 N_VDD_M1009_d N_A_152_89#_M1009_g N_A_27_115#_M1023_d N_VDD_M1023_b
+ PHIGHVT L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1011 A_386_617# N_D_M1011_g N_VDD_M1011_s N_VDD_M1023_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.2
+ SB=75003.7 A=0.45 P=6.3 MULT=1
MM1013 N_A_152_89#_M1013_d N_CK_M1013_g A_386_617# N_VDD_M1023_b PHIGHVT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75000.5 SB=75003.3 A=0.45 P=6.3 MULT=1
MM1018 A_578_617# N_A_428_89#_M1018_g N_A_152_89#_M1013_d N_VDD_M1023_b PHIGHVT
+ L=0.15 W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75001.1 SB=75002.7 A=0.45 P=6.3 MULT=1
MM1017 N_VDD_M1017_d N_A_27_115#_M1017_g A_578_617# N_VDD_M1023_b PHIGHVT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.5
+ SB=75002.4 A=0.45 P=6.3 MULT=1
MM1007 A_736_617# N_A_27_115#_M1007_g N_VDD_M1017_d N_VDD_M1023_b PHIGHVT L=0.15
+ W=3 AD=0.315 AS=0.42 PD=3.21 PS=3.28 NRD=3.2702 NRS=0 M=1 R=20 SA=75001.9
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1025 N_A_808_115#_M1025_d N_A_428_89#_M1025_g A_736_617# N_VDD_M1023_b PHIGHVT
+ L=0.15 W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75002.3 SB=75001.6 A=0.45 P=6.3 MULT=1
MM1000 A_928_617# N_CK_M1000_g N_A_808_115#_M1025_d N_VDD_M1023_b PHIGHVT L=0.15
+ W=3 AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20
+ SA=75002.9 SB=75001 A=0.45 P=6.3 MULT=1
MM1028 N_VDD_M1028_d N_A_970_89#_M1028_g A_928_617# N_VDD_M1023_b PHIGHVT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75003.3
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1019 N_A_428_89#_M1019_d N_CK_M1019_g N_VDD_M1028_d N_VDD_M1023_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.7
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1014 N_A_970_89#_M1014_d N_A_808_115#_M1014_g N_VDD_M1014_s N_VDD_M1023_b
+ PHIGHVT L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1029 N_VDD_M1029_d N_SN_M1029_g N_A_970_89#_M1014_d N_VDD_M1023_b PHIGHVT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.6 SB=75000.2 A=0.3 P=4.3 MULT=1
MM1001 N_VDD_M1001_d N_A_970_89#_M1001_g N_QN_M1001_s N_VDD_M1023_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1021 N_Q_M1021_d N_QN_M1021_g N_VDD_M1001_d N_VDD_M1023_b PHIGHVT L=0.15 W=3
+ AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX30_noxref N_GND_M1015_b N_VDD_M1023_b NWDIODE A=33.269 P=25.11
pX31_noxref noxref_23 SN SN PROBETYPE=1
pX32_noxref noxref_24 D D PROBETYPE=1
pX33_noxref noxref_25 CK CK PROBETYPE=1
pX34_noxref noxref_26 QN QN PROBETYPE=1
pX35_noxref noxref_27 Q Q PROBETYPE=1
c_1463 A_736_617# 0 1.57671e-19 $X=3.68 $Y=3.085
*
.include "sky130_osu_sc_18T_ls__dffs_1.pxi.spice"
*
.ends
*
*
