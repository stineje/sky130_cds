* File: sky130_osu_sc_12T_hs__or2_l.pxi.spice
* Created: Fri Nov 12 15:13:08 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__OR2_L%GND N_GND_M1003_s N_GND_M1000_d N_GND_M1003_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_19_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_HS__OR2_L%GND
x_PM_SKY130_OSU_SC_12T_HS__OR2_L%VDD N_VDD_M1004_d N_VDD_M1002_b N_VDD_c_38_p
+ N_VDD_c_42_p N_VDD_c_46_p VDD N_VDD_c_39_p PM_SKY130_OSU_SC_12T_HS__OR2_L%VDD
x_PM_SKY130_OSU_SC_12T_HS__OR2_L%B N_B_M1003_g N_B_M1002_g N_B_c_63_n N_B_c_64_n
+ B PM_SKY130_OSU_SC_12T_HS__OR2_L%B
x_PM_SKY130_OSU_SC_12T_HS__OR2_L%A N_A_M1000_g N_A_M1004_g N_A_c_93_n N_A_c_94_n
+ A PM_SKY130_OSU_SC_12T_HS__OR2_L%A
x_PM_SKY130_OSU_SC_12T_HS__OR2_L%A_27_605# N_A_27_605#_M1003_d
+ N_A_27_605#_M1002_s N_A_27_605#_M1001_g N_A_27_605#_M1005_g
+ N_A_27_605#_c_134_n N_A_27_605#_c_135_n N_A_27_605#_c_136_n
+ N_A_27_605#_c_148_n N_A_27_605#_c_151_n N_A_27_605#_c_152_n
+ N_A_27_605#_c_137_n N_A_27_605#_c_138_n N_A_27_605#_c_141_n
+ N_A_27_605#_c_142_n PM_SKY130_OSU_SC_12T_HS__OR2_L%A_27_605#
x_PM_SKY130_OSU_SC_12T_HS__OR2_L%Y N_Y_M1001_d N_Y_M1005_d N_Y_c_205_n
+ N_Y_c_208_n Y N_Y_c_210_n N_Y_c_211_n PM_SKY130_OSU_SC_12T_HS__OR2_L%Y
cc_1 N_GND_M1003_b N_B_M1003_g 0.121689f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.785
cc_2 N_GND_c_2_p N_B_M1003_g 0.00502587f $X=0.26 $Y=0.74 $X2=0.475 $Y2=0.785
cc_3 N_GND_c_3_p N_B_M1003_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.785
cc_4 N_GND_c_4_p N_B_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.785
cc_5 N_GND_M1003_b N_B_M1002_g 0.00488741f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.445
cc_6 N_GND_M1003_b N_B_c_63_n 0.0489195f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.565
cc_7 N_GND_M1003_b N_B_c_64_n 0.00390591f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.48
cc_8 N_GND_M1003_b B 0.0195655f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.48
cc_9 N_GND_M1003_b N_A_M1000_g 0.0693758f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.785
cc_10 N_GND_c_3_p N_A_M1000_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.785
cc_11 N_GND_c_11_p N_A_M1000_g 0.00308284f $X=1.12 $Y=0.74 $X2=0.905 $Y2=0.785
cc_12 N_GND_c_4_p N_A_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=0.785
cc_13 N_GND_M1003_b N_A_M1004_g 0.0177825f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.445
cc_14 N_GND_M1003_b N_A_c_93_n 0.0271998f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.275
cc_15 N_GND_M1003_b N_A_c_94_n 0.0021261f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.275
cc_16 N_GND_M1003_b A 0.0126158f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.48
cc_17 N_GND_M1003_b N_A_27_605#_M1001_g 0.0568175f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.785
cc_18 N_GND_c_11_p N_A_27_605#_M1001_g 0.00308284f $X=1.12 $Y=0.74 $X2=1.335
+ $Y2=0.785
cc_19 N_GND_c_19_p N_A_27_605#_M1001_g 0.00606474f $X=1.12 $Y=0.152 $X2=1.335
+ $Y2=0.785
cc_20 N_GND_c_4_p N_A_27_605#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=0.785
cc_21 N_GND_M1003_b N_A_27_605#_c_134_n 0.0364586f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=1.99
cc_22 N_GND_M1003_b N_A_27_605#_c_135_n 0.046655f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.7
cc_23 N_GND_M1003_b N_A_27_605#_c_136_n 0.0076832f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.835
cc_24 N_GND_M1003_b N_A_27_605#_c_137_n 0.00626981f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=2.935
cc_25 N_GND_M1003_b N_A_27_605#_c_138_n 0.0185591f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.74
cc_26 N_GND_c_3_p N_A_27_605#_c_138_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.74
cc_27 N_GND_c_4_p N_A_27_605#_c_138_n 0.00475776f $X=1.02 $Y=0.19 $X2=0.69
+ $Y2=0.74
cc_28 N_GND_M1003_b N_A_27_605#_c_141_n 0.0208326f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.825
cc_29 N_GND_M1003_b N_A_27_605#_c_142_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.825
cc_30 N_GND_M1003_b N_Y_c_205_n 0.0220167f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.74
cc_31 N_GND_c_19_p N_Y_c_205_n 0.00757793f $X=1.12 $Y=0.152 $X2=1.55 $Y2=0.74
cc_32 N_GND_c_4_p N_Y_c_205_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.74
cc_33 N_GND_M1003_b N_Y_c_208_n 0.0168357f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.48
cc_34 N_GND_M1003_b Y 0.039938f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.11
cc_35 N_GND_M1003_b N_Y_c_210_n 0.0157042f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.37
cc_36 N_GND_M1003_b N_Y_c_211_n 0.0141689f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.48
cc_37 N_VDD_M1002_b N_B_M1002_g 0.0303911f $X=-0.045 $Y=2.795 $X2=0.475
+ $Y2=3.445
cc_38 N_VDD_c_38_p N_B_M1002_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.445
cc_39 N_VDD_c_39_p N_B_M1002_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.445
cc_40 N_VDD_M1002_b N_A_M1004_g 0.0232721f $X=-0.045 $Y=2.795 $X2=0.905
+ $Y2=3.445
cc_41 N_VDD_c_38_p N_A_M1004_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.445
cc_42 N_VDD_c_42_p N_A_M1004_g 0.00354579f $X=1.12 $Y=3.615 $X2=0.905 $Y2=3.445
cc_43 N_VDD_c_39_p N_A_M1004_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.905 $Y2=3.445
cc_44 N_VDD_M1002_b N_A_27_605#_M1005_g 0.0251486f $X=-0.045 $Y=2.795 $X2=1.335
+ $Y2=3.445
cc_45 N_VDD_c_42_p N_A_27_605#_M1005_g 0.00354579f $X=1.12 $Y=3.615 $X2=1.335
+ $Y2=3.445
cc_46 N_VDD_c_46_p N_A_27_605#_M1005_g 0.00606474f $X=1.12 $Y=4.287 $X2=1.335
+ $Y2=3.445
cc_47 N_VDD_c_39_p N_A_27_605#_M1005_g 0.00468827f $X=1.02 $Y=4.25 $X2=1.335
+ $Y2=3.445
cc_48 N_VDD_M1002_b N_A_27_605#_c_136_n 0.00435501f $X=-0.045 $Y=2.795 $X2=1.352
+ $Y2=2.835
cc_49 N_VDD_M1002_b N_A_27_605#_c_148_n 0.00156053f $X=-0.045 $Y=2.795 $X2=0.26
+ $Y2=3.615
cc_50 N_VDD_c_38_p N_A_27_605#_c_148_n 0.00736239f $X=1.035 $Y=4.287 $X2=0.26
+ $Y2=3.615
cc_51 N_VDD_c_39_p N_A_27_605#_c_148_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26
+ $Y2=3.615
cc_52 N_VDD_M1002_b N_A_27_605#_c_151_n 0.00118949f $X=-0.045 $Y=2.795 $X2=0.525
+ $Y2=3.02
cc_53 N_VDD_M1002_b N_A_27_605#_c_152_n 0.00466538f $X=-0.045 $Y=2.795 $X2=0.345
+ $Y2=3.02
cc_54 N_VDD_M1002_b N_A_27_605#_c_137_n 0.00130531f $X=-0.045 $Y=2.795 $X2=0.61
+ $Y2=2.935
cc_55 N_VDD_M1002_b N_Y_c_208_n 0.0129685f $X=-0.045 $Y=2.795 $X2=1.55 $Y2=2.48
cc_56 N_VDD_c_46_p N_Y_c_208_n 0.00757793f $X=1.12 $Y=4.287 $X2=1.55 $Y2=2.48
cc_57 N_VDD_c_39_p N_Y_c_208_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.55 $Y2=2.48
cc_58 N_B_M1003_g N_A_M1000_g 0.0492988f $X=0.475 $Y=0.785 $X2=0.905 $Y2=0.785
cc_59 N_B_c_63_n N_A_M1004_g 0.0670255f $X=0.475 $Y=2.565 $X2=0.905 $Y2=3.445
cc_60 N_B_M1003_g N_A_c_93_n 0.0153344f $X=0.475 $Y=0.785 $X2=0.95 $Y2=2.275
cc_61 N_B_M1003_g N_A_c_94_n 5.05199e-19 $X=0.475 $Y=0.785 $X2=0.95 $Y2=2.275
cc_62 B A 0.0170852f $X=0.27 $Y=2.48 $X2=0.95 $Y2=2.48
cc_63 N_B_M1002_g N_A_27_605#_c_151_n 0.0158924f $X=0.475 $Y=3.445 $X2=0.525
+ $Y2=3.02
cc_64 N_B_c_63_n N_A_27_605#_c_151_n 0.00172264f $X=0.475 $Y=2.565 $X2=0.525
+ $Y2=3.02
cc_65 N_B_c_64_n N_A_27_605#_c_151_n 5.12056e-19 $X=0.27 $Y=2.48 $X2=0.525
+ $Y2=3.02
cc_66 B N_A_27_605#_c_151_n 0.00560865f $X=0.27 $Y=2.48 $X2=0.525 $Y2=3.02
cc_67 N_B_c_63_n N_A_27_605#_c_152_n 0.00169997f $X=0.475 $Y=2.565 $X2=0.345
+ $Y2=3.02
cc_68 N_B_c_64_n N_A_27_605#_c_152_n 0.0105955f $X=0.27 $Y=2.48 $X2=0.345
+ $Y2=3.02
cc_69 B N_A_27_605#_c_152_n 0.00146821f $X=0.27 $Y=2.48 $X2=0.345 $Y2=3.02
cc_70 N_B_M1003_g N_A_27_605#_c_137_n 0.0222319f $X=0.475 $Y=0.785 $X2=0.61
+ $Y2=2.935
cc_71 N_B_M1002_g N_A_27_605#_c_137_n 0.00967013f $X=0.475 $Y=3.445 $X2=0.61
+ $Y2=2.935
cc_72 N_B_c_63_n N_A_27_605#_c_137_n 0.00750666f $X=0.475 $Y=2.565 $X2=0.61
+ $Y2=2.935
cc_73 N_B_c_64_n N_A_27_605#_c_137_n 0.0208906f $X=0.27 $Y=2.48 $X2=0.61
+ $Y2=2.935
cc_74 B N_A_27_605#_c_137_n 0.00282146f $X=0.27 $Y=2.48 $X2=0.61 $Y2=2.935
cc_75 N_B_M1003_g N_A_27_605#_c_138_n 0.0179929f $X=0.475 $Y=0.785 $X2=0.69
+ $Y2=0.74
cc_76 N_B_M1003_g N_A_27_605#_c_142_n 0.0113001f $X=0.475 $Y=0.785 $X2=0.65
+ $Y2=1.825
cc_77 N_A_M1000_g N_A_27_605#_M1001_g 0.0423877f $X=0.905 $Y=0.785 $X2=1.335
+ $Y2=0.785
cc_78 N_A_M1000_g N_A_27_605#_c_134_n 0.0119161f $X=0.905 $Y=0.785 $X2=1.37
+ $Y2=1.99
cc_79 N_A_M1004_g N_A_27_605#_c_135_n 0.00948064f $X=0.905 $Y=3.445 $X2=1.352
+ $Y2=2.7
cc_80 N_A_c_93_n N_A_27_605#_c_135_n 0.0206139f $X=0.95 $Y=2.275 $X2=1.352
+ $Y2=2.7
cc_81 N_A_c_94_n N_A_27_605#_c_135_n 0.00278895f $X=0.95 $Y=2.275 $X2=1.352
+ $Y2=2.7
cc_82 A N_A_27_605#_c_135_n 0.00109846f $X=0.95 $Y=2.48 $X2=1.352 $Y2=2.7
cc_83 N_A_M1004_g N_A_27_605#_c_136_n 0.0377642f $X=0.905 $Y=3.445 $X2=1.352
+ $Y2=2.835
cc_84 N_A_M1004_g N_A_27_605#_c_151_n 0.00457566f $X=0.905 $Y=3.445 $X2=0.525
+ $Y2=3.02
cc_85 N_A_M1000_g N_A_27_605#_c_137_n 0.00429604f $X=0.905 $Y=0.785 $X2=0.61
+ $Y2=2.935
cc_86 N_A_M1004_g N_A_27_605#_c_137_n 0.00860585f $X=0.905 $Y=3.445 $X2=0.61
+ $Y2=2.935
cc_87 N_A_c_93_n N_A_27_605#_c_137_n 0.00205758f $X=0.95 $Y=2.275 $X2=0.61
+ $Y2=2.935
cc_88 N_A_c_94_n N_A_27_605#_c_137_n 0.030681f $X=0.95 $Y=2.275 $X2=0.61
+ $Y2=2.935
cc_89 A N_A_27_605#_c_137_n 0.00287859f $X=0.95 $Y=2.48 $X2=0.61 $Y2=2.935
cc_90 N_A_M1000_g N_A_27_605#_c_138_n 0.0179929f $X=0.905 $Y=0.785 $X2=0.69
+ $Y2=0.74
cc_91 N_A_M1000_g N_A_27_605#_c_141_n 0.0154849f $X=0.905 $Y=0.785 $X2=1.43
+ $Y2=1.825
cc_92 N_A_c_93_n N_A_27_605#_c_141_n 0.00276813f $X=0.95 $Y=2.275 $X2=1.43
+ $Y2=1.825
cc_93 N_A_c_94_n N_A_27_605#_c_141_n 0.0104443f $X=0.95 $Y=2.275 $X2=1.43
+ $Y2=1.825
cc_94 A N_A_27_605#_c_141_n 0.00820853f $X=0.95 $Y=2.48 $X2=1.43 $Y2=1.825
cc_95 N_A_c_94_n N_Y_c_208_n 0.00445016f $X=0.95 $Y=2.275 $X2=1.55 $Y2=2.48
cc_96 A N_Y_c_208_n 9.44517e-19 $X=0.95 $Y=2.48 $X2=1.55 $Y2=2.48
cc_97 N_A_M1000_g Y 6.73508e-19 $X=0.905 $Y=0.785 $X2=1.555 $Y2=2.11
cc_98 N_A_c_94_n Y 0.00825539f $X=0.95 $Y=2.275 $X2=1.555 $Y2=2.11
cc_99 N_A_M1000_g N_Y_c_210_n 0.00102215f $X=0.905 $Y=0.785 $X2=1.55 $Y2=1.37
cc_100 N_A_c_94_n N_Y_c_211_n 9.31495e-19 $X=0.95 $Y=2.275 $X2=1.55 $Y2=2.48
cc_101 A N_Y_c_211_n 0.0197623f $X=0.95 $Y=2.48 $X2=1.55 $Y2=2.48
cc_102 N_A_27_605#_c_151_n A_110_605# 0.00500895f $X=0.525 $Y=3.02 $X2=0.55
+ $Y2=3.025
cc_103 N_A_27_605#_M1001_g N_Y_c_205_n 0.0178582f $X=1.335 $Y=0.785 $X2=1.55
+ $Y2=0.74
cc_104 N_A_27_605#_c_134_n N_Y_c_205_n 0.00168f $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=0.74
cc_105 N_A_27_605#_c_141_n N_Y_c_205_n 0.00530006f $X=1.43 $Y=1.825 $X2=1.55
+ $Y2=0.74
cc_106 N_A_27_605#_M1005_g N_Y_c_208_n 0.0159552f $X=1.335 $Y=3.445 $X2=1.55
+ $Y2=2.48
cc_107 N_A_27_605#_c_134_n N_Y_c_208_n 0.00125776f $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=2.48
cc_108 N_A_27_605#_c_135_n N_Y_c_208_n 0.0148241f $X=1.352 $Y=2.7 $X2=1.55
+ $Y2=2.48
cc_109 N_A_27_605#_c_141_n N_Y_c_208_n 0.00273485f $X=1.43 $Y=1.825 $X2=1.55
+ $Y2=2.48
cc_110 N_A_27_605#_M1001_g Y 0.00406656f $X=1.335 $Y=0.785 $X2=1.555 $Y2=2.11
cc_111 N_A_27_605#_c_134_n Y 0.00704613f $X=1.37 $Y=1.99 $X2=1.555 $Y2=2.11
cc_112 N_A_27_605#_c_135_n Y 0.00892438f $X=1.352 $Y=2.7 $X2=1.555 $Y2=2.11
cc_113 N_A_27_605#_c_141_n Y 0.0151477f $X=1.43 $Y=1.825 $X2=1.555 $Y2=2.11
cc_114 N_A_27_605#_M1001_g N_Y_c_210_n 0.00715333f $X=1.335 $Y=0.785 $X2=1.55
+ $Y2=1.37
cc_115 N_A_27_605#_c_134_n N_Y_c_210_n 0.00154864f $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=1.37
cc_116 N_A_27_605#_c_141_n N_Y_c_210_n 0.00238892f $X=1.43 $Y=1.825 $X2=1.55
+ $Y2=1.37
cc_117 N_A_27_605#_c_134_n N_Y_c_211_n 4.58687e-19 $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=2.48
cc_118 N_A_27_605#_c_135_n N_Y_c_211_n 0.00579834f $X=1.352 $Y=2.7 $X2=1.55
+ $Y2=2.48
cc_119 N_A_27_605#_c_141_n N_Y_c_211_n 0.00181779f $X=1.43 $Y=1.825 $X2=1.55
+ $Y2=2.48
