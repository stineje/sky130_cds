* File: sky130_osu_sc_12T_ls__buf_8.pxi.spice
* Created: Fri Nov 12 15:35:30 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__BUF_8%GND N_GND_M1007_d N_GND_M1001_s N_GND_M1010_s
+ N_GND_M1013_s N_GND_M1017_s N_GND_M1007_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p
+ N_GND_c_15_p N_GND_c_24_p N_GND_c_30_p N_GND_c_37_p N_GND_c_44_p N_GND_c_51_p
+ N_GND_c_57_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_LS__BUF_8%GND
x_PM_SKY130_OSU_SC_12T_LS__BUF_8%VDD N_VDD_M1005_d N_VDD_M1003_s N_VDD_M1006_s
+ N_VDD_M1011_s N_VDD_M1016_s N_VDD_M1005_b N_VDD_c_131_p N_VDD_c_132_p
+ N_VDD_c_141_p N_VDD_c_146_p N_VDD_c_153_p N_VDD_c_158_p N_VDD_c_164_p
+ N_VDD_c_169_p N_VDD_c_175_p N_VDD_c_180_p VDD N_VDD_c_133_p
+ PM_SKY130_OSU_SC_12T_LS__BUF_8%VDD
x_PM_SKY130_OSU_SC_12T_LS__BUF_8%A N_A_M1007_g N_A_M1005_g N_A_c_217_n
+ N_A_c_218_n A PM_SKY130_OSU_SC_12T_LS__BUF_8%A
x_PM_SKY130_OSU_SC_12T_LS__BUF_8%A_27_115# N_A_27_115#_M1007_s
+ N_A_27_115#_M1005_s N_A_27_115#_M1000_g N_A_27_115#_c_321_n
+ N_A_27_115#_M1002_g N_A_27_115#_c_256_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_325_n N_A_27_115#_M1003_g N_A_27_115#_c_261_n
+ N_A_27_115#_c_263_n N_A_27_115#_c_264_n N_A_27_115#_c_265_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_333_n N_A_27_115#_M1004_g
+ N_A_27_115#_c_270_n N_A_27_115#_c_271_n N_A_27_115#_M1010_g
+ N_A_27_115#_c_338_n N_A_27_115#_M1006_g N_A_27_115#_c_276_n
+ N_A_27_115#_c_278_n N_A_27_115#_M1012_g N_A_27_115#_c_283_n
+ N_A_27_115#_c_344_n N_A_27_115#_M1009_g N_A_27_115#_c_284_n
+ N_A_27_115#_c_285_n N_A_27_115#_M1013_g N_A_27_115#_c_349_n
+ N_A_27_115#_M1011_g N_A_27_115#_c_290_n N_A_27_115#_c_292_n
+ N_A_27_115#_M1014_g N_A_27_115#_c_355_n N_A_27_115#_M1015_g
+ N_A_27_115#_c_297_n N_A_27_115#_c_298_n N_A_27_115#_M1017_g
+ N_A_27_115#_c_360_n N_A_27_115#_M1016_g N_A_27_115#_c_303_n
+ N_A_27_115#_c_304_n N_A_27_115#_c_305_n N_A_27_115#_c_306_n
+ N_A_27_115#_c_307_n N_A_27_115#_c_308_n N_A_27_115#_c_309_n
+ N_A_27_115#_c_310_n N_A_27_115#_c_311_n N_A_27_115#_c_312_n
+ N_A_27_115#_c_313_n N_A_27_115#_c_316_n N_A_27_115#_c_317_n
+ N_A_27_115#_c_319_n N_A_27_115#_c_320_n
+ PM_SKY130_OSU_SC_12T_LS__BUF_8%A_27_115#
x_PM_SKY130_OSU_SC_12T_LS__BUF_8%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1012_d
+ N_Y_M1014_d N_Y_M1002_d N_Y_M1004_d N_Y_M1009_d N_Y_M1015_d N_Y_c_484_n
+ N_Y_c_537_n N_Y_c_488_n N_Y_c_540_n N_Y_c_493_n N_Y_c_543_n N_Y_c_498_n
+ N_Y_c_546_n N_Y_c_502_n N_Y_c_506_n Y N_Y_c_508_n N_Y_c_550_n N_Y_c_512_n
+ N_Y_c_513_n N_Y_c_517_n N_Y_c_552_n N_Y_c_521_n N_Y_c_522_n N_Y_c_523_n
+ N_Y_c_527_n N_Y_c_555_n N_Y_c_531_n N_Y_c_532_n N_Y_c_536_n
+ PM_SKY130_OSU_SC_12T_LS__BUF_8%Y
cc_1 N_GND_M1007_b N_A_M1007_g 0.0588914f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1007_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_A_M1007_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.475 $Y2=0.835
cc_4 N_GND_c_4_p N_A_M1007_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.475 $Y2=0.835
cc_5 N_GND_M1007_b N_A_M1005_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_6 N_GND_M1007_b N_A_c_217_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_7 N_GND_M1007_b N_A_c_218_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2
cc_8 N_GND_M1007_b N_A_27_115#_M1000_g 0.0207501f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.835
cc_9 N_GND_c_3_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.755 $X2=0.905
+ $Y2=0.835
cc_10 N_GND_c_10_p N_A_27_115#_M1000_g 0.00606474f $X=1.465 $Y=0.152 $X2=0.905
+ $Y2=0.835
cc_11 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.905
+ $Y2=0.835
cc_12 N_GND_M1007_b N_A_27_115#_c_256_n 0.0479182f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.38
cc_13 N_GND_M1007_b N_A_27_115#_M1001_g 0.020212f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.835
cc_14 N_GND_c_10_p N_A_27_115#_M1001_g 0.00606474f $X=1.465 $Y=0.152 $X2=1.335
+ $Y2=0.835
cc_15 N_GND_c_15_p N_A_27_115#_M1001_g 0.00311745f $X=1.55 $Y=0.755 $X2=1.335
+ $Y2=0.835
cc_16 N_GND_c_4_p N_A_27_115#_M1001_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.335
+ $Y2=0.835
cc_17 N_GND_M1007_b N_A_27_115#_c_261_n 0.0215078f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=1.365
cc_18 N_GND_c_15_p N_A_27_115#_c_261_n 0.00256938f $X=1.55 $Y=0.755 $X2=1.69
+ $Y2=1.365
cc_19 N_GND_M1007_b N_A_27_115#_c_263_n 0.0429274f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=1.365
cc_20 N_GND_M1007_b N_A_27_115#_c_264_n 0.0158747f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.455
cc_21 N_GND_M1007_b N_A_27_115#_c_265_n 0.0196789f $X=-0.045 $Y=0 $X2=1.41
+ $Y2=2.455
cc_22 N_GND_M1007_b N_A_27_115#_M1008_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.835
cc_23 N_GND_c_15_p N_A_27_115#_M1008_g 0.00311745f $X=1.55 $Y=0.755 $X2=1.765
+ $Y2=0.835
cc_24 N_GND_c_24_p N_A_27_115#_M1008_g 0.00606474f $X=2.325 $Y=0.152 $X2=1.765
+ $Y2=0.835
cc_25 N_GND_c_4_p N_A_27_115#_M1008_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.765
+ $Y2=0.835
cc_26 N_GND_M1007_b N_A_27_115#_c_270_n 0.0195339f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.365
cc_27 N_GND_M1007_b N_A_27_115#_c_271_n 0.0107618f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.455
cc_28 N_GND_M1007_b N_A_27_115#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.835
cc_29 N_GND_c_24_p N_A_27_115#_M1010_g 0.00606474f $X=2.325 $Y=0.152 $X2=2.195
+ $Y2=0.835
cc_30 N_GND_c_30_p N_A_27_115#_M1010_g 0.00311745f $X=2.41 $Y=0.755 $X2=2.195
+ $Y2=0.835
cc_31 N_GND_c_4_p N_A_27_115#_M1010_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.195
+ $Y2=0.835
cc_32 N_GND_M1007_b N_A_27_115#_c_276_n 0.0165886f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.365
cc_33 N_GND_c_30_p N_A_27_115#_c_276_n 0.00256938f $X=2.41 $Y=0.755 $X2=2.55
+ $Y2=1.365
cc_34 N_GND_M1007_b N_A_27_115#_c_278_n 0.0109555f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.455
cc_35 N_GND_M1007_b N_A_27_115#_M1012_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.835
cc_36 N_GND_c_30_p N_A_27_115#_M1012_g 0.00311745f $X=2.41 $Y=0.755 $X2=2.625
+ $Y2=0.835
cc_37 N_GND_c_37_p N_A_27_115#_M1012_g 0.00606474f $X=3.185 $Y=0.152 $X2=2.625
+ $Y2=0.835
cc_38 N_GND_c_4_p N_A_27_115#_M1012_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.625
+ $Y2=0.835
cc_39 N_GND_M1007_b N_A_27_115#_c_283_n 0.0668243f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.38
cc_40 N_GND_M1007_b N_A_27_115#_c_284_n 0.0195339f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.365
cc_41 N_GND_M1007_b N_A_27_115#_c_285_n 0.0107618f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.455
cc_42 N_GND_M1007_b N_A_27_115#_M1013_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.835
cc_43 N_GND_c_37_p N_A_27_115#_M1013_g 0.00606474f $X=3.185 $Y=0.152 $X2=3.055
+ $Y2=0.835
cc_44 N_GND_c_44_p N_A_27_115#_M1013_g 0.00311745f $X=3.27 $Y=0.755 $X2=3.055
+ $Y2=0.835
cc_45 N_GND_c_4_p N_A_27_115#_M1013_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.055
+ $Y2=0.835
cc_46 N_GND_M1007_b N_A_27_115#_c_290_n 0.0215078f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.365
cc_47 N_GND_c_44_p N_A_27_115#_c_290_n 0.00256938f $X=3.27 $Y=0.755 $X2=3.41
+ $Y2=1.365
cc_48 N_GND_M1007_b N_A_27_115#_c_292_n 0.0158747f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.455
cc_49 N_GND_M1007_b N_A_27_115#_M1014_g 0.020212f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=0.835
cc_50 N_GND_c_44_p N_A_27_115#_M1014_g 0.00311745f $X=3.27 $Y=0.755 $X2=3.485
+ $Y2=0.835
cc_51 N_GND_c_51_p N_A_27_115#_M1014_g 0.00606474f $X=4.045 $Y=0.152 $X2=3.485
+ $Y2=0.835
cc_52 N_GND_c_4_p N_A_27_115#_M1014_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.485
+ $Y2=0.835
cc_53 N_GND_M1007_b N_A_27_115#_c_297_n 0.0385034f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.365
cc_54 N_GND_M1007_b N_A_27_115#_c_298_n 0.0221499f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.455
cc_55 N_GND_M1007_b N_A_27_115#_M1017_g 0.0264941f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=0.835
cc_56 N_GND_c_51_p N_A_27_115#_M1017_g 0.00606474f $X=4.045 $Y=0.152 $X2=3.915
+ $Y2=0.835
cc_57 N_GND_c_57_p N_A_27_115#_M1017_g 0.00502587f $X=4.13 $Y=0.755 $X2=3.915
+ $Y2=0.835
cc_58 N_GND_c_4_p N_A_27_115#_M1017_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.915
+ $Y2=0.835
cc_59 N_GND_M1007_b N_A_27_115#_c_303_n 0.0106787f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.365
cc_60 N_GND_M1007_b N_A_27_115#_c_304_n 0.00890086f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.455
cc_61 N_GND_M1007_b N_A_27_115#_c_305_n 0.0106787f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.365
cc_62 N_GND_M1007_b N_A_27_115#_c_306_n 0.00890086f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.455
cc_63 N_GND_M1007_b N_A_27_115#_c_307_n 0.0023879f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.365
cc_64 N_GND_M1007_b N_A_27_115#_c_308_n 7.16371e-19 $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.455
cc_65 N_GND_M1007_b N_A_27_115#_c_309_n 0.0106787f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.365
cc_66 N_GND_M1007_b N_A_27_115#_c_310_n 0.00890086f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.455
cc_67 N_GND_M1007_b N_A_27_115#_c_311_n 0.0106787f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.365
cc_68 N_GND_M1007_b N_A_27_115#_c_312_n 0.00890086f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.455
cc_69 N_GND_M1007_b N_A_27_115#_c_313_n 0.0142265f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_70 N_GND_c_2_p N_A_27_115#_c_313_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_71 N_GND_c_4_p N_A_27_115#_c_313_n 0.00476261f $X=3.74 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_72 N_GND_M1007_b N_A_27_115#_c_316_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=2.955
cc_73 N_GND_M1007_b N_A_27_115#_c_317_n 0.013728f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.455
cc_74 N_GND_c_3_p N_A_27_115#_c_317_n 0.00702738f $X=0.69 $Y=0.755 $X2=0.88
+ $Y2=1.455
cc_75 N_GND_M1007_b N_A_27_115#_c_319_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.455
cc_76 N_GND_M1007_b N_A_27_115#_c_320_n 0.00592383f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.455
cc_77 N_GND_M1007_b N_Y_c_484_n 0.00154299f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.755
cc_78 N_GND_c_10_p N_Y_c_484_n 0.00718527f $X=1.465 $Y=0.152 $X2=1.12 $Y2=0.755
cc_79 N_GND_c_15_p N_Y_c_484_n 8.14297e-19 $X=1.55 $Y=0.755 $X2=1.12 $Y2=0.755
cc_80 N_GND_c_4_p N_Y_c_484_n 0.0047139f $X=3.74 $Y=0.19 $X2=1.12 $Y2=0.755
cc_81 N_GND_M1007_b N_Y_c_488_n 0.00154299f $X=-0.045 $Y=0 $X2=1.98 $Y2=0.755
cc_82 N_GND_c_15_p N_Y_c_488_n 8.14297e-19 $X=1.55 $Y=0.755 $X2=1.98 $Y2=0.755
cc_83 N_GND_c_24_p N_Y_c_488_n 0.00738926f $X=2.325 $Y=0.152 $X2=1.98 $Y2=0.755
cc_84 N_GND_c_30_p N_Y_c_488_n 8.14297e-19 $X=2.41 $Y=0.755 $X2=1.98 $Y2=0.755
cc_85 N_GND_c_4_p N_Y_c_488_n 0.0047139f $X=3.74 $Y=0.19 $X2=1.98 $Y2=0.755
cc_86 N_GND_M1007_b N_Y_c_493_n 0.00154299f $X=-0.045 $Y=0 $X2=2.84 $Y2=0.755
cc_87 N_GND_c_30_p N_Y_c_493_n 8.14297e-19 $X=2.41 $Y=0.755 $X2=2.84 $Y2=0.755
cc_88 N_GND_c_37_p N_Y_c_493_n 0.00731228f $X=3.185 $Y=0.152 $X2=2.84 $Y2=0.755
cc_89 N_GND_c_44_p N_Y_c_493_n 8.14297e-19 $X=3.27 $Y=0.755 $X2=2.84 $Y2=0.755
cc_90 N_GND_c_4_p N_Y_c_493_n 0.0047139f $X=3.74 $Y=0.19 $X2=2.84 $Y2=0.755
cc_91 N_GND_M1007_b N_Y_c_498_n 0.00154299f $X=-0.045 $Y=0 $X2=3.7 $Y2=0.755
cc_92 N_GND_c_44_p N_Y_c_498_n 8.14297e-19 $X=3.27 $Y=0.755 $X2=3.7 $Y2=0.755
cc_93 N_GND_c_51_p N_Y_c_498_n 0.00718527f $X=4.045 $Y=0.152 $X2=3.7 $Y2=0.755
cc_94 N_GND_c_4_p N_Y_c_498_n 0.0047139f $X=3.74 $Y=0.19 $X2=3.7 $Y2=0.755
cc_95 N_GND_M1007_b N_Y_c_502_n 0.00244441f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.115
cc_96 N_GND_c_3_p N_Y_c_502_n 0.00134236f $X=0.69 $Y=0.755 $X2=1.12 $Y2=1.115
cc_97 N_GND_c_10_p N_Y_c_502_n 0.00245319f $X=1.465 $Y=0.152 $X2=1.12 $Y2=1.115
cc_98 N_GND_c_15_p N_Y_c_502_n 7.53951e-19 $X=1.55 $Y=0.755 $X2=1.12 $Y2=1.115
cc_99 N_GND_M1007_b N_Y_c_506_n 0.00329802f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.365
cc_100 N_GND_M1007_b Y 0.0126399f $X=-0.045 $Y=0 $X2=1.055 $Y2=1.79
cc_101 N_GND_M1001_s N_Y_c_508_n 0.0100329f $X=1.41 $Y=0.575 $X2=1.835 $Y2=1
cc_102 N_GND_c_10_p N_Y_c_508_n 0.0028844f $X=1.465 $Y=0.152 $X2=1.835 $Y2=1
cc_103 N_GND_c_15_p N_Y_c_508_n 0.0142303f $X=1.55 $Y=0.755 $X2=1.835 $Y2=1
cc_104 N_GND_c_24_p N_Y_c_508_n 0.0028844f $X=2.325 $Y=0.152 $X2=1.835 $Y2=1
cc_105 N_GND_M1007_b N_Y_c_512_n 0.0437239f $X=-0.045 $Y=0 $X2=1.98 $Y2=2.365
cc_106 N_GND_M1010_s N_Y_c_513_n 0.0100329f $X=2.27 $Y=0.575 $X2=2.695 $Y2=1
cc_107 N_GND_c_24_p N_Y_c_513_n 0.0028844f $X=2.325 $Y=0.152 $X2=2.695 $Y2=1
cc_108 N_GND_c_30_p N_Y_c_513_n 0.0142303f $X=2.41 $Y=0.755 $X2=2.695 $Y2=1
cc_109 N_GND_c_37_p N_Y_c_513_n 0.0028844f $X=3.185 $Y=0.152 $X2=2.695 $Y2=1
cc_110 N_GND_M1007_b N_Y_c_517_n 0.00409378f $X=-0.045 $Y=0 $X2=2.125 $Y2=1
cc_111 N_GND_c_15_p N_Y_c_517_n 7.53951e-19 $X=1.55 $Y=0.755 $X2=2.125 $Y2=1
cc_112 N_GND_c_24_p N_Y_c_517_n 0.00245319f $X=2.325 $Y=0.152 $X2=2.125 $Y2=1
cc_113 N_GND_c_30_p N_Y_c_517_n 7.53951e-19 $X=2.41 $Y=0.755 $X2=2.125 $Y2=1
cc_114 N_GND_M1007_b N_Y_c_521_n 0.00560779f $X=-0.045 $Y=0 $X2=2.125 $Y2=2.48
cc_115 N_GND_M1007_b N_Y_c_522_n 0.0575129f $X=-0.045 $Y=0 $X2=2.84 $Y2=2.365
cc_116 N_GND_M1013_s N_Y_c_523_n 0.0100329f $X=3.13 $Y=0.575 $X2=3.555 $Y2=1
cc_117 N_GND_c_37_p N_Y_c_523_n 0.0028844f $X=3.185 $Y=0.152 $X2=3.555 $Y2=1
cc_118 N_GND_c_44_p N_Y_c_523_n 0.0142303f $X=3.27 $Y=0.755 $X2=3.555 $Y2=1
cc_119 N_GND_c_51_p N_Y_c_523_n 0.0028844f $X=4.045 $Y=0.152 $X2=3.555 $Y2=1
cc_120 N_GND_M1007_b N_Y_c_527_n 0.00409378f $X=-0.045 $Y=0 $X2=2.985 $Y2=1
cc_121 N_GND_c_30_p N_Y_c_527_n 7.53951e-19 $X=2.41 $Y=0.755 $X2=2.985 $Y2=1
cc_122 N_GND_c_37_p N_Y_c_527_n 0.00245319f $X=3.185 $Y=0.152 $X2=2.985 $Y2=1
cc_123 N_GND_c_44_p N_Y_c_527_n 7.53951e-19 $X=3.27 $Y=0.755 $X2=2.985 $Y2=1
cc_124 N_GND_M1007_b N_Y_c_531_n 0.00485078f $X=-0.045 $Y=0 $X2=2.985 $Y2=2.48
cc_125 N_GND_M1007_b N_Y_c_532_n 0.00409378f $X=-0.045 $Y=0 $X2=3.7 $Y2=1.115
cc_126 N_GND_c_44_p N_Y_c_532_n 7.53951e-19 $X=3.27 $Y=0.755 $X2=3.7 $Y2=1.115
cc_127 N_GND_c_51_p N_Y_c_532_n 0.00245319f $X=4.045 $Y=0.152 $X2=3.7 $Y2=1.115
cc_128 N_GND_c_57_p N_Y_c_532_n 0.00134236f $X=4.13 $Y=0.755 $X2=3.7 $Y2=1.115
cc_129 N_GND_M1007_b N_Y_c_536_n 0.0800785f $X=-0.045 $Y=0 $X2=3.7 $Y2=2.365
cc_130 N_VDD_M1005_b N_A_M1005_g 0.0245629f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_131 N_VDD_c_131_p N_A_M1005_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_132 N_VDD_c_132_p N_A_M1005_g 0.00337744f $X=0.69 $Y=3.635 $X2=0.475
+ $Y2=3.235
cc_133 N_VDD_c_133_p N_A_M1005_g 0.00468827f $X=3.74 $Y=4.25 $X2=0.475 $Y2=3.235
cc_134 N_VDD_M1005_d N_A_c_218_n 0.00628533f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2
cc_135 N_VDD_M1005_b N_A_c_218_n 0.00328912f $X=-0.045 $Y=2.425 $X2=0.635 $Y2=2
cc_136 N_VDD_c_132_p N_A_c_218_n 0.00264661f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2
cc_137 N_VDD_M1005_d A 0.00797576f $X=0.55 $Y=2.605 $X2=0.635 $Y2=2.85
cc_138 N_VDD_c_132_p A 0.00510982f $X=0.69 $Y=3.635 $X2=0.635 $Y2=2.85
cc_139 N_VDD_M1005_b N_A_27_115#_c_321_n 0.014249f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.53
cc_140 N_VDD_c_132_p N_A_27_115#_c_321_n 0.00337744f $X=0.69 $Y=3.635 $X2=0.905
+ $Y2=2.53
cc_141 N_VDD_c_141_p N_A_27_115#_c_321_n 0.00606474f $X=1.465 $Y=4.287 $X2=0.905
+ $Y2=2.53
cc_142 N_VDD_c_133_p N_A_27_115#_c_321_n 0.00468827f $X=3.74 $Y=4.25 $X2=0.905
+ $Y2=2.53
cc_143 N_VDD_M1005_b N_A_27_115#_c_325_n 0.0141063f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.53
cc_144 N_VDD_c_132_p N_A_27_115#_c_325_n 3.67508e-19 $X=0.69 $Y=3.635 $X2=1.335
+ $Y2=2.53
cc_145 N_VDD_c_141_p N_A_27_115#_c_325_n 0.00610567f $X=1.465 $Y=4.287 $X2=1.335
+ $Y2=2.53
cc_146 N_VDD_c_146_p N_A_27_115#_c_325_n 0.0035715f $X=1.55 $Y=2.955 $X2=1.335
+ $Y2=2.53
cc_147 N_VDD_c_133_p N_A_27_115#_c_325_n 0.00470215f $X=3.74 $Y=4.25 $X2=1.335
+ $Y2=2.53
cc_148 N_VDD_M1005_b N_A_27_115#_c_264_n 0.00647677f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.455
cc_149 N_VDD_c_146_p N_A_27_115#_c_264_n 0.00364479f $X=1.55 $Y=2.955 $X2=1.69
+ $Y2=2.455
cc_150 N_VDD_M1005_b N_A_27_115#_c_265_n 0.0113915f $X=-0.045 $Y=2.425 $X2=1.41
+ $Y2=2.455
cc_151 N_VDD_M1005_b N_A_27_115#_c_333_n 0.0137901f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.53
cc_152 N_VDD_c_146_p N_A_27_115#_c_333_n 0.00337744f $X=1.55 $Y=2.955 $X2=1.765
+ $Y2=2.53
cc_153 N_VDD_c_153_p N_A_27_115#_c_333_n 0.00606474f $X=2.325 $Y=4.287 $X2=1.765
+ $Y2=2.53
cc_154 N_VDD_c_133_p N_A_27_115#_c_333_n 0.00468827f $X=3.74 $Y=4.25 $X2=1.765
+ $Y2=2.53
cc_155 N_VDD_M1005_b N_A_27_115#_c_271_n 0.00596183f $X=-0.045 $Y=2.425 $X2=2.12
+ $Y2=2.455
cc_156 N_VDD_M1005_b N_A_27_115#_c_338_n 0.0137901f $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.53
cc_157 N_VDD_c_153_p N_A_27_115#_c_338_n 0.00606474f $X=2.325 $Y=4.287 $X2=2.195
+ $Y2=2.53
cc_158 N_VDD_c_158_p N_A_27_115#_c_338_n 0.00337744f $X=2.41 $Y=2.955 $X2=2.195
+ $Y2=2.53
cc_159 N_VDD_c_133_p N_A_27_115#_c_338_n 0.00468827f $X=3.74 $Y=4.25 $X2=2.195
+ $Y2=2.53
cc_160 N_VDD_M1005_b N_A_27_115#_c_278_n 0.00647677f $X=-0.045 $Y=2.425 $X2=2.55
+ $Y2=2.455
cc_161 N_VDD_c_158_p N_A_27_115#_c_278_n 0.00364479f $X=2.41 $Y=2.955 $X2=2.55
+ $Y2=2.455
cc_162 N_VDD_M1005_b N_A_27_115#_c_344_n 0.0137901f $X=-0.045 $Y=2.425 $X2=2.625
+ $Y2=2.53
cc_163 N_VDD_c_158_p N_A_27_115#_c_344_n 0.00337744f $X=2.41 $Y=2.955 $X2=2.625
+ $Y2=2.53
cc_164 N_VDD_c_164_p N_A_27_115#_c_344_n 0.00606474f $X=3.185 $Y=4.287 $X2=2.625
+ $Y2=2.53
cc_165 N_VDD_c_133_p N_A_27_115#_c_344_n 0.00468827f $X=3.74 $Y=4.25 $X2=2.625
+ $Y2=2.53
cc_166 N_VDD_M1005_b N_A_27_115#_c_285_n 0.00596183f $X=-0.045 $Y=2.425 $X2=2.98
+ $Y2=2.455
cc_167 N_VDD_M1005_b N_A_27_115#_c_349_n 0.0137901f $X=-0.045 $Y=2.425 $X2=3.055
+ $Y2=2.53
cc_168 N_VDD_c_164_p N_A_27_115#_c_349_n 0.00606474f $X=3.185 $Y=4.287 $X2=3.055
+ $Y2=2.53
cc_169 N_VDD_c_169_p N_A_27_115#_c_349_n 0.00337744f $X=3.27 $Y=2.955 $X2=3.055
+ $Y2=2.53
cc_170 N_VDD_c_133_p N_A_27_115#_c_349_n 0.00468827f $X=3.74 $Y=4.25 $X2=3.055
+ $Y2=2.53
cc_171 N_VDD_M1005_b N_A_27_115#_c_292_n 0.00647677f $X=-0.045 $Y=2.425 $X2=3.41
+ $Y2=2.455
cc_172 N_VDD_c_169_p N_A_27_115#_c_292_n 0.00364479f $X=3.27 $Y=2.955 $X2=3.41
+ $Y2=2.455
cc_173 N_VDD_M1005_b N_A_27_115#_c_355_n 0.0137901f $X=-0.045 $Y=2.425 $X2=3.485
+ $Y2=2.53
cc_174 N_VDD_c_169_p N_A_27_115#_c_355_n 0.00337744f $X=3.27 $Y=2.955 $X2=3.485
+ $Y2=2.53
cc_175 N_VDD_c_175_p N_A_27_115#_c_355_n 0.00606474f $X=4.045 $Y=4.287 $X2=3.485
+ $Y2=2.53
cc_176 N_VDD_c_133_p N_A_27_115#_c_355_n 0.00468827f $X=3.74 $Y=4.25 $X2=3.485
+ $Y2=2.53
cc_177 N_VDD_M1005_b N_A_27_115#_c_298_n 0.0134369f $X=-0.045 $Y=2.425 $X2=3.84
+ $Y2=2.455
cc_178 N_VDD_M1005_b N_A_27_115#_c_360_n 0.0166569f $X=-0.045 $Y=2.425 $X2=3.915
+ $Y2=2.53
cc_179 N_VDD_c_175_p N_A_27_115#_c_360_n 0.00606474f $X=4.045 $Y=4.287 $X2=3.915
+ $Y2=2.53
cc_180 N_VDD_c_180_p N_A_27_115#_c_360_n 0.00636672f $X=4.13 $Y=2.955 $X2=3.915
+ $Y2=2.53
cc_181 N_VDD_c_133_p N_A_27_115#_c_360_n 0.00468827f $X=3.74 $Y=4.25 $X2=3.915
+ $Y2=2.53
cc_182 N_VDD_M1005_b N_A_27_115#_c_304_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=1.765 $Y2=2.455
cc_183 N_VDD_M1005_b N_A_27_115#_c_306_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=2.195 $Y2=2.455
cc_184 N_VDD_M1005_b N_A_27_115#_c_308_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=2.625 $Y2=2.455
cc_185 N_VDD_M1005_b N_A_27_115#_c_310_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=3.055 $Y2=2.455
cc_186 N_VDD_M1005_b N_A_27_115#_c_312_n 0.00167153f $X=-0.045 $Y=2.425
+ $X2=3.485 $Y2=2.455
cc_187 N_VDD_M1005_b N_A_27_115#_c_316_n 0.00996008f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=2.955
cc_188 N_VDD_c_131_p N_A_27_115#_c_316_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=2.955
cc_189 N_VDD_c_133_p N_A_27_115#_c_316_n 0.00476261f $X=3.74 $Y=4.25 $X2=0.26
+ $Y2=2.955
cc_190 N_VDD_M1005_b N_Y_c_537_n 0.00290209f $X=-0.045 $Y=2.425 $X2=1.12
+ $Y2=2.48
cc_191 N_VDD_c_141_p N_Y_c_537_n 0.00734006f $X=1.465 $Y=4.287 $X2=1.12 $Y2=2.48
cc_192 N_VDD_c_133_p N_Y_c_537_n 0.00475776f $X=3.74 $Y=4.25 $X2=1.12 $Y2=2.48
cc_193 N_VDD_M1005_b N_Y_c_540_n 0.00337919f $X=-0.045 $Y=2.425 $X2=1.98
+ $Y2=2.48
cc_194 N_VDD_c_153_p N_Y_c_540_n 0.00754406f $X=2.325 $Y=4.287 $X2=1.98 $Y2=2.48
cc_195 N_VDD_c_133_p N_Y_c_540_n 0.00475776f $X=3.74 $Y=4.25 $X2=1.98 $Y2=2.48
cc_196 N_VDD_M1005_b N_Y_c_543_n 0.00337919f $X=-0.045 $Y=2.425 $X2=2.84
+ $Y2=2.48
cc_197 N_VDD_c_164_p N_Y_c_543_n 0.00746708f $X=3.185 $Y=4.287 $X2=2.84 $Y2=2.48
cc_198 N_VDD_c_133_p N_Y_c_543_n 0.00475776f $X=3.74 $Y=4.25 $X2=2.84 $Y2=2.48
cc_199 N_VDD_M1005_b N_Y_c_546_n 0.00337919f $X=-0.045 $Y=2.425 $X2=3.7 $Y2=2.48
cc_200 N_VDD_c_175_p N_Y_c_546_n 0.00734006f $X=4.045 $Y=4.287 $X2=3.7 $Y2=2.48
cc_201 N_VDD_c_133_p N_Y_c_546_n 0.00475776f $X=3.74 $Y=4.25 $X2=3.7 $Y2=2.48
cc_202 N_VDD_M1005_b N_Y_c_506_n 0.00409378f $X=-0.045 $Y=2.425 $X2=1.12
+ $Y2=2.365
cc_203 N_VDD_M1005_b N_Y_c_550_n 0.00520877f $X=-0.045 $Y=2.425 $X2=1.835
+ $Y2=2.48
cc_204 N_VDD_c_146_p N_Y_c_550_n 0.0090257f $X=1.55 $Y=2.955 $X2=1.835 $Y2=2.48
cc_205 N_VDD_M1005_b N_Y_c_552_n 0.00520877f $X=-0.045 $Y=2.425 $X2=2.695
+ $Y2=2.48
cc_206 N_VDD_c_158_p N_Y_c_552_n 0.0090257f $X=2.41 $Y=2.955 $X2=2.695 $Y2=2.48
cc_207 N_VDD_M1005_b N_Y_c_521_n 0.00409378f $X=-0.045 $Y=2.425 $X2=2.125
+ $Y2=2.48
cc_208 N_VDD_M1005_b N_Y_c_555_n 0.00520877f $X=-0.045 $Y=2.425 $X2=3.555
+ $Y2=2.48
cc_209 N_VDD_c_169_p N_Y_c_555_n 0.0090257f $X=3.27 $Y=2.955 $X2=3.555 $Y2=2.48
cc_210 N_VDD_M1005_b N_Y_c_531_n 0.00409378f $X=-0.045 $Y=2.425 $X2=2.985
+ $Y2=2.48
cc_211 N_VDD_M1005_b N_Y_c_536_n 0.00409378f $X=-0.045 $Y=2.425 $X2=3.7
+ $Y2=2.365
cc_212 A N_A_27_115#_M1005_s 0.00410657f $X=0.635 $Y=2.85 $X2=0.135 $Y2=2.605
cc_213 N_A_M1007_g N_A_27_115#_M1000_g 0.0342527f $X=0.475 $Y=0.835 $X2=0.905
+ $Y2=0.835
cc_214 A N_A_27_115#_c_321_n 0.00419145f $X=0.635 $Y=2.85 $X2=0.905 $Y2=2.53
cc_215 N_A_M1007_g N_A_27_115#_c_256_n 0.00260138f $X=0.475 $Y=0.835 $X2=1.18
+ $Y2=2.38
cc_216 N_A_M1005_g N_A_27_115#_c_256_n 0.00209773f $X=0.475 $Y=3.235 $X2=1.18
+ $Y2=2.38
cc_217 N_A_c_217_n N_A_27_115#_c_256_n 0.0139096f $X=0.635 $Y=2 $X2=1.18
+ $Y2=2.38
cc_218 N_A_c_218_n N_A_27_115#_c_256_n 0.00361737f $X=0.635 $Y=2 $X2=1.18
+ $Y2=2.38
cc_219 N_A_M1005_g N_A_27_115#_c_265_n 0.0485392f $X=0.475 $Y=3.235 $X2=1.41
+ $Y2=2.455
cc_220 N_A_c_218_n N_A_27_115#_c_265_n 0.00477416f $X=0.635 $Y=2 $X2=1.41
+ $Y2=2.455
cc_221 N_A_M1007_g N_A_27_115#_c_313_n 0.0124465f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.755
cc_222 N_A_M1007_g N_A_27_115#_c_316_n 0.0330322f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=2.955
cc_223 N_A_c_218_n N_A_27_115#_c_316_n 0.0548951f $X=0.635 $Y=2 $X2=0.26
+ $Y2=2.955
cc_224 A N_A_27_115#_c_316_n 0.0155137f $X=0.635 $Y=2.85 $X2=0.26 $Y2=2.955
cc_225 N_A_M1007_g N_A_27_115#_c_317_n 0.0207696f $X=0.475 $Y=0.835 $X2=0.88
+ $Y2=1.455
cc_226 N_A_c_217_n N_A_27_115#_c_317_n 0.00273049f $X=0.635 $Y=2 $X2=0.88
+ $Y2=1.455
cc_227 N_A_c_218_n N_A_27_115#_c_317_n 0.00886797f $X=0.635 $Y=2 $X2=0.88
+ $Y2=1.455
cc_228 N_A_M1007_g N_A_27_115#_c_320_n 6.59135e-19 $X=0.475 $Y=0.835 $X2=0.965
+ $Y2=1.455
cc_229 N_A_c_218_n N_Y_c_537_n 0.0135622f $X=0.635 $Y=2 $X2=1.12 $Y2=2.48
cc_230 A N_Y_c_537_n 0.00731851f $X=0.635 $Y=2.85 $X2=1.12 $Y2=2.48
cc_231 N_A_M1007_g N_Y_c_502_n 8.01483e-19 $X=0.475 $Y=0.835 $X2=1.12 $Y2=1.115
cc_232 N_A_c_218_n N_Y_c_506_n 0.00677552f $X=0.635 $Y=2 $X2=1.12 $Y2=2.365
cc_233 N_A_M1007_g Y 0.00310306f $X=0.475 $Y=0.835 $X2=1.055 $Y2=1.79
cc_234 N_A_c_217_n Y 0.00441844f $X=0.635 $Y=2 $X2=1.055 $Y2=1.79
cc_235 N_A_c_218_n Y 0.0200396f $X=0.635 $Y=2 $X2=1.055 $Y2=1.79
cc_236 N_A_27_115#_M1000_g N_Y_c_484_n 0.00182852f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_237 N_A_27_115#_M1001_g N_Y_c_484_n 0.00182852f $X=1.335 $Y=0.835 $X2=1.12
+ $Y2=0.755
cc_238 N_A_27_115#_c_263_n N_Y_c_484_n 0.00296072f $X=1.41 $Y=1.365 $X2=1.12
+ $Y2=0.755
cc_239 N_A_27_115#_c_320_n N_Y_c_484_n 7.29965e-19 $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=0.755
cc_240 N_A_27_115#_c_321_n N_Y_c_537_n 0.00138273f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_241 N_A_27_115#_c_325_n N_Y_c_537_n 0.00233646f $X=1.335 $Y=2.53 $X2=1.12
+ $Y2=2.48
cc_242 N_A_27_115#_c_265_n N_Y_c_537_n 0.0126676f $X=1.41 $Y=2.455 $X2=1.12
+ $Y2=2.48
cc_243 N_A_27_115#_M1008_g N_Y_c_488_n 0.00182852f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=0.755
cc_244 N_A_27_115#_c_270_n N_Y_c_488_n 0.00274041f $X=2.12 $Y=1.365 $X2=1.98
+ $Y2=0.755
cc_245 N_A_27_115#_M1010_g N_Y_c_488_n 0.00182852f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=0.755
cc_246 N_A_27_115#_c_333_n N_Y_c_540_n 0.00233646f $X=1.765 $Y=2.53 $X2=1.98
+ $Y2=2.48
cc_247 N_A_27_115#_c_271_n N_Y_c_540_n 0.0138847f $X=2.12 $Y=2.455 $X2=1.98
+ $Y2=2.48
cc_248 N_A_27_115#_c_338_n N_Y_c_540_n 0.00233646f $X=2.195 $Y=2.53 $X2=1.98
+ $Y2=2.48
cc_249 N_A_27_115#_M1012_g N_Y_c_493_n 0.00182852f $X=2.625 $Y=0.835 $X2=2.84
+ $Y2=0.755
cc_250 N_A_27_115#_c_284_n N_Y_c_493_n 0.00274041f $X=2.98 $Y=1.365 $X2=2.84
+ $Y2=0.755
cc_251 N_A_27_115#_M1013_g N_Y_c_493_n 0.00182852f $X=3.055 $Y=0.835 $X2=2.84
+ $Y2=0.755
cc_252 N_A_27_115#_c_344_n N_Y_c_543_n 0.00233646f $X=2.625 $Y=2.53 $X2=2.84
+ $Y2=2.48
cc_253 N_A_27_115#_c_285_n N_Y_c_543_n 0.0138847f $X=2.98 $Y=2.455 $X2=2.84
+ $Y2=2.48
cc_254 N_A_27_115#_c_349_n N_Y_c_543_n 0.00233646f $X=3.055 $Y=2.53 $X2=2.84
+ $Y2=2.48
cc_255 N_A_27_115#_M1014_g N_Y_c_498_n 0.00182852f $X=3.485 $Y=0.835 $X2=3.7
+ $Y2=0.755
cc_256 N_A_27_115#_c_297_n N_Y_c_498_n 0.00274041f $X=3.84 $Y=1.365 $X2=3.7
+ $Y2=0.755
cc_257 N_A_27_115#_M1017_g N_Y_c_498_n 0.00182852f $X=3.915 $Y=0.835 $X2=3.7
+ $Y2=0.755
cc_258 N_A_27_115#_c_355_n N_Y_c_546_n 0.00233646f $X=3.485 $Y=2.53 $X2=3.7
+ $Y2=2.48
cc_259 N_A_27_115#_c_298_n N_Y_c_546_n 0.013404f $X=3.84 $Y=2.455 $X2=3.7
+ $Y2=2.48
cc_260 N_A_27_115#_c_360_n N_Y_c_546_n 0.00233646f $X=3.915 $Y=2.53 $X2=3.7
+ $Y2=2.48
cc_261 N_A_27_115#_M1000_g N_Y_c_502_n 0.00480694f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=1.115
cc_262 N_A_27_115#_M1001_g N_Y_c_502_n 0.00201073f $X=1.335 $Y=0.835 $X2=1.12
+ $Y2=1.115
cc_263 N_A_27_115#_c_320_n N_Y_c_502_n 0.00278861f $X=0.965 $Y=1.455 $X2=1.12
+ $Y2=1.115
cc_264 N_A_27_115#_c_321_n N_Y_c_506_n 0.00120715f $X=0.905 $Y=2.53 $X2=1.12
+ $Y2=2.365
cc_265 N_A_27_115#_c_256_n N_Y_c_506_n 0.00215118f $X=1.18 $Y=2.38 $X2=1.12
+ $Y2=2.365
cc_266 N_A_27_115#_c_325_n N_Y_c_506_n 0.00113627f $X=1.335 $Y=2.53 $X2=1.12
+ $Y2=2.365
cc_267 N_A_27_115#_c_265_n N_Y_c_506_n 0.00372325f $X=1.41 $Y=2.455 $X2=1.12
+ $Y2=2.365
cc_268 N_A_27_115#_M1000_g Y 0.00251111f $X=0.905 $Y=0.835 $X2=1.055 $Y2=1.79
cc_269 N_A_27_115#_c_256_n Y 0.0314621f $X=1.18 $Y=2.38 $X2=1.055 $Y2=1.79
cc_270 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=0.835 $X2=1.055 $Y2=1.79
cc_271 N_A_27_115#_c_263_n Y 0.0166018f $X=1.41 $Y=1.365 $X2=1.055 $Y2=1.79
cc_272 N_A_27_115#_c_317_n Y 8.73078e-19 $X=0.88 $Y=1.455 $X2=1.055 $Y2=1.79
cc_273 N_A_27_115#_c_320_n Y 0.0121742f $X=0.965 $Y=1.455 $X2=1.055 $Y2=1.79
cc_274 N_A_27_115#_M1001_g N_Y_c_508_n 0.00908832f $X=1.335 $Y=0.835 $X2=1.835
+ $Y2=1
cc_275 N_A_27_115#_c_261_n N_Y_c_508_n 0.00213861f $X=1.69 $Y=1.365 $X2=1.835
+ $Y2=1
cc_276 N_A_27_115#_M1008_g N_Y_c_508_n 0.00873177f $X=1.765 $Y=0.835 $X2=1.835
+ $Y2=1
cc_277 N_A_27_115#_c_325_n N_Y_c_550_n 0.00639369f $X=1.335 $Y=2.53 $X2=1.835
+ $Y2=2.48
cc_278 N_A_27_115#_c_264_n N_Y_c_550_n 0.0125005f $X=1.69 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_279 N_A_27_115#_c_265_n N_Y_c_550_n 0.00627763f $X=1.41 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_280 N_A_27_115#_c_333_n N_Y_c_550_n 0.00639369f $X=1.765 $Y=2.53 $X2=1.835
+ $Y2=2.48
cc_281 N_A_27_115#_c_304_n N_Y_c_550_n 0.00580646f $X=1.765 $Y=2.455 $X2=1.835
+ $Y2=2.48
cc_282 N_A_27_115#_c_263_n N_Y_c_512_n 0.013329f $X=1.41 $Y=1.365 $X2=1.98
+ $Y2=2.365
cc_283 N_A_27_115#_M1008_g N_Y_c_512_n 0.00251111f $X=1.765 $Y=0.835 $X2=1.98
+ $Y2=2.365
cc_284 N_A_27_115#_c_270_n N_Y_c_512_n 0.0178059f $X=2.12 $Y=1.365 $X2=1.98
+ $Y2=2.365
cc_285 N_A_27_115#_M1010_g N_Y_c_512_n 0.00251111f $X=2.195 $Y=0.835 $X2=1.98
+ $Y2=2.365
cc_286 N_A_27_115#_c_283_n N_Y_c_512_n 0.0137936f $X=2.625 $Y=2.38 $X2=1.98
+ $Y2=2.365
cc_287 N_A_27_115#_M1010_g N_Y_c_513_n 0.00873177f $X=2.195 $Y=0.835 $X2=2.695
+ $Y2=1
cc_288 N_A_27_115#_c_276_n N_Y_c_513_n 0.00213861f $X=2.55 $Y=1.365 $X2=2.695
+ $Y2=1
cc_289 N_A_27_115#_M1012_g N_Y_c_513_n 0.00938169f $X=2.625 $Y=0.835 $X2=2.695
+ $Y2=1
cc_290 N_A_27_115#_M1008_g N_Y_c_517_n 0.00198614f $X=1.765 $Y=0.835 $X2=2.125
+ $Y2=1
cc_291 N_A_27_115#_M1010_g N_Y_c_517_n 0.00198614f $X=2.195 $Y=0.835 $X2=2.125
+ $Y2=1
cc_292 N_A_27_115#_c_338_n N_Y_c_552_n 0.00639369f $X=2.195 $Y=2.53 $X2=2.695
+ $Y2=2.48
cc_293 N_A_27_115#_c_278_n N_Y_c_552_n 0.0130313f $X=2.55 $Y=2.455 $X2=2.695
+ $Y2=2.48
cc_294 N_A_27_115#_c_344_n N_Y_c_552_n 0.00639369f $X=2.625 $Y=2.53 $X2=2.695
+ $Y2=2.48
cc_295 N_A_27_115#_c_306_n N_Y_c_552_n 0.00580646f $X=2.195 $Y=2.455 $X2=2.695
+ $Y2=2.48
cc_296 N_A_27_115#_c_308_n N_Y_c_552_n 0.00666531f $X=2.625 $Y=2.455 $X2=2.695
+ $Y2=2.48
cc_297 N_A_27_115#_c_333_n N_Y_c_521_n 0.00113627f $X=1.765 $Y=2.53 $X2=2.125
+ $Y2=2.48
cc_298 N_A_27_115#_c_271_n N_Y_c_521_n 0.00364679f $X=2.12 $Y=2.455 $X2=2.125
+ $Y2=2.48
cc_299 N_A_27_115#_c_338_n N_Y_c_521_n 0.00113627f $X=2.195 $Y=2.53 $X2=2.125
+ $Y2=2.48
cc_300 N_A_27_115#_c_304_n N_Y_c_521_n 6.99501e-19 $X=1.765 $Y=2.455 $X2=2.125
+ $Y2=2.48
cc_301 N_A_27_115#_c_306_n N_Y_c_521_n 6.99501e-19 $X=2.195 $Y=2.455 $X2=2.125
+ $Y2=2.48
cc_302 N_A_27_115#_M1012_g N_Y_c_522_n 0.00251111f $X=2.625 $Y=0.835 $X2=2.84
+ $Y2=2.365
cc_303 N_A_27_115#_c_283_n N_Y_c_522_n 0.017762f $X=2.625 $Y=2.38 $X2=2.84
+ $Y2=2.365
cc_304 N_A_27_115#_c_284_n N_Y_c_522_n 0.0178059f $X=2.98 $Y=1.365 $X2=2.84
+ $Y2=2.365
cc_305 N_A_27_115#_M1013_g N_Y_c_522_n 0.00251111f $X=3.055 $Y=0.835 $X2=2.84
+ $Y2=2.365
cc_306 N_A_27_115#_M1013_g N_Y_c_523_n 0.00873177f $X=3.055 $Y=0.835 $X2=3.555
+ $Y2=1
cc_307 N_A_27_115#_c_290_n N_Y_c_523_n 0.00213861f $X=3.41 $Y=1.365 $X2=3.555
+ $Y2=1
cc_308 N_A_27_115#_M1014_g N_Y_c_523_n 0.00873177f $X=3.485 $Y=0.835 $X2=3.555
+ $Y2=1
cc_309 N_A_27_115#_M1012_g N_Y_c_527_n 0.00201073f $X=2.625 $Y=0.835 $X2=2.985
+ $Y2=1
cc_310 N_A_27_115#_M1013_g N_Y_c_527_n 0.00198614f $X=3.055 $Y=0.835 $X2=2.985
+ $Y2=1
cc_311 N_A_27_115#_c_349_n N_Y_c_555_n 0.00639369f $X=3.055 $Y=2.53 $X2=3.555
+ $Y2=2.48
cc_312 N_A_27_115#_c_292_n N_Y_c_555_n 0.0125005f $X=3.41 $Y=2.455 $X2=3.555
+ $Y2=2.48
cc_313 N_A_27_115#_c_355_n N_Y_c_555_n 0.00639369f $X=3.485 $Y=2.53 $X2=3.555
+ $Y2=2.48
cc_314 N_A_27_115#_c_310_n N_Y_c_555_n 0.00580646f $X=3.055 $Y=2.455 $X2=3.555
+ $Y2=2.48
cc_315 N_A_27_115#_c_312_n N_Y_c_555_n 0.00580646f $X=3.485 $Y=2.455 $X2=3.555
+ $Y2=2.48
cc_316 N_A_27_115#_c_283_n N_Y_c_531_n 8.30534e-19 $X=2.625 $Y=2.38 $X2=2.985
+ $Y2=2.48
cc_317 N_A_27_115#_c_344_n N_Y_c_531_n 0.00113627f $X=2.625 $Y=2.53 $X2=2.985
+ $Y2=2.48
cc_318 N_A_27_115#_c_285_n N_Y_c_531_n 0.00364679f $X=2.98 $Y=2.455 $X2=2.985
+ $Y2=2.48
cc_319 N_A_27_115#_c_349_n N_Y_c_531_n 0.00113627f $X=3.055 $Y=2.53 $X2=2.985
+ $Y2=2.48
cc_320 N_A_27_115#_c_308_n N_Y_c_531_n 6.59375e-19 $X=2.625 $Y=2.455 $X2=2.985
+ $Y2=2.48
cc_321 N_A_27_115#_c_310_n N_Y_c_531_n 6.99501e-19 $X=3.055 $Y=2.455 $X2=2.985
+ $Y2=2.48
cc_322 N_A_27_115#_M1014_g N_Y_c_532_n 0.00198614f $X=3.485 $Y=0.835 $X2=3.7
+ $Y2=1.115
cc_323 N_A_27_115#_M1017_g N_Y_c_532_n 0.00878256f $X=3.915 $Y=0.835 $X2=3.7
+ $Y2=1.115
cc_324 N_A_27_115#_M1014_g N_Y_c_536_n 0.00251111f $X=3.485 $Y=0.835 $X2=3.7
+ $Y2=2.365
cc_325 N_A_27_115#_c_355_n N_Y_c_536_n 0.00113627f $X=3.485 $Y=2.53 $X2=3.7
+ $Y2=2.365
cc_326 N_A_27_115#_c_297_n N_Y_c_536_n 0.0170354f $X=3.84 $Y=1.365 $X2=3.7
+ $Y2=2.365
cc_327 N_A_27_115#_c_298_n N_Y_c_536_n 0.00966211f $X=3.84 $Y=2.455 $X2=3.7
+ $Y2=2.365
cc_328 N_A_27_115#_M1017_g N_Y_c_536_n 0.00251111f $X=3.915 $Y=0.835 $X2=3.7
+ $Y2=2.365
cc_329 N_A_27_115#_c_360_n N_Y_c_536_n 0.0031083f $X=3.915 $Y=2.53 $X2=3.7
+ $Y2=2.365
cc_330 N_A_27_115#_c_312_n N_Y_c_536_n 6.99501e-19 $X=3.485 $Y=2.455 $X2=3.7
+ $Y2=2.365
