* File: sky130_osu_sc_15T_hs__addh_l.pxi.spice
* Created: Fri Nov 12 14:26:33 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%GND N_GND_M1006_d N_GND_M1001_d N_GND_M1006_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_25_p N_GND_c_9_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_15T_HS__ADDH_L%GND
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%VDD N_VDD_M1002_d N_VDD_M1003_d N_VDD_M1011_d
+ N_VDD_M1003_b N_VDD_c_97_p N_VDD_c_98_p N_VDD_c_111_p N_VDD_c_119_p
+ N_VDD_c_101_p N_VDD_c_104_p N_VDD_c_106_p VDD N_VDD_c_99_p
+ PM_SKY130_OSU_SC_15T_HS__ADDH_L%VDD
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%CON N_CON_M1004_d N_CON_M1002_s N_CON_M1000_d
+ N_CON_M1006_g N_CON_M1003_g N_CON_c_158_n N_CON_c_159_n N_CON_c_161_n
+ N_CON_c_162_n N_CON_c_179_n N_CON_c_163_n N_CON_c_164_n N_CON_c_165_n
+ N_CON_c_166_n N_CON_c_184_n N_CON_c_167_n N_CON_c_168_n N_CON_c_170_n
+ N_CON_c_172_n CON PM_SKY130_OSU_SC_15T_HS__ADDH_L%CON
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%B N_B_M1007_g N_B_M1010_g N_B_M1004_g
+ N_B_M1013_g N_B_c_290_n N_B_c_292_n N_B_c_293_n N_B_c_295_n N_B_c_296_n
+ N_B_c_297_n B PM_SKY130_OSU_SC_15T_HS__ADDH_L%B
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%A N_A_M1008_g N_A_M1011_g N_A_M1000_g
+ N_A_M1005_g N_A_c_391_n N_A_c_392_n N_A_c_393_n N_A_c_394_n N_A_c_395_n A
+ N_A_c_397_n PM_SKY130_OSU_SC_15T_HS__ADDH_L%A
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%A_208_565# N_A_208_565#_M1008_d
+ N_A_208_565#_M1010_d N_A_208_565#_c_471_n N_A_208_565#_c_472_n
+ N_A_208_565#_M1012_g N_A_208_565#_c_474_n N_A_208_565#_c_475_n
+ N_A_208_565#_M1001_g N_A_208_565#_c_480_n N_A_208_565#_c_482_n
+ N_A_208_565#_M1009_g N_A_208_565#_M1002_g N_A_208_565#_c_486_n
+ N_A_208_565#_c_487_n N_A_208_565#_c_501_n N_A_208_565#_c_504_n
+ N_A_208_565#_c_507_n N_A_208_565#_c_488_n N_A_208_565#_c_491_n
+ N_A_208_565#_c_492_n PM_SKY130_OSU_SC_15T_HS__ADDH_L%A_208_565#
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%S N_S_M1006_s N_S_M1003_s N_S_c_586_n
+ N_S_c_593_n S N_S_c_591_n N_S_c_598_n PM_SKY130_OSU_SC_15T_HS__ADDH_L%S
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%CO N_CO_M1001_s N_CO_M1012_d N_CO_c_617_n
+ N_CO_c_625_n N_CO_c_620_n N_CO_c_622_n N_CO_c_623_n CO
+ PM_SKY130_OSU_SC_15T_HS__ADDH_L%CO
x_PM_SKY130_OSU_SC_15T_HS__ADDH_L%A_570_115# N_A_570_115#_M1009_d
+ N_A_570_115#_M1005_d N_A_570_115#_c_675_n N_A_570_115#_c_670_n
+ N_A_570_115#_c_672_n PM_SKY130_OSU_SC_15T_HS__ADDH_L%A_570_115#
cc_1 N_GND_M1006_b N_CON_M1006_g 0.0359014f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_CON_M1006_g 0.00606474f $X=0.665 $Y=0.152 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_CON_M1006_g 0.00882091f $X=0.75 $Y=0.74 $X2=0.475 $Y2=0.85
cc_4 N_GND_c_4_p N_CON_M1006_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.475 $Y2=0.85
cc_5 N_GND_M1006_b N_CON_M1003_g 0.060974f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.195
cc_6 N_GND_M1006_b N_CON_c_158_n 0.0413643f $X=-0.045 $Y=0 $X2=0.35 $Y2=1.59
cc_7 N_GND_M1006_b N_CON_c_159_n 0.00877401f $X=-0.045 $Y=0 $X2=0.635 $Y2=1.59
cc_8 N_GND_c_3_p N_CON_c_159_n 0.00248867f $X=0.75 $Y=0.74 $X2=0.635 $Y2=1.59
cc_9 N_GND_c_9_p N_CON_c_161_n 0.00470352f $X=2.56 $Y=0.74 $X2=2.62 $Y2=1.675
cc_10 N_GND_M1006_b N_CON_c_162_n 0.0155029f $X=-0.045 $Y=0 $X2=2.62 $Y2=2.605
cc_11 N_GND_M1006_b N_CON_c_163_n 0.0100275f $X=-0.045 $Y=0 $X2=3.335 $Y2=1.59
cc_12 N_GND_M1006_b N_CON_c_164_n 0.0112921f $X=-0.045 $Y=0 $X2=3.755 $Y2=2.69
cc_13 N_GND_M1006_b N_CON_c_165_n 0.00433753f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.505
cc_14 N_GND_M1006_b N_CON_c_166_n 0.00195909f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.065
cc_15 N_GND_M1006_b N_CON_c_167_n 2.79926e-19 $X=-0.045 $Y=0 $X2=2.62 $Y2=2.69
cc_16 N_GND_M1006_b N_CON_c_168_n 0.0196394f $X=-0.045 $Y=0 $X2=2.475 $Y2=1.59
cc_17 N_GND_c_3_p N_CON_c_168_n 0.00166299f $X=0.75 $Y=0.74 $X2=2.475 $Y2=1.59
cc_18 N_GND_M1006_b N_CON_c_170_n 0.0133709f $X=-0.045 $Y=0 $X2=0.78 $Y2=1.59
cc_19 N_GND_c_3_p N_CON_c_170_n 0.00391282f $X=0.75 $Y=0.74 $X2=0.78 $Y2=1.59
cc_20 N_GND_M1006_b N_CON_c_172_n 0.00474051f $X=-0.045 $Y=0 $X2=2.62 $Y2=1.59
cc_21 N_GND_c_9_p N_CON_c_172_n 0.00612077f $X=2.56 $Y=0.74 $X2=2.62 $Y2=1.59
cc_22 N_GND_M1006_b CON 0.00668459f $X=-0.045 $Y=0 $X2=3.42 $Y2=1.59
cc_23 N_GND_M1006_b N_B_M1007_g 0.0292341f $X=-0.045 $Y=0 $X2=0.965 $Y2=0.995
cc_24 N_GND_c_3_p N_B_M1007_g 0.00318344f $X=0.75 $Y=0.74 $X2=0.965 $Y2=0.995
cc_25 N_GND_c_25_p N_B_M1007_g 0.00606474f $X=2.475 $Y=0.152 $X2=0.965 $Y2=0.995
cc_26 N_GND_c_4_p N_B_M1007_g 0.00468827f $X=3.74 $Y=0.19 $X2=0.965 $Y2=0.995
cc_27 N_GND_M1006_b N_B_M1010_g 0.0282323f $X=-0.045 $Y=0 $X2=0.965 $Y2=3.825
cc_28 N_GND_M1006_b N_B_M1004_g 0.0334167f $X=-0.045 $Y=0 $X2=3.205 $Y2=0.995
cc_29 N_GND_c_4_p N_B_M1004_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.205 $Y2=0.995
cc_30 N_GND_M1006_b N_B_M1013_g 0.0272084f $X=-0.045 $Y=0 $X2=3.265 $Y2=3.825
cc_31 N_GND_M1006_b N_B_c_290_n 0.0278498f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.96
cc_32 N_GND_c_3_p N_B_c_290_n 0.00118315f $X=0.75 $Y=0.74 $X2=0.905 $Y2=1.96
cc_33 N_GND_M1006_b N_B_c_292_n 0.0299556f $X=-0.045 $Y=0 $X2=3.205 $Y2=1.96
cc_34 N_GND_M1006_b N_B_c_293_n 0.00405307f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.96
cc_35 N_GND_c_3_p N_B_c_293_n 0.00111247f $X=0.75 $Y=0.74 $X2=0.905 $Y2=1.96
cc_36 N_GND_M1006_b N_B_c_295_n 0.00365598f $X=-0.045 $Y=0 $X2=3.205 $Y2=1.96
cc_37 N_GND_M1006_b N_B_c_296_n 0.00204225f $X=-0.045 $Y=0 $X2=1.05 $Y2=1.96
cc_38 N_GND_M1006_b N_B_c_297_n 0.0175444f $X=-0.045 $Y=0 $X2=3.06 $Y2=1.96
cc_39 N_GND_M1006_b B 0.00164195f $X=-0.045 $Y=0 $X2=3.21 $Y2=1.96
cc_40 N_GND_M1006_b N_A_M1008_g 0.050508f $X=-0.045 $Y=0 $X2=1.325 $Y2=0.995
cc_41 N_GND_c_25_p N_A_M1008_g 0.00606474f $X=2.475 $Y=0.152 $X2=1.325 $Y2=0.995
cc_42 N_GND_c_4_p N_A_M1008_g 0.00468827f $X=3.74 $Y=0.19 $X2=1.325 $Y2=0.995
cc_43 N_GND_M1006_b N_A_M1011_g 0.00835457f $X=-0.045 $Y=0 $X2=1.395 $Y2=3.825
cc_44 N_GND_M1006_b N_A_M1000_g 0.0108664f $X=-0.045 $Y=0 $X2=3.625 $Y2=3.825
cc_45 N_GND_M1006_b N_A_M1005_g 0.0755267f $X=-0.045 $Y=0 $X2=3.635 $Y2=0.995
cc_46 N_GND_c_4_p N_A_M1005_g 0.00468827f $X=3.74 $Y=0.19 $X2=3.635 $Y2=0.995
cc_47 N_GND_M1006_b N_A_c_391_n 0.0253796f $X=-0.045 $Y=0 $X2=1.385 $Y2=2.33
cc_48 N_GND_M1006_b N_A_c_392_n 0.034256f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.33
cc_49 N_GND_M1006_b N_A_c_393_n 9.49347e-19 $X=-0.045 $Y=0 $X2=1.385 $Y2=2.33
cc_50 N_GND_M1006_b N_A_c_394_n 0.00995238f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.33
cc_51 N_GND_M1006_b N_A_c_395_n 0.00430309f $X=-0.045 $Y=0 $X2=1.53 $Y2=2.33
cc_52 N_GND_M1006_b A 0.00380188f $X=-0.045 $Y=0 $X2=3.685 $Y2=2.33
cc_53 N_GND_M1006_b N_A_c_397_n 0.0115252f $X=-0.045 $Y=0 $X2=3.54 $Y2=2.33
cc_54 N_GND_M1006_b N_A_208_565#_c_471_n 0.0381678f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=1.86
cc_55 N_GND_M1006_b N_A_208_565#_c_472_n 0.0270254f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=2.335
cc_56 N_GND_M1006_b N_A_208_565#_M1012_g 0.00928694f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=4.195
cc_57 N_GND_M1006_b N_A_208_565#_c_474_n 0.0168875f $X=-0.045 $Y=0 $X2=2.21
+ $Y2=1.565
cc_58 N_GND_M1006_b N_A_208_565#_c_475_n 0.0616052f $X=-0.045 $Y=0 $X2=2.76
+ $Y2=2.41
cc_59 N_GND_M1006_b N_A_208_565#_M1001_g 0.0318047f $X=-0.045 $Y=0 $X2=2.285
+ $Y2=0.895
cc_60 N_GND_c_25_p N_A_208_565#_M1001_g 0.00606474f $X=2.475 $Y=0.152 $X2=2.285
+ $Y2=0.895
cc_61 N_GND_c_9_p N_A_208_565#_M1001_g 0.00868712f $X=2.56 $Y=0.74 $X2=2.285
+ $Y2=0.895
cc_62 N_GND_c_4_p N_A_208_565#_M1001_g 0.00468827f $X=3.74 $Y=0.19 $X2=2.285
+ $Y2=0.895
cc_63 N_GND_M1006_b N_A_208_565#_c_480_n 0.0273212f $X=-0.045 $Y=0 $X2=2.7
+ $Y2=1.565
cc_64 N_GND_c_9_p N_A_208_565#_c_480_n 0.00319024f $X=2.56 $Y=0.74 $X2=2.7
+ $Y2=1.565
cc_65 N_GND_M1006_b N_A_208_565#_c_482_n 0.0209741f $X=-0.045 $Y=0 $X2=2.775
+ $Y2=1.49
cc_66 N_GND_c_9_p N_A_208_565#_c_482_n 0.00163921f $X=2.56 $Y=0.74 $X2=2.775
+ $Y2=1.49
cc_67 N_GND_c_4_p N_A_208_565#_c_482_n 0.00468827f $X=3.74 $Y=0.19 $X2=2.775
+ $Y2=1.49
cc_68 N_GND_M1006_b N_A_208_565#_M1002_g 0.00900107f $X=-0.045 $Y=0 $X2=2.835
+ $Y2=3.825
cc_69 N_GND_M1006_b N_A_208_565#_c_486_n 0.00492701f $X=-0.045 $Y=0 $X2=1.885
+ $Y2=2.41
cc_70 N_GND_M1006_b N_A_208_565#_c_487_n 0.00608465f $X=-0.045 $Y=0 $X2=2.285
+ $Y2=1.565
cc_71 N_GND_M1006_b N_A_208_565#_c_488_n 0.00396179f $X=-0.045 $Y=0 $X2=1.54
+ $Y2=0.74
cc_72 N_GND_c_25_p N_A_208_565#_c_488_n 0.00741243f $X=2.475 $Y=0.152 $X2=1.54
+ $Y2=0.74
cc_73 N_GND_c_4_p N_A_208_565#_c_488_n 0.00476261f $X=3.74 $Y=0.19 $X2=1.54
+ $Y2=0.74
cc_74 N_GND_M1006_b N_A_208_565#_c_491_n 0.0137594f $X=-0.045 $Y=0 $X2=1.725
+ $Y2=2.665
cc_75 N_GND_M1006_b N_A_208_565#_c_492_n 0.00684174f $X=-0.045 $Y=0 $X2=1.725
+ $Y2=1.695
cc_76 N_GND_M1006_b N_S_c_586_n 0.00704303f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.825
cc_77 N_GND_c_2_p N_S_c_586_n 0.00736239f $X=0.665 $Y=0.152 $X2=0.26 $Y2=0.825
cc_78 N_GND_c_3_p N_S_c_586_n 0.0165502f $X=0.75 $Y=0.74 $X2=0.26 $Y2=0.825
cc_79 N_GND_c_4_p N_S_c_586_n 0.00476261f $X=3.74 $Y=0.19 $X2=0.26 $Y2=0.825
cc_80 N_GND_M1006_b S 0.063433f $X=-0.045 $Y=0 $X2=0.25 $Y2=2.125
cc_81 N_GND_M1006_b N_S_c_591_n 0.0121294f $X=-0.045 $Y=0 $X2=0.26 $Y2=1.215
cc_82 N_GND_c_3_p N_S_c_591_n 0.00348655f $X=0.75 $Y=0.74 $X2=0.26 $Y2=1.215
cc_83 N_GND_M1006_b N_CO_c_617_n 0.0015547f $X=-0.045 $Y=0 $X2=2.07 $Y2=0.825
cc_84 N_GND_c_25_p N_CO_c_617_n 0.00746729f $X=2.475 $Y=0.152 $X2=2.07 $Y2=0.825
cc_85 N_GND_c_4_p N_CO_c_617_n 0.0047312f $X=3.74 $Y=0.19 $X2=2.07 $Y2=0.825
cc_86 N_GND_M1006_b N_CO_c_620_n 0.00150848f $X=-0.045 $Y=0 $X2=2.175 $Y2=1.215
cc_87 N_GND_c_9_p N_CO_c_620_n 0.00695566f $X=2.56 $Y=0.74 $X2=2.175 $Y2=1.215
cc_88 N_GND_M1006_b N_CO_c_622_n 0.00130468f $X=-0.045 $Y=0 $X2=2.175 $Y2=2.7
cc_89 N_GND_M1006_b N_CO_c_623_n 0.0163213f $X=-0.045 $Y=0 $X2=2.137 $Y2=2.615
cc_90 N_GND_M1006_b CO 0.00219851f $X=-0.045 $Y=0 $X2=2.175 $Y2=2.7
cc_91 N_GND_M1006_b N_A_570_115#_c_670_n 0.0652319f $X=-0.045 $Y=0 $X2=3.765
+ $Y2=0.56
cc_92 N_GND_c_4_p N_A_570_115#_c_670_n 0.024842f $X=3.74 $Y=0.19 $X2=3.765
+ $Y2=0.56
cc_93 N_GND_M1006_b N_A_570_115#_c_672_n 0.0145317f $X=-0.045 $Y=0 $X2=3.075
+ $Y2=0.56
cc_94 N_GND_c_9_p N_A_570_115#_c_672_n 0.0062002f $X=2.56 $Y=0.74 $X2=3.075
+ $Y2=0.56
cc_95 N_GND_c_4_p N_A_570_115#_c_672_n 0.00506617f $X=3.74 $Y=0.19 $X2=3.075
+ $Y2=0.56
cc_96 N_VDD_M1003_b N_CON_M1003_g 0.0752803f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=4.195
cc_97 N_VDD_c_97_p N_CON_M1003_g 0.00496961f $X=0.665 $Y=5.397 $X2=0.475
+ $Y2=4.195
cc_98 N_VDD_c_98_p N_CON_M1003_g 0.0195001f $X=0.75 $Y=3.215 $X2=0.475 $Y2=4.195
cc_99 N_VDD_c_99_p N_CON_M1003_g 0.00429146f $X=3.74 $Y=5.36 $X2=0.475 $Y2=4.195
cc_100 N_VDD_M1003_b N_CON_c_179_n 0.00290115f $X=-0.045 $Y=2.645 $X2=2.62
+ $Y2=3.215
cc_101 N_VDD_c_101_p N_CON_c_179_n 0.00469914f $X=2.965 $Y=5.397 $X2=2.62
+ $Y2=3.215
cc_102 N_VDD_c_99_p N_CON_c_179_n 0.00435496f $X=3.74 $Y=5.36 $X2=2.62 $Y2=3.215
cc_103 N_VDD_M1003_b N_CON_c_164_n 0.0218832f $X=-0.045 $Y=2.645 $X2=3.755
+ $Y2=2.69
cc_104 N_VDD_c_104_p N_CON_c_164_n 0.0121906f $X=3.05 $Y=3.215 $X2=3.755
+ $Y2=2.69
cc_105 N_VDD_M1003_b N_CON_c_184_n 0.00419737f $X=-0.045 $Y=2.645 $X2=3.84
+ $Y2=3.215
cc_106 N_VDD_c_106_p N_CON_c_184_n 0.00452684f $X=3.74 $Y=5.33 $X2=3.84
+ $Y2=3.215
cc_107 N_VDD_c_99_p N_CON_c_184_n 0.00435496f $X=3.74 $Y=5.36 $X2=3.84 $Y2=3.215
cc_108 N_VDD_M1003_b N_CON_c_167_n 0.00108117f $X=-0.045 $Y=2.645 $X2=2.62
+ $Y2=2.69
cc_109 N_VDD_M1003_b N_B_M1010_g 0.0216302f $X=-0.045 $Y=2.645 $X2=0.965
+ $Y2=3.825
cc_110 N_VDD_c_98_p N_B_M1010_g 0.00373151f $X=0.75 $Y=3.215 $X2=0.965 $Y2=3.825
cc_111 N_VDD_c_111_p N_B_M1010_g 0.00496961f $X=1.525 $Y=5.397 $X2=0.965
+ $Y2=3.825
cc_112 N_VDD_c_99_p N_B_M1010_g 0.00429146f $X=3.74 $Y=5.36 $X2=0.965 $Y2=3.825
cc_113 N_VDD_M1003_b N_B_M1013_g 0.0185755f $X=-0.045 $Y=2.645 $X2=3.265
+ $Y2=3.825
cc_114 N_VDD_c_104_p N_B_M1013_g 0.00354579f $X=3.05 $Y=3.215 $X2=3.265
+ $Y2=3.825
cc_115 N_VDD_c_106_p N_B_M1013_g 0.00496961f $X=3.74 $Y=5.33 $X2=3.265 $Y2=3.825
cc_116 N_VDD_c_99_p N_B_M1013_g 0.00429146f $X=3.74 $Y=5.36 $X2=3.265 $Y2=3.825
cc_117 N_VDD_M1003_b N_A_M1011_g 0.0197771f $X=-0.045 $Y=2.645 $X2=1.395
+ $Y2=3.825
cc_118 N_VDD_c_111_p N_A_M1011_g 0.00496961f $X=1.525 $Y=5.397 $X2=1.395
+ $Y2=3.825
cc_119 N_VDD_c_119_p N_A_M1011_g 0.00373151f $X=1.61 $Y=3.555 $X2=1.395
+ $Y2=3.825
cc_120 N_VDD_c_99_p N_A_M1011_g 0.00429146f $X=3.74 $Y=5.36 $X2=1.395 $Y2=3.825
cc_121 N_VDD_M1003_b N_A_M1000_g 0.0243418f $X=-0.045 $Y=2.645 $X2=3.625
+ $Y2=3.825
cc_122 N_VDD_c_106_p N_A_M1000_g 0.00496961f $X=3.74 $Y=5.33 $X2=3.625 $Y2=3.825
cc_123 N_VDD_c_99_p N_A_M1000_g 0.00429146f $X=3.74 $Y=5.36 $X2=3.625 $Y2=3.825
cc_124 N_VDD_M1003_b N_A_208_565#_M1012_g 0.0679203f $X=-0.045 $Y=2.645
+ $X2=1.885 $Y2=4.195
cc_125 N_VDD_c_119_p N_A_208_565#_M1012_g 0.0162477f $X=1.61 $Y=3.555 $X2=1.885
+ $Y2=4.195
cc_126 N_VDD_c_101_p N_A_208_565#_M1012_g 0.00496961f $X=2.965 $Y=5.397
+ $X2=1.885 $Y2=4.195
cc_127 N_VDD_c_99_p N_A_208_565#_M1012_g 0.00429146f $X=3.74 $Y=5.36 $X2=1.885
+ $Y2=4.195
cc_128 N_VDD_M1003_b N_A_208_565#_M1002_g 0.0252169f $X=-0.045 $Y=2.645
+ $X2=2.835 $Y2=3.825
cc_129 N_VDD_c_101_p N_A_208_565#_M1002_g 0.00496961f $X=2.965 $Y=5.397
+ $X2=2.835 $Y2=3.825
cc_130 N_VDD_c_104_p N_A_208_565#_M1002_g 0.00354579f $X=3.05 $Y=3.215 $X2=2.835
+ $Y2=3.825
cc_131 N_VDD_c_99_p N_A_208_565#_M1002_g 0.00429146f $X=3.74 $Y=5.36 $X2=2.835
+ $Y2=3.825
cc_132 N_VDD_M1003_b N_A_208_565#_c_501_n 0.00198641f $X=-0.045 $Y=2.645
+ $X2=1.18 $Y2=3.555
cc_133 N_VDD_c_111_p N_A_208_565#_c_501_n 0.00456907f $X=1.525 $Y=5.397 $X2=1.18
+ $Y2=3.555
cc_134 N_VDD_c_99_p N_A_208_565#_c_501_n 0.00434939f $X=3.74 $Y=5.36 $X2=1.18
+ $Y2=3.555
cc_135 N_VDD_M1011_d N_A_208_565#_c_504_n 0.00483849f $X=1.47 $Y=2.825 $X2=1.64
+ $Y2=2.75
cc_136 N_VDD_M1003_b N_A_208_565#_c_504_n 0.00578065f $X=-0.045 $Y=2.645
+ $X2=1.64 $Y2=2.75
cc_137 N_VDD_c_119_p N_A_208_565#_c_504_n 0.00659105f $X=1.61 $Y=3.555 $X2=1.64
+ $Y2=2.75
cc_138 N_VDD_M1003_b N_A_208_565#_c_507_n 0.00518782f $X=-0.045 $Y=2.645
+ $X2=1.265 $Y2=2.75
cc_139 N_VDD_M1003_b N_A_208_565#_c_491_n 3.89739e-19 $X=-0.045 $Y=2.645
+ $X2=1.725 $Y2=2.665
cc_140 N_VDD_M1003_b N_S_c_593_n 0.027267f $X=-0.045 $Y=2.645 $X2=0.26 $Y2=3.07
cc_141 N_VDD_c_97_p N_S_c_593_n 0.00452684f $X=0.665 $Y=5.397 $X2=0.26 $Y2=3.07
cc_142 N_VDD_c_98_p N_S_c_593_n 0.0532241f $X=0.75 $Y=3.215 $X2=0.26 $Y2=3.07
cc_143 N_VDD_c_99_p N_S_c_593_n 0.00435496f $X=3.74 $Y=5.36 $X2=0.26 $Y2=3.07
cc_144 N_VDD_M1003_b S 0.0165608f $X=-0.045 $Y=2.645 $X2=0.25 $Y2=2.125
cc_145 N_VDD_M1003_b N_S_c_598_n 0.0173138f $X=-0.045 $Y=2.645 $X2=0.26 $Y2=3.07
cc_146 N_VDD_c_98_p N_S_c_598_n 0.0056248f $X=0.75 $Y=3.215 $X2=0.26 $Y2=3.07
cc_147 N_VDD_M1003_b N_CO_c_625_n 0.0206443f $X=-0.045 $Y=2.645 $X2=2.1
+ $Y2=3.895
cc_148 N_VDD_c_119_p N_CO_c_625_n 0.0409245f $X=1.61 $Y=3.555 $X2=2.1 $Y2=3.895
cc_149 N_VDD_c_101_p N_CO_c_625_n 0.00475705f $X=2.965 $Y=5.397 $X2=2.1
+ $Y2=3.895
cc_150 N_VDD_c_99_p N_CO_c_625_n 0.00435496f $X=3.74 $Y=5.36 $X2=2.1 $Y2=3.895
cc_151 N_VDD_M1003_b N_CO_c_622_n 0.00360959f $X=-0.045 $Y=2.645 $X2=2.175
+ $Y2=2.7
cc_152 N_VDD_M1003_b CO 0.0105263f $X=-0.045 $Y=2.645 $X2=2.175 $Y2=2.7
cc_153 N_CON_M1006_g N_B_M1007_g 0.033689f $X=0.475 $Y=0.85 $X2=0.965 $Y2=0.995
cc_154 N_CON_c_159_n N_B_M1007_g 0.00317949f $X=0.635 $Y=1.59 $X2=0.965
+ $Y2=0.995
cc_155 N_CON_c_168_n N_B_M1007_g 0.0103705f $X=2.475 $Y=1.59 $X2=0.965 $Y2=0.995
cc_156 N_CON_c_170_n N_B_M1007_g 9.80511e-19 $X=0.78 $Y=1.59 $X2=0.965 $Y2=0.995
cc_157 N_CON_M1003_g N_B_M1010_g 0.0622958f $X=0.475 $Y=4.195 $X2=0.965
+ $Y2=3.825
cc_158 N_CON_c_162_n N_B_M1004_g 0.00298059f $X=2.62 $Y=2.605 $X2=3.205
+ $Y2=0.995
cc_159 N_CON_c_163_n N_B_M1004_g 0.0120887f $X=3.335 $Y=1.59 $X2=3.205 $Y2=0.995
cc_160 N_CON_c_166_n N_B_M1004_g 0.00288927f $X=3.42 $Y=1.065 $X2=3.205
+ $Y2=0.995
cc_161 N_CON_c_172_n N_B_M1004_g 4.76806e-19 $X=2.62 $Y=1.59 $X2=3.205 $Y2=0.995
cc_162 CON N_B_M1004_g 0.00638136f $X=3.42 $Y=1.59 $X2=3.205 $Y2=0.995
cc_163 N_CON_c_162_n N_B_M1013_g 0.00509671f $X=2.62 $Y=2.605 $X2=3.265
+ $Y2=3.825
cc_164 N_CON_c_164_n N_B_M1013_g 0.0160357f $X=3.755 $Y=2.69 $X2=3.265 $Y2=3.825
cc_165 N_CON_M1003_g N_B_c_290_n 0.0198105f $X=0.475 $Y=4.195 $X2=0.905 $Y2=1.96
cc_166 N_CON_c_168_n N_B_c_290_n 0.0017113f $X=2.475 $Y=1.59 $X2=0.905 $Y2=1.96
cc_167 N_CON_c_162_n N_B_c_292_n 0.00527976f $X=2.62 $Y=2.605 $X2=3.205 $Y2=1.96
cc_168 N_CON_c_163_n N_B_c_292_n 0.00297725f $X=3.335 $Y=1.59 $X2=3.205 $Y2=1.96
cc_169 N_CON_c_164_n N_B_c_292_n 0.00235541f $X=3.755 $Y=2.69 $X2=3.205 $Y2=1.96
cc_170 CON N_B_c_292_n 0.00117979f $X=3.42 $Y=1.59 $X2=3.205 $Y2=1.96
cc_171 N_CON_M1003_g N_B_c_293_n 0.00376362f $X=0.475 $Y=4.195 $X2=0.905
+ $Y2=1.96
cc_172 N_CON_c_168_n N_B_c_293_n 0.00349538f $X=2.475 $Y=1.59 $X2=0.905 $Y2=1.96
cc_173 N_CON_c_170_n N_B_c_293_n 7.89715e-19 $X=0.78 $Y=1.59 $X2=0.905 $Y2=1.96
cc_174 N_CON_c_162_n N_B_c_295_n 0.00612449f $X=2.62 $Y=2.605 $X2=3.205 $Y2=1.96
cc_175 N_CON_c_163_n N_B_c_295_n 0.0159093f $X=3.335 $Y=1.59 $X2=3.205 $Y2=1.96
cc_176 N_CON_c_164_n N_B_c_295_n 0.00416532f $X=3.755 $Y=2.69 $X2=3.205 $Y2=1.96
cc_177 N_CON_c_165_n N_B_c_295_n 0.00205373f $X=3.42 $Y=1.505 $X2=3.205 $Y2=1.96
cc_178 CON N_B_c_295_n 9.81883e-19 $X=3.42 $Y=1.59 $X2=3.205 $Y2=1.96
cc_179 N_CON_M1003_g N_B_c_296_n 3.21736e-19 $X=0.475 $Y=4.195 $X2=1.05 $Y2=1.96
cc_180 N_CON_c_168_n N_B_c_296_n 0.024704f $X=2.475 $Y=1.59 $X2=1.05 $Y2=1.96
cc_181 N_CON_c_170_n N_B_c_296_n 0.00206194f $X=0.78 $Y=1.59 $X2=1.05 $Y2=1.96
cc_182 N_CON_c_162_n N_B_c_297_n 0.0139114f $X=2.62 $Y=2.605 $X2=3.06 $Y2=1.96
cc_183 N_CON_c_163_n N_B_c_297_n 0.0132985f $X=3.335 $Y=1.59 $X2=3.06 $Y2=1.96
cc_184 N_CON_c_168_n N_B_c_297_n 0.116608f $X=2.475 $Y=1.59 $X2=3.06 $Y2=1.96
cc_185 N_CON_c_172_n N_B_c_297_n 0.0254758f $X=2.62 $Y=1.59 $X2=3.06 $Y2=1.96
cc_186 N_CON_c_162_n B 0.00223952f $X=2.62 $Y=2.605 $X2=3.21 $Y2=1.96
cc_187 N_CON_c_163_n B 0.00321159f $X=3.335 $Y=1.59 $X2=3.21 $Y2=1.96
cc_188 CON B 0.0176994f $X=3.42 $Y=1.59 $X2=3.21 $Y2=1.96
cc_189 N_CON_c_168_n N_A_M1008_g 0.0102813f $X=2.475 $Y=1.59 $X2=1.325 $Y2=0.995
cc_190 N_CON_c_164_n N_A_M1000_g 0.015762f $X=3.755 $Y=2.69 $X2=3.625 $Y2=3.825
cc_191 N_CON_c_184_n N_A_M1000_g 0.00669003f $X=3.84 $Y=3.215 $X2=3.625
+ $Y2=3.825
cc_192 N_CON_c_165_n N_A_M1005_g 0.00402015f $X=3.42 $Y=1.505 $X2=3.635
+ $Y2=0.995
cc_193 N_CON_c_166_n N_A_M1005_g 0.00288927f $X=3.42 $Y=1.065 $X2=3.635
+ $Y2=0.995
cc_194 CON N_A_M1005_g 0.010636f $X=3.42 $Y=1.59 $X2=3.635 $Y2=0.995
cc_195 N_CON_c_164_n N_A_c_392_n 0.00303009f $X=3.755 $Y=2.69 $X2=3.685 $Y2=2.33
cc_196 N_CON_c_164_n N_A_c_394_n 0.0189273f $X=3.755 $Y=2.69 $X2=3.685 $Y2=2.33
cc_197 CON N_A_c_394_n 3.86961e-19 $X=3.42 $Y=1.59 $X2=3.685 $Y2=2.33
cc_198 N_CON_c_164_n A 0.00711502f $X=3.755 $Y=2.69 $X2=3.685 $Y2=2.33
cc_199 CON A 0.00132366f $X=3.42 $Y=1.59 $X2=3.685 $Y2=2.33
cc_200 N_CON_c_162_n N_A_c_397_n 0.0228953f $X=2.62 $Y=2.605 $X2=3.54 $Y2=2.33
cc_201 N_CON_c_164_n N_A_c_397_n 0.0305931f $X=3.755 $Y=2.69 $X2=3.54 $Y2=2.33
cc_202 N_CON_c_165_n N_A_c_397_n 8.38986e-19 $X=3.42 $Y=1.505 $X2=3.54 $Y2=2.33
cc_203 CON N_A_c_397_n 0.0098042f $X=3.42 $Y=1.59 $X2=3.54 $Y2=2.33
cc_204 N_CON_c_168_n N_A_208_565#_c_471_n 0.0103721f $X=2.475 $Y=1.59 $X2=1.885
+ $Y2=1.86
cc_205 N_CON_c_168_n N_A_208_565#_c_474_n 0.00229041f $X=2.475 $Y=1.59 $X2=2.21
+ $Y2=1.565
cc_206 N_CON_c_162_n N_A_208_565#_c_475_n 0.0141245f $X=2.62 $Y=2.605 $X2=2.76
+ $Y2=2.41
cc_207 N_CON_c_163_n N_A_208_565#_c_475_n 0.00257529f $X=3.335 $Y=1.59 $X2=2.76
+ $Y2=2.41
cc_208 N_CON_c_172_n N_A_208_565#_M1001_g 2.41495e-19 $X=2.62 $Y=1.59 $X2=2.285
+ $Y2=0.895
cc_209 N_CON_c_161_n N_A_208_565#_c_480_n 0.00929899f $X=2.62 $Y=1.675 $X2=2.7
+ $Y2=1.565
cc_210 N_CON_c_163_n N_A_208_565#_c_480_n 0.0101401f $X=3.335 $Y=1.59 $X2=2.7
+ $Y2=1.565
cc_211 N_CON_c_168_n N_A_208_565#_c_480_n 0.00553403f $X=2.475 $Y=1.59 $X2=2.7
+ $Y2=1.565
cc_212 N_CON_c_172_n N_A_208_565#_c_480_n 0.00162604f $X=2.62 $Y=1.59 $X2=2.7
+ $Y2=1.565
cc_213 N_CON_c_172_n N_A_208_565#_c_482_n 0.00294886f $X=2.62 $Y=1.59 $X2=2.775
+ $Y2=1.49
cc_214 N_CON_c_162_n N_A_208_565#_M1002_g 0.0046186f $X=2.62 $Y=2.605 $X2=2.835
+ $Y2=3.825
cc_215 N_CON_c_179_n N_A_208_565#_M1002_g 0.00669003f $X=2.62 $Y=3.215 $X2=2.835
+ $Y2=3.825
cc_216 N_CON_c_164_n N_A_208_565#_M1002_g 0.0162813f $X=3.755 $Y=2.69 $X2=2.835
+ $Y2=3.825
cc_217 N_CON_c_168_n N_A_208_565#_c_487_n 0.00467421f $X=2.475 $Y=1.59 $X2=2.285
+ $Y2=1.565
cc_218 N_CON_c_168_n N_A_208_565#_c_488_n 0.0108903f $X=2.475 $Y=1.59 $X2=1.54
+ $Y2=0.74
cc_219 N_CON_c_168_n N_A_208_565#_c_492_n 0.0233954f $X=2.475 $Y=1.59 $X2=1.725
+ $Y2=1.695
cc_220 N_CON_M1006_g N_S_c_586_n 0.00734808f $X=0.475 $Y=0.85 $X2=0.26 $Y2=0.825
cc_221 N_CON_c_158_n N_S_c_586_n 0.00243007f $X=0.35 $Y=1.59 $X2=0.26 $Y2=0.825
cc_222 N_CON_c_159_n N_S_c_586_n 0.00919709f $X=0.635 $Y=1.59 $X2=0.26 $Y2=0.825
cc_223 N_CON_M1003_g N_S_c_593_n 0.0168927f $X=0.475 $Y=4.195 $X2=0.26 $Y2=3.07
cc_224 N_CON_M1006_g S 0.00219688f $X=0.475 $Y=0.85 $X2=0.25 $Y2=2.125
cc_225 N_CON_M1003_g S 0.026126f $X=0.475 $Y=4.195 $X2=0.25 $Y2=2.125
cc_226 N_CON_c_158_n S 0.0074247f $X=0.35 $Y=1.59 $X2=0.25 $Y2=2.125
cc_227 N_CON_c_159_n S 0.0144314f $X=0.635 $Y=1.59 $X2=0.25 $Y2=2.125
cc_228 N_CON_c_170_n S 0.0220567f $X=0.78 $Y=1.59 $X2=0.25 $Y2=2.125
cc_229 N_CON_M1006_g N_S_c_591_n 0.00595114f $X=0.475 $Y=0.85 $X2=0.26 $Y2=1.215
cc_230 N_CON_c_158_n N_S_c_591_n 0.00148757f $X=0.35 $Y=1.59 $X2=0.26 $Y2=1.215
cc_231 N_CON_c_159_n N_S_c_591_n 0.00260285f $X=0.635 $Y=1.59 $X2=0.26 $Y2=1.215
cc_232 N_CON_M1003_g N_S_c_598_n 0.0054567f $X=0.475 $Y=4.195 $X2=0.26 $Y2=3.07
cc_233 N_CON_c_179_n N_CO_c_625_n 0.0878891f $X=2.62 $Y=3.215 $X2=2.1 $Y2=3.895
cc_234 N_CON_c_168_n N_CO_c_620_n 0.00506454f $X=2.475 $Y=1.59 $X2=2.175
+ $Y2=1.215
cc_235 N_CON_c_179_n N_CO_c_622_n 3.73019e-19 $X=2.62 $Y=3.215 $X2=2.175 $Y2=2.7
cc_236 N_CON_c_161_n N_CO_c_623_n 0.00670709f $X=2.62 $Y=1.675 $X2=2.137
+ $Y2=2.615
cc_237 N_CON_c_162_n N_CO_c_623_n 0.0448782f $X=2.62 $Y=2.605 $X2=2.137
+ $Y2=2.615
cc_238 N_CON_c_167_n N_CO_c_623_n 0.00730853f $X=2.62 $Y=2.69 $X2=2.137
+ $Y2=2.615
cc_239 N_CON_c_168_n N_CO_c_623_n 0.0121795f $X=2.475 $Y=1.59 $X2=2.137
+ $Y2=2.615
cc_240 N_CON_c_172_n N_CO_c_623_n 0.00207393f $X=2.62 $Y=1.59 $X2=2.137
+ $Y2=2.615
cc_241 N_CON_c_162_n CO 5.70376e-19 $X=2.62 $Y=2.605 $X2=2.175 $Y2=2.7
cc_242 N_CON_c_179_n CO 0.00122973f $X=2.62 $Y=3.215 $X2=2.175 $Y2=2.7
cc_243 N_CON_c_167_n CO 0.00605606f $X=2.62 $Y=2.69 $X2=2.175 $Y2=2.7
cc_244 N_CON_c_163_n N_A_570_115#_c_675_n 0.0101003f $X=3.335 $Y=1.59 $X2=2.99
+ $Y2=0.74
cc_245 N_CON_M1004_d N_A_570_115#_c_670_n 0.00176461f $X=3.28 $Y=0.575 $X2=3.765
+ $Y2=0.56
cc_246 N_CON_c_166_n N_A_570_115#_c_670_n 0.0130031f $X=3.42 $Y=1.065 $X2=3.765
+ $Y2=0.56
cc_247 N_B_M1007_g N_A_M1008_g 0.0639188f $X=0.965 $Y=0.995 $X2=1.325 $Y2=0.995
cc_248 N_B_c_293_n N_A_M1008_g 0.00121678f $X=0.905 $Y=1.96 $X2=1.325 $Y2=0.995
cc_249 N_B_c_296_n N_A_M1008_g 7.94897e-19 $X=1.05 $Y=1.96 $X2=1.325 $Y2=0.995
cc_250 N_B_c_297_n N_A_M1008_g 0.00595709f $X=3.06 $Y=1.96 $X2=1.325 $Y2=0.995
cc_251 N_B_M1010_g N_A_M1011_g 0.0405421f $X=0.965 $Y=3.825 $X2=1.395 $Y2=3.825
cc_252 N_B_M1004_g N_A_M1005_g 0.0414265f $X=3.205 $Y=0.995 $X2=3.635 $Y2=0.995
cc_253 N_B_c_292_n N_A_M1005_g 0.022402f $X=3.205 $Y=1.96 $X2=3.635 $Y2=0.995
cc_254 N_B_c_295_n N_A_M1005_g 0.00376362f $X=3.205 $Y=1.96 $X2=3.635 $Y2=0.995
cc_255 B N_A_M1005_g 9.23221e-19 $X=3.21 $Y=1.96 $X2=3.635 $Y2=0.995
cc_256 N_B_c_290_n N_A_c_391_n 0.0639188f $X=0.905 $Y=1.96 $X2=1.385 $Y2=2.33
cc_257 N_B_c_297_n N_A_c_391_n 7.99243e-19 $X=3.06 $Y=1.96 $X2=1.385 $Y2=2.33
cc_258 N_B_M1013_g N_A_c_392_n 0.168643f $X=3.265 $Y=3.825 $X2=3.685 $Y2=2.33
cc_259 N_B_M1010_g N_A_c_393_n 0.00286993f $X=0.965 $Y=3.825 $X2=1.385 $Y2=2.33
cc_260 N_B_c_297_n N_A_c_393_n 0.00428104f $X=3.06 $Y=1.96 $X2=1.385 $Y2=2.33
cc_261 N_B_M1013_g N_A_c_394_n 0.00278747f $X=3.265 $Y=3.825 $X2=3.685 $Y2=2.33
cc_262 N_B_M1010_g N_A_c_395_n 0.00405562f $X=0.965 $Y=3.825 $X2=1.53 $Y2=2.33
cc_263 N_B_c_297_n N_A_c_395_n 0.0263377f $X=3.06 $Y=1.96 $X2=1.53 $Y2=2.33
cc_264 N_B_M1013_g A 7.94897e-19 $X=3.265 $Y=3.825 $X2=3.685 $Y2=2.33
cc_265 N_B_M1013_g N_A_c_397_n 0.00633265f $X=3.265 $Y=3.825 $X2=3.54 $Y2=2.33
cc_266 N_B_c_292_n N_A_c_397_n 0.00210214f $X=3.205 $Y=1.96 $X2=3.54 $Y2=2.33
cc_267 N_B_c_295_n N_A_c_397_n 0.00225835f $X=3.205 $Y=1.96 $X2=3.54 $Y2=2.33
cc_268 N_B_c_297_n N_A_c_397_n 0.128931f $X=3.06 $Y=1.96 $X2=3.54 $Y2=2.33
cc_269 B N_A_c_397_n 0.0270107f $X=3.21 $Y=1.96 $X2=3.54 $Y2=2.33
cc_270 N_B_c_297_n N_A_208_565#_c_472_n 0.00725075f $X=3.06 $Y=1.96 $X2=1.885
+ $Y2=2.335
cc_271 N_B_c_297_n N_A_208_565#_c_474_n 0.00119779f $X=3.06 $Y=1.96 $X2=2.21
+ $Y2=1.565
cc_272 N_B_M1013_g N_A_208_565#_c_475_n 0.0381911f $X=3.265 $Y=3.825 $X2=2.76
+ $Y2=2.41
cc_273 N_B_c_297_n N_A_208_565#_c_475_n 0.00176131f $X=3.06 $Y=1.96 $X2=2.76
+ $Y2=2.41
cc_274 N_B_M1004_g N_A_208_565#_c_482_n 0.022187f $X=3.205 $Y=0.995 $X2=2.775
+ $Y2=1.49
cc_275 N_B_M1010_g N_A_208_565#_c_507_n 0.00507079f $X=0.965 $Y=3.825 $X2=1.265
+ $Y2=2.75
cc_276 N_B_c_297_n N_A_208_565#_c_507_n 0.0051538f $X=3.06 $Y=1.96 $X2=1.265
+ $Y2=2.75
cc_277 N_B_c_293_n N_A_208_565#_c_491_n 0.00316158f $X=0.905 $Y=1.96 $X2=1.725
+ $Y2=2.665
cc_278 N_B_c_296_n N_A_208_565#_c_491_n 0.00129846f $X=1.05 $Y=1.96 $X2=1.725
+ $Y2=2.665
cc_279 N_B_c_297_n N_A_208_565#_c_491_n 0.0153226f $X=3.06 $Y=1.96 $X2=1.725
+ $Y2=2.665
cc_280 N_B_c_296_n N_A_208_565#_c_492_n 5.15761e-19 $X=1.05 $Y=1.96 $X2=1.725
+ $Y2=1.695
cc_281 N_B_c_297_n N_A_208_565#_c_492_n 0.00890945f $X=3.06 $Y=1.96 $X2=1.725
+ $Y2=1.695
cc_282 N_B_M1007_g S 4.21151e-19 $X=0.965 $Y=0.995 $X2=0.25 $Y2=2.125
cc_283 N_B_c_293_n S 0.00429487f $X=0.905 $Y=1.96 $X2=0.25 $Y2=2.125
cc_284 N_B_c_296_n S 0.0134542f $X=1.05 $Y=1.96 $X2=0.25 $Y2=2.125
cc_285 N_B_M1007_g N_S_c_591_n 3.27178e-19 $X=0.965 $Y=0.995 $X2=0.26 $Y2=1.215
cc_286 N_B_c_297_n N_CO_c_623_n 0.0136552f $X=3.06 $Y=1.96 $X2=2.137 $Y2=2.615
cc_287 N_B_M1004_g N_A_570_115#_c_670_n 0.012637f $X=3.205 $Y=0.995 $X2=3.765
+ $Y2=0.56
cc_288 N_A_M1008_g N_A_208_565#_c_471_n 0.0164301f $X=1.325 $Y=0.995 $X2=1.885
+ $Y2=1.86
cc_289 N_A_M1008_g N_A_208_565#_c_472_n 0.00833244f $X=1.325 $Y=0.995 $X2=1.885
+ $Y2=2.335
cc_290 N_A_c_391_n N_A_208_565#_c_472_n 0.0147848f $X=1.385 $Y=2.33 $X2=1.885
+ $Y2=2.335
cc_291 N_A_c_397_n N_A_208_565#_c_472_n 0.00210973f $X=3.54 $Y=2.33 $X2=1.885
+ $Y2=2.335
cc_292 N_A_M1011_g N_A_208_565#_M1012_g 0.0513848f $X=1.395 $Y=3.825 $X2=1.885
+ $Y2=4.195
cc_293 N_A_c_397_n N_A_208_565#_c_475_n 0.0139241f $X=3.54 $Y=2.33 $X2=2.76
+ $Y2=2.41
cc_294 N_A_c_397_n N_A_208_565#_c_486_n 0.00700381f $X=3.54 $Y=2.33 $X2=1.885
+ $Y2=2.41
cc_295 N_A_M1011_g N_A_208_565#_c_504_n 0.0147914f $X=1.395 $Y=3.825 $X2=1.64
+ $Y2=2.75
cc_296 N_A_c_391_n N_A_208_565#_c_504_n 0.00348735f $X=1.385 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_297 N_A_c_393_n N_A_208_565#_c_504_n 0.0111584f $X=1.385 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_298 N_A_c_395_n N_A_208_565#_c_504_n 0.00509311f $X=1.53 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_299 N_A_c_397_n N_A_208_565#_c_504_n 0.00467069f $X=3.54 $Y=2.33 $X2=1.64
+ $Y2=2.75
cc_300 N_A_c_391_n N_A_208_565#_c_507_n 7.25782e-19 $X=1.385 $Y=2.33 $X2=1.265
+ $Y2=2.75
cc_301 N_A_c_395_n N_A_208_565#_c_507_n 0.00124978f $X=1.53 $Y=2.33 $X2=1.265
+ $Y2=2.75
cc_302 N_A_M1008_g N_A_208_565#_c_488_n 0.00607295f $X=1.325 $Y=0.995 $X2=1.54
+ $Y2=0.74
cc_303 N_A_M1008_g N_A_208_565#_c_491_n 0.00392362f $X=1.325 $Y=0.995 $X2=1.725
+ $Y2=2.665
cc_304 N_A_M1011_g N_A_208_565#_c_491_n 0.00360042f $X=1.395 $Y=3.825 $X2=1.725
+ $Y2=2.665
cc_305 N_A_c_391_n N_A_208_565#_c_491_n 0.00193142f $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_306 N_A_c_393_n N_A_208_565#_c_491_n 0.0224238f $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_307 N_A_c_395_n N_A_208_565#_c_491_n 0.00168305f $X=1.53 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_308 N_A_c_397_n N_A_208_565#_c_491_n 0.0185059f $X=3.54 $Y=2.33 $X2=1.725
+ $Y2=2.665
cc_309 N_A_M1008_g N_A_208_565#_c_492_n 0.00736605f $X=1.325 $Y=0.995 $X2=1.725
+ $Y2=1.695
cc_310 N_A_c_391_n N_A_208_565#_c_492_n 0.00175929f $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=1.695
cc_311 N_A_c_393_n N_A_208_565#_c_492_n 2.52704e-19 $X=1.385 $Y=2.33 $X2=1.725
+ $Y2=1.695
cc_312 N_A_c_397_n N_CO_c_622_n 0.00105312f $X=3.54 $Y=2.33 $X2=2.175 $Y2=2.7
cc_313 N_A_c_397_n N_CO_c_623_n 0.0133702f $X=3.54 $Y=2.33 $X2=2.137 $Y2=2.615
cc_314 N_A_c_397_n CO 0.0346374f $X=3.54 $Y=2.33 $X2=2.175 $Y2=2.7
cc_315 N_A_M1005_g N_A_570_115#_c_670_n 0.0135957f $X=3.635 $Y=0.995 $X2=3.765
+ $Y2=0.56
cc_316 N_A_208_565#_c_488_n N_CO_c_617_n 0.0232208f $X=1.54 $Y=0.74 $X2=2.07
+ $Y2=0.825
cc_317 N_A_208_565#_c_474_n N_CO_c_620_n 0.00410169f $X=2.21 $Y=1.565 $X2=2.175
+ $Y2=1.215
cc_318 N_A_208_565#_M1001_g N_CO_c_620_n 0.00814843f $X=2.285 $Y=0.895 $X2=2.175
+ $Y2=1.215
cc_319 N_A_208_565#_c_482_n N_CO_c_620_n 2.32977e-19 $X=2.775 $Y=1.49 $X2=2.175
+ $Y2=1.215
cc_320 N_A_208_565#_c_488_n N_CO_c_620_n 0.00744736f $X=1.54 $Y=0.74 $X2=2.175
+ $Y2=1.215
cc_321 N_A_208_565#_M1012_g N_CO_c_622_n 0.0331071f $X=1.885 $Y=4.195 $X2=2.175
+ $Y2=2.7
cc_322 N_A_208_565#_c_475_n N_CO_c_622_n 0.00140819f $X=2.76 $Y=2.41 $X2=2.175
+ $Y2=2.7
cc_323 N_A_208_565#_c_504_n N_CO_c_622_n 0.0107786f $X=1.64 $Y=2.75 $X2=2.175
+ $Y2=2.7
cc_324 N_A_208_565#_c_491_n N_CO_c_622_n 0.00298908f $X=1.725 $Y=2.665 $X2=2.175
+ $Y2=2.7
cc_325 N_A_208_565#_c_471_n N_CO_c_623_n 0.0106746f $X=1.885 $Y=1.86 $X2=2.137
+ $Y2=2.615
cc_326 N_A_208_565#_M1012_g N_CO_c_623_n 0.00273706f $X=1.885 $Y=4.195 $X2=2.137
+ $Y2=2.615
cc_327 N_A_208_565#_c_474_n N_CO_c_623_n 0.00787523f $X=2.21 $Y=1.565 $X2=2.137
+ $Y2=2.615
cc_328 N_A_208_565#_c_475_n N_CO_c_623_n 0.0137108f $X=2.76 $Y=2.41 $X2=2.137
+ $Y2=2.615
cc_329 N_A_208_565#_M1001_g N_CO_c_623_n 0.00669606f $X=2.285 $Y=0.895 $X2=2.137
+ $Y2=2.615
cc_330 N_A_208_565#_c_482_n N_CO_c_623_n 9.34664e-19 $X=2.775 $Y=1.49 $X2=2.137
+ $Y2=2.615
cc_331 N_A_208_565#_M1002_g N_CO_c_623_n 8.14457e-19 $X=2.835 $Y=3.825 $X2=2.137
+ $Y2=2.615
cc_332 N_A_208_565#_c_487_n N_CO_c_623_n 0.0035441f $X=2.285 $Y=1.565 $X2=2.137
+ $Y2=2.615
cc_333 N_A_208_565#_c_488_n N_CO_c_623_n 0.00797516f $X=1.54 $Y=0.74 $X2=2.137
+ $Y2=2.615
cc_334 N_A_208_565#_c_491_n N_CO_c_623_n 0.0354244f $X=1.725 $Y=2.665 $X2=2.137
+ $Y2=2.615
cc_335 N_A_208_565#_c_492_n N_CO_c_623_n 0.0222011f $X=1.725 $Y=1.695 $X2=2.137
+ $Y2=2.615
cc_336 N_A_208_565#_M1012_g CO 7.58429e-19 $X=1.885 $Y=4.195 $X2=2.175 $Y2=2.7
cc_337 N_A_208_565#_c_475_n CO 0.0027071f $X=2.76 $Y=2.41 $X2=2.175 $Y2=2.7
cc_338 N_A_208_565#_c_504_n CO 0.00111652f $X=1.64 $Y=2.75 $X2=2.175 $Y2=2.7
cc_339 N_A_208_565#_c_491_n CO 0.0012063f $X=1.725 $Y=2.665 $X2=2.175 $Y2=2.7
cc_340 N_A_208_565#_c_482_n N_A_570_115#_c_672_n 9.82882e-19 $X=2.775 $Y=1.49
+ $X2=3.075 $Y2=0.56
