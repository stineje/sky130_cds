magic
tech sky130A
magscale 1 2
timestamp 1612373886
<< nwell >>
rect -9 529 638 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 238 115 268 243
rect 358 115 388 243
rect 430 115 460 243
rect 516 115 546 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 238 565 268 965
rect 358 565 388 965
rect 430 565 460 965
rect 516 565 546 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 165 166 243
rect 110 131 121 165
rect 155 131 166 165
rect 110 115 166 131
rect 196 115 238 243
rect 268 215 358 243
rect 268 131 279 215
rect 347 131 358 215
rect 268 115 358 131
rect 388 115 430 243
rect 460 165 516 243
rect 460 131 471 165
rect 505 131 516 165
rect 460 115 516 131
rect 546 215 599 243
rect 546 131 557 215
rect 591 131 599 215
rect 546 115 599 131
<< pdiff >>
rect 27 949 80 965
rect 27 605 35 949
rect 69 605 80 949
rect 27 565 80 605
rect 110 949 166 965
rect 110 605 121 949
rect 155 605 166 949
rect 110 565 166 605
rect 196 565 238 965
rect 268 949 358 965
rect 268 605 279 949
rect 347 605 358 949
rect 268 565 358 605
rect 388 565 430 965
rect 460 949 516 965
rect 460 605 471 949
rect 505 605 516 949
rect 460 565 516 605
rect 546 949 599 965
rect 546 606 557 949
rect 591 606 599 949
rect 546 565 599 606
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 165
rect 279 131 347 215
rect 471 131 505 165
rect 557 131 591 215
<< pdiffc >>
rect 35 605 69 949
rect 121 605 155 949
rect 279 605 347 949
rect 471 605 505 949
rect 557 606 591 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 238 965 268 991
rect 358 965 388 991
rect 430 965 460 991
rect 516 965 546 991
rect 80 550 110 565
rect 70 520 110 550
rect 70 308 100 520
rect 166 459 196 565
rect 142 443 196 459
rect 142 409 152 443
rect 186 409 196 443
rect 142 393 196 409
rect 238 534 268 565
rect 238 518 292 534
rect 238 484 248 518
rect 282 484 292 518
rect 238 468 292 484
rect 142 335 196 351
rect 142 308 152 335
rect 70 301 152 308
rect 186 301 196 335
rect 70 278 196 301
rect 80 243 110 278
rect 166 243 196 278
rect 238 243 268 468
rect 358 459 388 565
rect 430 550 460 565
rect 516 550 546 565
rect 430 520 546 550
rect 358 443 472 459
rect 358 429 428 443
rect 418 409 428 429
rect 462 409 472 443
rect 418 393 472 409
rect 516 351 546 520
rect 326 335 380 351
rect 326 301 336 335
rect 370 308 380 335
rect 479 335 546 351
rect 479 308 489 335
rect 370 301 388 308
rect 326 285 388 301
rect 358 243 388 285
rect 430 301 489 308
rect 523 301 546 335
rect 430 278 546 301
rect 430 243 460 278
rect 516 243 546 278
rect 80 89 110 115
rect 166 89 196 115
rect 238 89 268 115
rect 358 89 388 115
rect 430 89 460 115
rect 516 89 546 115
<< polycont >>
rect 152 409 186 443
rect 248 484 282 518
rect 152 301 186 335
rect 428 409 462 443
rect 336 301 370 335
rect 489 301 523 335
<< locali >>
rect 0 1089 638 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 638 1089
rect 35 949 69 965
rect 35 443 69 605
rect 121 949 155 1049
rect 279 949 347 965
rect 121 589 155 605
rect 268 631 279 637
rect 302 597 347 605
rect 279 589 347 597
rect 471 949 505 1049
rect 471 589 505 605
rect 557 949 591 965
rect 557 518 591 606
rect 232 484 248 518
rect 282 484 591 518
rect 35 409 152 443
rect 186 409 370 443
rect 35 215 69 409
rect 152 335 186 351
rect 336 335 370 409
rect 152 261 186 301
rect 268 231 302 301
rect 336 285 370 301
rect 412 409 428 443
rect 462 409 478 443
rect 412 261 446 409
rect 489 335 523 351
rect 489 285 523 301
rect 268 215 347 231
rect 268 197 279 215
rect 35 115 69 131
rect 121 165 155 181
rect 121 61 155 131
rect 557 215 591 484
rect 279 115 347 131
rect 471 165 505 181
rect 471 61 505 131
rect 557 115 591 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 638 61
rect 0 0 638 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 268 605 279 631
rect 279 605 302 631
rect 268 597 302 605
rect 152 227 186 261
rect 268 301 302 335
rect 489 301 523 335
rect 412 227 446 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
<< metal1 >>
rect 0 1089 638 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 638 1089
rect 0 1049 638 1055
rect 256 631 314 637
rect 256 597 268 631
rect 302 597 314 631
rect 256 591 314 597
rect 268 341 302 591
rect 256 335 314 341
rect 477 335 535 341
rect 256 301 268 335
rect 302 301 314 335
rect 455 301 489 335
rect 523 301 535 335
rect 256 295 314 301
rect 477 295 535 301
rect 140 261 198 267
rect 400 261 458 267
rect 140 227 152 261
rect 186 227 412 261
rect 446 227 458 261
rect 140 221 198 227
rect 400 221 458 227
rect 0 55 638 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 638 55
rect 0 0 638 21
<< labels >>
rlabel viali 506 318 506 318 1 B
port 2 n
rlabel metal1 284 375 284 375 1 Y
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
rlabel viali 170 244 170 244 1 A
port 1 n
<< end >>
