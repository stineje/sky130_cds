* File: sky130_osu_sc_18T_hs__and2_1.pxi.spice
* Created: Thu Oct 29 17:05:45 2020
* 
x_PM_SKY130_OSU_SC_18T_HS__AND2_1%GND N_GND_M1003_d N_GND_M1005_b N_GND_c_2_p
+ N_GND_c_8_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_HS__AND2_1%GND
x_PM_SKY130_OSU_SC_18T_HS__AND2_1%VDD N_VDD_M1004_s N_VDD_M1000_d N_VDD_M1004_b
+ N_VDD_c_38_p N_VDD_c_49_p N_VDD_c_39_p N_VDD_c_57_p VDD N_VDD_c_40_p
+ PM_SKY130_OSU_SC_18T_HS__AND2_1%VDD
x_PM_SKY130_OSU_SC_18T_HS__AND2_1%A N_A_M1005_g N_A_M1004_g A N_A_c_69_n
+ N_A_c_70_n PM_SKY130_OSU_SC_18T_HS__AND2_1%A
x_PM_SKY130_OSU_SC_18T_HS__AND2_1%B N_B_M1003_g N_B_M1000_g B N_B_c_104_n
+ N_B_c_105_n PM_SKY130_OSU_SC_18T_HS__AND2_1%B
x_PM_SKY130_OSU_SC_18T_HS__AND2_1%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1004_d N_A_27_115#_M1002_g N_A_27_115#_M1001_g
+ N_A_27_115#_c_142_n N_A_27_115#_c_143_n N_A_27_115#_c_144_n
+ N_A_27_115#_c_145_n N_A_27_115#_c_148_n N_A_27_115#_c_149_n
+ N_A_27_115#_c_158_n N_A_27_115#_c_150_n N_A_27_115#_c_152_n
+ N_A_27_115#_c_153_n N_A_27_115#_c_174_n
+ PM_SKY130_OSU_SC_18T_HS__AND2_1%A_27_115#
x_PM_SKY130_OSU_SC_18T_HS__AND2_1%Y N_Y_M1002_d N_Y_M1001_d Y N_Y_c_209_n
+ N_Y_c_211_n N_Y_c_212_n N_Y_c_213_n PM_SKY130_OSU_SC_18T_HS__AND2_1%Y
cc_1 N_GND_M1005_b N_A_M1005_g 0.0806078f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1005_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1005_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.475 $Y2=1.075
cc_4 N_GND_M1005_b N_A_c_69_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.765
cc_5 N_GND_M1005_b N_A_c_70_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_6 N_GND_M1005_b N_B_M1003_g 0.0460664f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_7 N_GND_c_2_p N_B_M1003_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=1.075
cc_8 N_GND_c_8_p N_B_M1003_g 0.00376152f $X=1.05 $Y=0.825 $X2=0.835 $Y2=1.075
cc_9 N_GND_c_3_p N_B_M1003_g 0.00468827f $X=1.02 $Y=0.17 $X2=0.835 $Y2=1.075
cc_10 N_GND_M1005_b N_B_M1000_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_11 N_GND_M1005_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.96
cc_12 N_GND_M1005_b N_B_c_104_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_13 N_GND_M1005_b N_B_c_105_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_14 N_GND_M1005_b N_A_27_115#_M1002_g 0.0346079f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_15 N_GND_c_8_p N_A_27_115#_M1002_g 0.0103278f $X=1.05 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_16 N_GND_c_3_p N_A_27_115#_M1002_g 0.00468827f $X=1.02 $Y=0.17 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_M1005_b N_A_27_115#_c_142_n 0.0373102f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.1
cc_18 N_GND_M1005_b N_A_27_115#_c_143_n 0.0470206f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.81
cc_19 N_GND_M1005_b N_A_27_115#_c_144_n 0.0076653f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.96
cc_20 N_GND_M1005_b N_A_27_115#_c_145_n 0.0143389f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_21 N_GND_c_2_p N_A_27_115#_c_145_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_22 N_GND_c_3_p N_A_27_115#_c_145_n 0.00476261f $X=1.02 $Y=0.17 $X2=0.26
+ $Y2=0.825
cc_23 N_GND_M1005_b N_A_27_115#_c_148_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.935
cc_24 N_GND_M1005_b N_A_27_115#_c_149_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.935
cc_25 N_GND_M1005_b N_A_27_115#_c_150_n 0.0240789f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_26 N_GND_c_8_p N_A_27_115#_c_150_n 0.00704977f $X=1.05 $Y=0.825 $X2=1.43
+ $Y2=1.935
cc_27 N_GND_M1005_b N_A_27_115#_c_152_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.935
cc_28 N_GND_M1005_b N_A_27_115#_c_153_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.545
cc_29 N_GND_M1005_b Y 0.0401139f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_30 N_GND_M1005_b N_Y_c_209_n 0.0121687f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.48
cc_31 N_GND_c_8_p N_Y_c_209_n 0.00119317f $X=1.05 $Y=0.825 $X2=1.55 $Y2=1.48
cc_32 N_GND_M1005_b N_Y_c_211_n 0.0141689f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_33 N_GND_M1005_b N_Y_c_212_n 0.0163869f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_34 N_GND_M1005_b N_Y_c_213_n 0.00913846f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_35 N_GND_c_8_p N_Y_c_213_n 0.0187614f $X=1.05 $Y=0.825 $X2=1.55 $Y2=0.825
cc_36 N_GND_c_3_p N_Y_c_213_n 0.00476261f $X=1.02 $Y=0.17 $X2=1.55 $Y2=0.825
cc_37 N_VDD_M1004_b N_A_M1004_g 0.0189471f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_38 N_VDD_c_38_p N_A_M1004_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_39 N_VDD_c_39_p N_A_M1004_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=4.585
cc_40 N_VDD_c_40_p N_A_M1004_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.475 $Y2=4.585
cc_41 N_VDD_M1004_s A 0.00742066f $X=0.135 $Y=3.085 $X2=0.275 $Y2=3.33
cc_42 N_VDD_M1004_b A 0.00970321f $X=-0.045 $Y=2.905 $X2=0.275 $Y2=3.33
cc_43 N_VDD_c_38_p A 0.00434783f $X=0.26 $Y=4.135 $X2=0.275 $Y2=3.33
cc_44 N_VDD_M1004_s N_A_c_69_n 0.0127298f $X=0.135 $Y=3.085 $X2=0.27 $Y2=2.765
cc_45 N_VDD_M1004_b N_A_c_69_n 0.00612103f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.765
cc_46 N_VDD_c_38_p N_A_c_69_n 0.00370742f $X=0.26 $Y=4.135 $X2=0.27 $Y2=2.765
cc_47 N_VDD_M1004_b N_A_c_70_n 0.0111025f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=2.765
cc_48 N_VDD_M1004_b N_B_M1000_g 0.0187476f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_49 N_VDD_c_49_p N_B_M1000_g 0.00354579f $X=1.12 $Y=3.795 $X2=0.905 $Y2=4.585
cc_50 N_VDD_c_39_p N_B_M1000_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=4.585
cc_51 N_VDD_c_40_p N_B_M1000_g 0.00468827f $X=1.02 $Y=6.49 $X2=0.905 $Y2=4.585
cc_52 N_VDD_M1004_b B 0.00856863f $X=-0.045 $Y=2.905 $X2=0.955 $Y2=2.96
cc_53 N_VDD_c_49_p B 0.00240671f $X=1.12 $Y=3.795 $X2=0.955 $Y2=2.96
cc_54 N_VDD_M1004_b N_B_c_104_n 0.00170274f $X=-0.045 $Y=2.905 $X2=0.95
+ $Y2=2.425
cc_55 N_VDD_M1004_b N_A_27_115#_c_144_n 0.0267233f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.96
cc_56 N_VDD_c_49_p N_A_27_115#_c_144_n 0.00354579f $X=1.12 $Y=3.795 $X2=1.352
+ $Y2=2.96
cc_57 N_VDD_c_57_p N_A_27_115#_c_144_n 0.00606474f $X=1.12 $Y=6.507 $X2=1.352
+ $Y2=2.96
cc_58 N_VDD_c_40_p N_A_27_115#_c_144_n 0.00468827f $X=1.02 $Y=6.49 $X2=1.352
+ $Y2=2.96
cc_59 N_VDD_M1004_b N_A_27_115#_c_158_n 0.00155118f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=3.795
cc_60 N_VDD_c_39_p N_A_27_115#_c_158_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69
+ $Y2=3.795
cc_61 N_VDD_c_40_p N_A_27_115#_c_158_n 0.00475776f $X=1.02 $Y=6.49 $X2=0.69
+ $Y2=3.795
cc_62 N_VDD_M1004_b N_A_27_115#_c_153_n 8.22047e-19 $X=-0.045 $Y=2.905 $X2=0.65
+ $Y2=3.545
cc_63 N_VDD_M1004_b N_Y_c_212_n 0.0100094f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.59
cc_64 N_VDD_c_57_p N_Y_c_212_n 0.00757793f $X=1.12 $Y=6.507 $X2=1.55 $Y2=2.59
cc_65 N_VDD_c_40_p N_Y_c_212_n 0.00476261f $X=1.02 $Y=6.49 $X2=1.55 $Y2=2.59
cc_66 N_A_M1005_g N_B_M1003_g 0.129148f $X=0.475 $Y=1.075 $X2=0.835 $Y2=1.075
cc_67 N_A_M1005_g N_B_M1000_g 0.0498038f $X=0.475 $Y=1.075 $X2=0.905 $Y2=4.585
cc_68 N_A_M1005_g N_B_c_104_n 7.8234e-19 $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.425
cc_69 N_A_M1005_g N_A_27_115#_c_145_n 0.0158058f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_70 N_A_M1005_g N_A_27_115#_c_148_n 0.0160984f $X=0.475 $Y=1.075 $X2=0.525
+ $Y2=1.935
cc_71 N_A_c_69_n N_A_27_115#_c_148_n 2.65873e-19 $X=0.27 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_72 N_A_c_70_n N_A_27_115#_c_148_n 0.00117122f $X=0.475 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_73 N_A_c_69_n N_A_27_115#_c_149_n 0.0055861f $X=0.27 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_74 N_A_c_70_n N_A_27_115#_c_149_n 0.00133457f $X=0.475 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_75 N_A_M1005_g N_A_27_115#_c_152_n 0.00322084f $X=0.475 $Y=1.075 $X2=0.61
+ $Y2=1.935
cc_76 N_A_M1005_g N_A_27_115#_c_153_n 0.0265302f $X=0.475 $Y=1.075 $X2=0.65
+ $Y2=3.545
cc_77 N_A_M1004_g N_A_27_115#_c_153_n 0.0140172f $X=0.475 $Y=4.585 $X2=0.65
+ $Y2=3.545
cc_78 A N_A_27_115#_c_153_n 0.00758489f $X=0.275 $Y=3.33 $X2=0.65 $Y2=3.545
cc_79 N_A_c_69_n N_A_27_115#_c_153_n 0.0456533f $X=0.27 $Y=2.765 $X2=0.65
+ $Y2=3.545
cc_80 N_A_c_70_n N_A_27_115#_c_153_n 0.00766302f $X=0.475 $Y=2.765 $X2=0.65
+ $Y2=3.545
cc_81 N_A_M1004_g N_A_27_115#_c_174_n 0.00884152f $X=0.475 $Y=4.585 $X2=0.65
+ $Y2=3.715
cc_82 N_B_M1003_g N_A_27_115#_M1002_g 0.0347278f $X=0.835 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_83 N_B_M1003_g N_A_27_115#_c_142_n 0.0104742f $X=0.835 $Y=1.075 $X2=1.37
+ $Y2=2.1
cc_84 N_B_M1000_g N_A_27_115#_c_143_n 0.00773101f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.81
cc_85 N_B_c_104_n N_A_27_115#_c_143_n 0.0033451f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.81
cc_86 N_B_c_105_n N_A_27_115#_c_143_n 0.0206104f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.81
cc_87 N_B_M1000_g N_A_27_115#_c_144_n 0.0395234f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.96
cc_88 B N_A_27_115#_c_144_n 0.0037561f $X=0.955 $Y=2.96 $X2=1.352 $Y2=2.96
cc_89 N_B_c_104_n N_A_27_115#_c_144_n 0.00156524f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.96
cc_90 N_B_M1003_g N_A_27_115#_c_150_n 0.0182215f $X=0.835 $Y=1.075 $X2=1.43
+ $Y2=1.935
cc_91 N_B_c_104_n N_A_27_115#_c_150_n 0.0101796f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_92 N_B_c_105_n N_A_27_115#_c_150_n 0.00258465f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_93 N_B_M1003_g N_A_27_115#_c_153_n 0.00755919f $X=0.835 $Y=1.075 $X2=0.65
+ $Y2=3.545
cc_94 N_B_M1000_g N_A_27_115#_c_153_n 0.0133197f $X=0.905 $Y=4.585 $X2=0.65
+ $Y2=3.545
cc_95 B N_A_27_115#_c_153_n 0.00866797f $X=0.955 $Y=2.96 $X2=0.65 $Y2=3.545
cc_96 N_B_c_104_n N_A_27_115#_c_153_n 0.0541375f $X=0.95 $Y=2.425 $X2=0.65
+ $Y2=3.545
cc_97 B N_A_27_115#_c_174_n 0.00286715f $X=0.955 $Y=2.96 $X2=0.65 $Y2=3.715
cc_98 N_B_M1003_g Y 6.71108e-19 $X=0.835 $Y=1.075 $X2=1.555 $Y2=2.22
cc_99 N_B_c_104_n Y 0.00695761f $X=0.95 $Y=2.425 $X2=1.555 $Y2=2.22
cc_100 N_B_M1003_g N_Y_c_209_n 7.96664e-19 $X=0.835 $Y=1.075 $X2=1.55 $Y2=1.48
cc_101 N_B_c_104_n N_Y_c_211_n 0.00532157f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_102 N_B_c_105_n N_Y_c_211_n 5.70769e-19 $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_103 B N_Y_c_212_n 0.00659455f $X=0.955 $Y=2.96 $X2=1.55 $Y2=2.59
cc_104 N_B_c_104_n N_Y_c_212_n 0.0153635f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_105 N_A_27_115#_M1002_g Y 0.00406656f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_106 N_A_27_115#_c_142_n Y 0.00711756f $X=1.37 $Y=2.1 $X2=1.555 $Y2=2.22
cc_107 N_A_27_115#_c_143_n Y 0.00892438f $X=1.352 $Y=2.81 $X2=1.555 $Y2=2.22
cc_108 N_A_27_115#_c_150_n Y 0.0152626f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_109 N_A_27_115#_M1002_g N_Y_c_209_n 0.00681195f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.48
cc_110 N_A_27_115#_c_142_n N_Y_c_209_n 0.00154864f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=1.48
cc_111 N_A_27_115#_c_150_n N_Y_c_209_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.48
cc_112 N_A_27_115#_c_142_n N_Y_c_211_n 4.58687e-19 $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_113 N_A_27_115#_c_143_n N_Y_c_211_n 0.00721849f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_114 N_A_27_115#_c_150_n N_Y_c_211_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_115 N_A_27_115#_c_142_n N_Y_c_212_n 0.00125776f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_116 N_A_27_115#_c_143_n N_Y_c_212_n 0.0115869f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_117 N_A_27_115#_c_144_n N_Y_c_212_n 0.00807887f $X=1.352 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_118 N_A_27_115#_c_150_n N_Y_c_212_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_119 N_A_27_115#_M1002_g N_Y_c_213_n 0.00580462f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_120 N_A_27_115#_c_142_n N_Y_c_213_n 0.00168f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=0.825
cc_121 N_A_27_115#_c_150_n N_Y_c_213_n 0.00510008f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
