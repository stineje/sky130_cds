* File: sky130_osu_sc_15T_ms__ant.spice
* Created: Fri Nov 12 14:40:57 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ms__ant.pex.spice"
.subckt sky130_osu_sc_15T_ms__ant  GND VDD A
* 
* A	A
* VDD	VDD
* GND	GND
MM1000 N_A_M1000_s N_A_M1000_g N_A_M1000_s N_GND_M1000_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_M1001_s N_VDD_M1001_b PSHORT L=0.15 W=2
+ AD=0.53 AS=0.53 PD=4.53 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.2
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX2_noxref N_GND_M1000_b N_VDD_M1001_b NWDIODE A=3.068 P=7.98
pX3_noxref noxref_4 A A PROBETYPE=1
*
.include "sky130_osu_sc_15T_ms__ant.pxi.spice"
*
.ends
*
*
