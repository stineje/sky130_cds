magic
tech sky130A
magscale 1 2
timestamp 1598479240
<< checkpaint >>
rect -1260 -1260 1261 1261
<< nwell >>
rect -9 581 728 1341
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
rect 338 617 368 1217
rect 424 617 454 1217
rect 510 617 540 1217
rect 596 617 626 1217
<< nmoslvt >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
rect 338 115 368 315
rect 424 115 454 315
rect 510 115 540 315
rect 596 115 626 315
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 166 315
rect 110 131 121 267
rect 155 131 166 267
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 267 338 315
rect 282 131 293 267
rect 327 131 338 267
rect 282 115 338 131
rect 368 267 424 315
rect 368 131 379 267
rect 413 131 424 267
rect 368 115 424 131
rect 454 267 510 315
rect 454 131 465 267
rect 499 131 510 267
rect 454 115 510 131
rect 540 267 596 315
rect 540 131 551 267
rect 585 131 596 267
rect 540 115 596 131
rect 626 267 679 315
rect 626 131 637 267
rect 671 131 679 267
rect 626 115 679 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 657 35 1201
rect 69 657 80 1201
rect 27 617 80 657
rect 110 1201 166 1217
rect 110 793 121 1201
rect 155 793 166 1201
rect 110 617 166 793
rect 196 1201 252 1217
rect 196 657 207 1201
rect 241 657 252 1201
rect 196 617 252 657
rect 282 1201 338 1217
rect 282 657 293 1201
rect 327 657 338 1201
rect 282 617 338 657
rect 368 1201 424 1217
rect 368 657 379 1201
rect 413 657 424 1201
rect 368 617 424 657
rect 454 1201 510 1217
rect 454 657 465 1201
rect 499 657 510 1201
rect 454 617 510 657
rect 540 1201 596 1217
rect 540 657 551 1201
rect 585 657 596 1201
rect 540 617 596 657
rect 626 1201 679 1217
rect 626 657 637 1201
rect 671 657 679 1201
rect 626 617 679 657
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 207 131 241 267
rect 293 131 327 267
rect 379 131 413 267
rect 465 131 499 267
rect 551 131 585 267
rect 637 131 671 267
<< pdiffc >>
rect 35 657 69 1201
rect 121 793 155 1201
rect 207 657 241 1201
rect 293 657 327 1201
rect 379 657 413 1201
rect 465 657 499 1201
rect 551 657 585 1201
rect 637 657 671 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1244
rect 338 1217 368 1243
rect 424 1217 454 1243
rect 510 1217 540 1243
rect 596 1217 626 1243
rect 80 529 110 617
rect 166 602 196 617
rect 252 602 282 617
rect 338 602 368 617
rect 424 602 454 617
rect 510 602 540 617
rect 596 602 626 617
rect 166 572 626 602
rect 80 513 154 529
rect 80 479 110 513
rect 144 479 154 513
rect 80 463 154 479
rect 80 315 110 463
rect 221 420 251 572
rect 166 404 251 420
rect 166 370 176 404
rect 210 384 251 404
rect 510 384 540 572
rect 210 370 626 384
rect 166 354 626 370
rect 166 315 196 354
rect 252 315 282 354
rect 338 315 368 354
rect 424 315 454 354
rect 510 315 540 354
rect 596 315 626 354
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
rect 338 89 368 115
rect 424 89 454 115
rect 510 89 540 115
rect 596 89 626 115
<< polycont >>
rect 110 479 144 513
rect 176 370 210 404
<< locali >>
rect 0 1305 726 1332
rect 0 1271 51 1305
rect 85 1271 187 1305
rect 221 1271 323 1305
rect 357 1271 459 1305
rect 493 1271 595 1305
rect 629 1271 726 1305
rect 35 1201 69 1217
rect 121 1201 155 1271
rect 121 777 155 793
rect 207 1201 241 1217
rect 35 404 69 657
rect 110 513 144 649
rect 207 609 241 657
rect 293 1201 327 1271
rect 293 641 327 657
rect 379 1201 413 1217
rect 379 609 413 657
rect 465 1201 499 1271
rect 465 641 499 657
rect 551 1201 585 1217
rect 551 609 585 657
rect 637 1201 671 1271
rect 637 641 671 657
rect 110 463 144 479
rect 176 404 210 420
rect 35 370 176 404
rect 35 267 69 370
rect 176 354 210 370
rect 35 115 69 131
rect 121 267 155 283
rect 121 61 155 131
rect 207 267 241 279
rect 207 115 241 131
rect 293 267 327 283
rect 293 61 327 131
rect 379 267 413 279
rect 379 115 413 131
rect 465 267 499 283
rect 465 61 499 131
rect 551 267 585 279
rect 551 115 585 131
rect 637 267 671 283
rect 637 61 671 131
rect 0 27 51 61
rect 85 27 187 61
rect 221 27 323 61
rect 357 27 459 61
rect 493 27 595 61
rect 629 27 726 61
rect 0 0 726 27
<< viali >>
rect 110 649 144 683
rect 207 575 241 609
rect 379 575 413 609
rect 551 575 585 609
rect 207 279 241 313
rect 379 279 413 313
rect 551 279 585 313
<< metal1 >>
rect 0 1271 726 1332
rect 98 683 156 689
rect 64 649 110 683
rect 144 649 156 683
rect 98 643 156 649
rect 195 609 253 615
rect 367 609 425 615
rect 539 609 597 615
rect 195 575 207 609
rect 241 575 379 609
rect 413 575 551 609
rect 585 575 597 609
rect 195 569 253 575
rect 367 569 425 575
rect 539 569 597 575
rect 207 319 241 569
rect 379 319 413 569
rect 551 319 585 569
rect 195 313 253 319
rect 367 313 425 319
rect 539 313 597 319
rect 195 279 207 313
rect 241 279 379 313
rect 413 279 551 313
rect 585 279 597 313
rect 195 273 253 279
rect 367 273 425 279
rect 539 273 597 279
rect 0 0 726 61
<< labels >>
rlabel metal1 127 666 127 666 1 A
port 1 n
rlabel metal1 211 454 211 454 1 Y
port 2 n
rlabel metal1 68 44 68 44 1 gnd
rlabel metal1 68 1288 68 1288 1 vdd
<< end >>
