* File: sky130_osu_sc_18T_ms__nand2_l.pxi.spice
* Created: Fri Nov 12 14:05:20 2021
* 
x_PM_SKY130_OSU_SC_18T_MS__NAND2_L%GND N_GND_M1000_d N_GND_M1001_b N_GND_c_2_p
+ N_GND_c_9_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_MS__NAND2_L%GND
x_PM_SKY130_OSU_SC_18T_MS__NAND2_L%VDD N_VDD_M1003_s N_VDD_M1002_d N_VDD_M1003_b
+ N_VDD_c_26_p N_VDD_c_27_p N_VDD_c_33_p VDD N_VDD_c_28_p
+ PM_SKY130_OSU_SC_18T_MS__NAND2_L%VDD
x_PM_SKY130_OSU_SC_18T_MS__NAND2_L%A N_A_M1001_g N_A_M1003_g N_A_c_44_n
+ N_A_c_45_n A PM_SKY130_OSU_SC_18T_MS__NAND2_L%A
x_PM_SKY130_OSU_SC_18T_MS__NAND2_L%B N_B_M1000_g N_B_M1002_g N_B_c_72_n
+ N_B_c_74_n N_B_c_75_n B PM_SKY130_OSU_SC_18T_MS__NAND2_L%B
x_PM_SKY130_OSU_SC_18T_MS__NAND2_L%Y N_Y_M1001_s N_Y_M1003_d N_Y_c_102_n
+ N_Y_c_105_n N_Y_c_106_n N_Y_c_107_n Y N_Y_c_109_n
+ PM_SKY130_OSU_SC_18T_MS__NAND2_L%Y
cc_1 N_GND_M1001_b N_A_M1001_g 0.105321f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.945
cc_3 N_GND_c_3_p N_A_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1001_b N_A_M1003_g 0.00342256f $X=-0.045 $Y=0 $X2=0.475 $Y2=5.085
cc_5 N_GND_M1001_b N_A_c_44_n 0.0490341f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.685
cc_6 N_GND_M1001_b N_A_c_45_n 0.00856875f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.685
cc_7 N_GND_M1001_b N_B_M1000_g 0.044779f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.945
cc_8 N_GND_c_2_p N_B_M1000_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.945
cc_9 N_GND_c_9_p N_B_M1000_g 0.00713292f $X=1.05 $Y=0.825 $X2=0.835 $Y2=0.945
cc_10 N_GND_c_3_p N_B_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.945
cc_11 N_GND_M1001_b N_B_M1002_g 0.0497877f $X=-0.045 $Y=0 $X2=0.905 $Y2=5.085
cc_12 N_GND_M1001_b N_B_c_72_n 0.0355341f $X=-0.045 $Y=0 $X2=0.915 $Y2=1.935
cc_13 N_GND_c_9_p N_B_c_72_n 0.00219428f $X=1.05 $Y=0.825 $X2=0.915 $Y2=1.935
cc_14 N_GND_M1001_b N_B_c_74_n 0.0293783f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.96
cc_15 N_GND_M1001_b N_B_c_75_n 0.0123076f $X=-0.045 $Y=0 $X2=1.06 $Y2=1.935
cc_16 N_GND_M1001_b B 0.00499588f $X=-0.045 $Y=0 $X2=1.06 $Y2=2.96
cc_17 N_GND_M1001_b N_Y_c_102_n 0.0125734f $X=-0.045 $Y=0 $X2=0.26 $Y2=0.825
cc_18 N_GND_c_2_p N_Y_c_102_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26 $Y2=0.825
cc_19 N_GND_c_3_p N_Y_c_102_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26 $Y2=0.825
cc_20 N_GND_M1001_b N_Y_c_105_n 0.00860362f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.59
cc_21 N_GND_M1001_b N_Y_c_106_n 0.0101912f $X=-0.045 $Y=0 $X2=0.605 $Y2=1.48
cc_22 N_GND_M1001_b N_Y_c_107_n 0.0242516f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.48
cc_23 N_GND_M1001_b Y 0.0166407f $X=-0.045 $Y=0 $X2=0.68 $Y2=2.35
cc_24 N_GND_M1001_b N_Y_c_109_n 0.00535447f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.59
cc_25 N_VDD_M1003_b N_A_M1003_g 0.0970858f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=5.085
cc_26 N_VDD_c_26_p N_A_M1003_g 0.00713292f $X=0.26 $Y=4.815 $X2=0.475 $Y2=5.085
cc_27 N_VDD_c_27_p N_A_M1003_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=5.085
cc_28 N_VDD_c_28_p N_A_M1003_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=5.085
cc_29 N_VDD_M1003_b N_A_c_45_n 0.0153337f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=2.685
cc_30 N_VDD_M1003_b A 0.0208751f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=3.33
cc_31 N_VDD_M1003_b N_B_M1002_g 0.104061f $X=-0.045 $Y=2.905 $X2=0.905 $Y2=5.085
cc_32 N_VDD_c_27_p N_B_M1002_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=5.085
cc_33 N_VDD_c_33_p N_B_M1002_g 0.00713292f $X=1.12 $Y=4.815 $X2=0.905 $Y2=5.085
cc_34 N_VDD_c_28_p N_B_M1002_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.905 $Y2=5.085
cc_35 N_VDD_M1003_b N_B_c_74_n 0.00391589f $X=-0.045 $Y=2.905 $X2=1.06 $Y2=2.96
cc_36 N_VDD_M1003_b B 0.0168801f $X=-0.045 $Y=2.905 $X2=1.06 $Y2=2.96
cc_37 N_VDD_M1003_b N_Y_c_105_n 0.027504f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.59
cc_38 N_VDD_c_27_p N_Y_c_105_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69 $Y2=2.59
cc_39 N_VDD_c_28_p N_Y_c_105_n 0.00475776f $X=1.02 $Y=6.47 $X2=0.69 $Y2=2.59
cc_40 N_A_M1001_g N_B_M1000_g 0.102948f $X=0.475 $Y=0.945 $X2=0.835 $Y2=0.945
cc_41 N_A_M1001_g N_B_M1002_g 0.105181f $X=0.475 $Y=0.945 $X2=0.905 $Y2=5.085
cc_42 N_A_M1001_g N_B_c_74_n 0.00248145f $X=0.475 $Y=0.945 $X2=1.06 $Y2=2.96
cc_43 N_A_M1001_g N_B_c_75_n 0.00282768f $X=0.475 $Y=0.945 $X2=1.06 $Y2=1.935
cc_44 N_A_M1001_g N_Y_c_102_n 0.0152627f $X=0.475 $Y=0.945 $X2=0.26 $Y2=0.825
cc_45 N_A_M1001_g N_Y_c_105_n 0.0253166f $X=0.475 $Y=0.945 $X2=0.69 $Y2=2.59
cc_46 N_A_c_45_n N_Y_c_105_n 0.0513069f $X=0.32 $Y=2.685 $X2=0.69 $Y2=2.59
cc_47 A N_Y_c_105_n 0.00831114f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.59
cc_48 N_A_M1001_g N_Y_c_106_n 0.0136921f $X=0.475 $Y=0.945 $X2=0.605 $Y2=1.48
cc_49 N_A_M1001_g N_Y_c_107_n 0.00393078f $X=0.475 $Y=0.945 $X2=0.405 $Y2=1.48
cc_50 N_A_M1001_g Y 0.0125133f $X=0.475 $Y=0.945 $X2=0.68 $Y2=2.35
cc_51 N_A_M1001_g N_Y_c_109_n 0.00216533f $X=0.475 $Y=0.945 $X2=0.69 $Y2=2.59
cc_52 N_A_c_44_n N_Y_c_109_n 0.00278592f $X=0.32 $Y=2.685 $X2=0.69 $Y2=2.59
cc_53 N_A_c_45_n N_Y_c_109_n 0.00474021f $X=0.32 $Y=2.685 $X2=0.69 $Y2=2.59
cc_54 A N_Y_c_109_n 0.00152954f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.59
cc_55 N_B_M1002_g N_Y_c_105_n 0.0309814f $X=0.905 $Y=5.085 $X2=0.69 $Y2=2.59
cc_56 N_B_c_74_n N_Y_c_105_n 0.0295869f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_57 N_B_c_75_n N_Y_c_105_n 5.24123e-19 $X=1.06 $Y=1.935 $X2=0.69 $Y2=2.59
cc_58 B N_Y_c_105_n 0.00831114f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_59 N_B_M1000_g N_Y_c_106_n 0.00853825f $X=0.835 $Y=0.945 $X2=0.605 $Y2=1.48
cc_60 N_B_M1000_g Y 0.00770103f $X=0.835 $Y=0.945 $X2=0.68 $Y2=2.35
cc_61 N_B_M1002_g Y 0.00539744f $X=0.905 $Y=5.085 $X2=0.68 $Y2=2.35
cc_62 N_B_c_72_n Y 0.00401356f $X=0.915 $Y=1.935 $X2=0.68 $Y2=2.35
cc_63 N_B_c_74_n Y 0.0183986f $X=1.06 $Y=2.96 $X2=0.68 $Y2=2.35
cc_64 N_B_c_75_n Y 0.0141623f $X=1.06 $Y=1.935 $X2=0.68 $Y2=2.35
cc_65 N_B_M1002_g N_Y_c_109_n 0.00341272f $X=0.905 $Y=5.085 $X2=0.69 $Y2=2.59
cc_66 N_B_c_72_n N_Y_c_109_n 0.00144278f $X=0.915 $Y=1.935 $X2=0.69 $Y2=2.59
cc_67 N_B_c_74_n N_Y_c_109_n 0.00640429f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
cc_68 N_B_c_75_n N_Y_c_109_n 0.00194461f $X=1.06 $Y=1.935 $X2=0.69 $Y2=2.59
cc_69 B N_Y_c_109_n 0.00280435f $X=1.06 $Y=2.96 $X2=0.69 $Y2=2.59
