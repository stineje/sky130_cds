* File: sky130_osu_sc_12T_ms__and2_l.pxi.spice
* Created: Fri Nov 12 15:20:51 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__AND2_L%GND N_GND_M1001_d N_GND_M1003_b N_GND_c_2_p
+ N_GND_c_9_p GND N_GND_c_3_p PM_SKY130_OSU_SC_12T_MS__AND2_L%GND
x_PM_SKY130_OSU_SC_12T_MS__AND2_L%VDD N_VDD_M1002_s N_VDD_M1004_d N_VDD_M1002_b
+ N_VDD_c_36_p N_VDD_c_37_p N_VDD_c_46_p N_VDD_c_52_p VDD N_VDD_c_38_p
+ PM_SKY130_OSU_SC_12T_MS__AND2_L%VDD
x_PM_SKY130_OSU_SC_12T_MS__AND2_L%A N_A_M1003_g N_A_M1002_g N_A_c_66_n
+ N_A_c_67_n A PM_SKY130_OSU_SC_12T_MS__AND2_L%A
x_PM_SKY130_OSU_SC_12T_MS__AND2_L%B N_B_M1001_g N_B_M1004_g N_B_c_101_n
+ N_B_c_102_n B PM_SKY130_OSU_SC_12T_MS__AND2_L%B
x_PM_SKY130_OSU_SC_12T_MS__AND2_L%A_27_115# N_A_27_115#_M1003_s
+ N_A_27_115#_M1002_d N_A_27_115#_M1000_g N_A_27_115#_M1005_g
+ N_A_27_115#_c_140_n N_A_27_115#_c_141_n N_A_27_115#_c_142_n
+ N_A_27_115#_c_143_n N_A_27_115#_c_146_n N_A_27_115#_c_147_n
+ N_A_27_115#_c_156_n N_A_27_115#_c_148_n N_A_27_115#_c_149_n
+ N_A_27_115#_c_150_n N_A_27_115#_c_160_n
+ PM_SKY130_OSU_SC_12T_MS__AND2_L%A_27_115#
x_PM_SKY130_OSU_SC_12T_MS__AND2_L%Y N_Y_M1000_d N_Y_M1005_d N_Y_c_208_n
+ N_Y_c_210_n Y N_Y_c_212_n N_Y_c_213_n PM_SKY130_OSU_SC_12T_MS__AND2_L%Y
cc_1 N_GND_M1003_b N_A_M1003_g 0.109036f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.755
cc_2 N_GND_c_2_p N_A_M1003_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.755
cc_3 N_GND_c_3_p N_A_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.755
cc_4 N_GND_M1003_b N_A_c_66_n 0.0391443f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.66
cc_5 N_GND_M1003_b N_A_c_67_n 0.00303836f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.48
cc_6 N_GND_M1003_b A 0.013676f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.485
cc_7 N_GND_M1003_b N_B_M1001_g 0.0744418f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.755
cc_8 N_GND_c_2_p N_B_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.755
cc_9 N_GND_c_9_p N_B_M1001_g 0.00319969f $X=1.05 $Y=0.74 $X2=0.835 $Y2=0.755
cc_10 N_GND_c_3_p N_B_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.835 $Y2=0.755
cc_11 N_GND_M1003_b N_B_M1004_g 0.0160032f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.445
cc_12 N_GND_M1003_b N_B_c_101_n 0.0331543f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.31
cc_13 N_GND_M1003_b N_B_c_102_n 0.00275487f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.31
cc_14 N_GND_M1003_b B 0.0078879f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.48
cc_15 N_GND_M1003_b N_A_27_115#_M1000_g 0.0635173f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.755
cc_16 N_GND_c_9_p N_A_27_115#_M1000_g 0.00584472f $X=1.05 $Y=0.74 $X2=1.335
+ $Y2=0.755
cc_17 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=0.755
cc_18 N_GND_M1003_b N_A_27_115#_c_140_n 0.0433374f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=1.99
cc_19 N_GND_M1003_b N_A_27_115#_c_141_n 0.0470152f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.7
cc_20 N_GND_M1003_b N_A_27_115#_c_142_n 0.0076832f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.85
cc_21 N_GND_M1003_b N_A_27_115#_c_143_n 0.0371775f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_22 N_GND_c_2_p N_A_27_115#_c_143_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_23 N_GND_c_3_p N_A_27_115#_c_143_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_24 N_GND_M1003_b N_A_27_115#_c_146_n 0.0022584f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.755
cc_25 N_GND_M1003_b N_A_27_115#_c_147_n 0.00906593f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.755
cc_26 N_GND_M1003_b N_A_27_115#_c_148_n 0.0252109f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.755
cc_27 N_GND_M1003_b N_A_27_115#_c_149_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.755
cc_28 N_GND_M1003_b N_A_27_115#_c_150_n 0.00693462f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.025
cc_29 N_GND_M1003_b N_Y_c_208_n 0.03243f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.74
cc_30 N_GND_c_3_p N_Y_c_208_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.74
cc_31 N_GND_M1003_b N_Y_c_210_n 0.0169214f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.48
cc_32 N_GND_M1003_b Y 0.0380962f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.11
cc_33 N_GND_M1003_b N_Y_c_212_n 0.0156693f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.37
cc_34 N_GND_M1003_b N_Y_c_213_n 0.0141861f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.48
cc_35 N_VDD_M1002_b N_A_M1002_g 0.0263651f $X=-0.045 $Y=2.795 $X2=0.475
+ $Y2=3.445
cc_36 N_VDD_c_36_p N_A_M1002_g 0.00713292f $X=0.26 $Y=3.275 $X2=0.475 $Y2=3.445
cc_37 N_VDD_c_37_p N_A_M1002_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.445
cc_38 N_VDD_c_38_p N_A_M1002_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.445
cc_39 N_VDD_M1002_b N_A_c_66_n 0.0127774f $X=-0.045 $Y=2.795 $X2=0.475 $Y2=2.66
cc_40 N_VDD_c_36_p N_A_c_66_n 0.00165206f $X=0.26 $Y=3.275 $X2=0.475 $Y2=2.66
cc_41 N_VDD_M1002_b N_A_c_67_n 0.00194065f $X=-0.045 $Y=2.795 $X2=0.27 $Y2=2.48
cc_42 N_VDD_c_36_p N_A_c_67_n 0.0109365f $X=0.26 $Y=3.275 $X2=0.27 $Y2=2.48
cc_43 N_VDD_c_36_p A 0.00121903f $X=0.26 $Y=3.275 $X2=0.27 $Y2=2.485
cc_44 N_VDD_M1002_b N_B_M1004_g 0.023266f $X=-0.045 $Y=2.795 $X2=0.905 $Y2=3.445
cc_45 N_VDD_c_37_p N_B_M1004_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.445
cc_46 N_VDD_c_46_p N_B_M1004_g 0.00354579f $X=1.12 $Y=3.275 $X2=0.905 $Y2=3.445
cc_47 N_VDD_c_38_p N_B_M1004_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.905 $Y2=3.445
cc_48 N_VDD_c_46_p N_B_c_101_n 0.00116158f $X=1.12 $Y=3.275 $X2=0.95 $Y2=2.31
cc_49 N_VDD_c_46_p B 0.00688801f $X=1.12 $Y=3.275 $X2=0.95 $Y2=2.48
cc_50 N_VDD_M1002_b N_A_27_115#_M1005_g 0.0243035f $X=-0.045 $Y=2.795 $X2=1.335
+ $Y2=3.445
cc_51 N_VDD_c_46_p N_A_27_115#_M1005_g 0.00354579f $X=1.12 $Y=3.275 $X2=1.335
+ $Y2=3.445
cc_52 N_VDD_c_52_p N_A_27_115#_M1005_g 0.00606474f $X=1.12 $Y=4.287 $X2=1.335
+ $Y2=3.445
cc_53 N_VDD_c_38_p N_A_27_115#_M1005_g 0.00468827f $X=1.02 $Y=4.25 $X2=1.335
+ $Y2=3.445
cc_54 N_VDD_M1002_b N_A_27_115#_c_142_n 0.0052627f $X=-0.045 $Y=2.795 $X2=1.352
+ $Y2=2.85
cc_55 N_VDD_M1002_b N_A_27_115#_c_156_n 0.00155118f $X=-0.045 $Y=2.795 $X2=0.69
+ $Y2=3.275
cc_56 N_VDD_c_37_p N_A_27_115#_c_156_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69
+ $Y2=3.275
cc_57 N_VDD_c_38_p N_A_27_115#_c_156_n 0.00475776f $X=1.02 $Y=4.25 $X2=0.69
+ $Y2=3.275
cc_58 N_VDD_M1002_b N_A_27_115#_c_150_n 0.00215047f $X=-0.045 $Y=2.795 $X2=0.65
+ $Y2=3.025
cc_59 N_VDD_M1002_b N_A_27_115#_c_160_n 0.0028529f $X=-0.045 $Y=2.795 $X2=0.65
+ $Y2=3.195
cc_60 N_VDD_M1002_b N_Y_c_210_n 0.0129676f $X=-0.045 $Y=2.795 $X2=1.55 $Y2=2.48
cc_61 N_VDD_c_52_p N_Y_c_210_n 0.00757793f $X=1.12 $Y=4.287 $X2=1.55 $Y2=2.48
cc_62 N_VDD_c_38_p N_Y_c_210_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.55 $Y2=2.48
cc_63 N_A_M1003_g N_B_M1001_g 0.124037f $X=0.475 $Y=0.755 $X2=0.835 $Y2=0.755
cc_64 N_A_M1003_g N_B_M1004_g 0.0324123f $X=0.475 $Y=0.755 $X2=0.905 $Y2=3.445
cc_65 N_A_M1003_g N_B_c_102_n 4.36797e-19 $X=0.475 $Y=0.755 $X2=0.95 $Y2=2.31
cc_66 A B 0.0168274f $X=0.27 $Y=2.485 $X2=0.95 $Y2=2.48
cc_67 N_A_M1003_g N_A_27_115#_c_143_n 0.0284873f $X=0.475 $Y=0.755 $X2=0.26
+ $Y2=0.74
cc_68 N_A_M1003_g N_A_27_115#_c_146_n 0.0133945f $X=0.475 $Y=0.755 $X2=0.525
+ $Y2=1.755
cc_69 N_A_c_66_n N_A_27_115#_c_146_n 8.11165e-19 $X=0.475 $Y=2.66 $X2=0.525
+ $Y2=1.755
cc_70 A N_A_27_115#_c_146_n 0.00481725f $X=0.27 $Y=2.485 $X2=0.525 $Y2=1.755
cc_71 N_A_c_66_n N_A_27_115#_c_147_n 0.00111032f $X=0.475 $Y=2.66 $X2=0.345
+ $Y2=1.755
cc_72 N_A_c_67_n N_A_27_115#_c_147_n 0.00345248f $X=0.27 $Y=2.48 $X2=0.345
+ $Y2=1.755
cc_73 A N_A_27_115#_c_147_n 0.00417148f $X=0.27 $Y=2.485 $X2=0.345 $Y2=1.755
cc_74 N_A_M1003_g N_A_27_115#_c_149_n 0.00322084f $X=0.475 $Y=0.755 $X2=0.61
+ $Y2=1.755
cc_75 N_A_M1003_g N_A_27_115#_c_150_n 0.0262426f $X=0.475 $Y=0.755 $X2=0.65
+ $Y2=3.025
cc_76 N_A_M1002_g N_A_27_115#_c_150_n 0.00943195f $X=0.475 $Y=3.445 $X2=0.65
+ $Y2=3.025
cc_77 N_A_c_66_n N_A_27_115#_c_150_n 0.00759169f $X=0.475 $Y=2.66 $X2=0.65
+ $Y2=3.025
cc_78 N_A_c_67_n N_A_27_115#_c_150_n 0.0275984f $X=0.27 $Y=2.48 $X2=0.65
+ $Y2=3.025
cc_79 A N_A_27_115#_c_150_n 0.00281638f $X=0.27 $Y=2.485 $X2=0.65 $Y2=3.025
cc_80 N_A_M1002_g N_A_27_115#_c_160_n 0.00355211f $X=0.475 $Y=3.445 $X2=0.65
+ $Y2=3.195
cc_81 N_B_M1001_g N_A_27_115#_M1000_g 0.0383396f $X=0.835 $Y=0.755 $X2=1.335
+ $Y2=0.755
cc_82 N_B_M1001_g N_A_27_115#_c_140_n 0.0125873f $X=0.835 $Y=0.755 $X2=1.37
+ $Y2=1.99
cc_83 N_B_M1004_g N_A_27_115#_c_141_n 0.00806858f $X=0.905 $Y=3.445 $X2=1.352
+ $Y2=2.7
cc_84 N_B_c_101_n N_A_27_115#_c_141_n 0.0211828f $X=0.95 $Y=2.31 $X2=1.352
+ $Y2=2.7
cc_85 N_B_c_102_n N_A_27_115#_c_141_n 0.00249959f $X=0.95 $Y=2.31 $X2=1.352
+ $Y2=2.7
cc_86 B N_A_27_115#_c_141_n 0.00106496f $X=0.95 $Y=2.48 $X2=1.352 $Y2=2.7
cc_87 N_B_M1004_g N_A_27_115#_c_142_n 0.0223151f $X=0.905 $Y=3.445 $X2=1.352
+ $Y2=2.85
cc_88 N_B_M1001_g N_A_27_115#_c_148_n 0.0170493f $X=0.835 $Y=0.755 $X2=1.43
+ $Y2=1.755
cc_89 N_B_c_101_n N_A_27_115#_c_148_n 0.00242951f $X=0.95 $Y=2.31 $X2=1.43
+ $Y2=1.755
cc_90 N_B_c_102_n N_A_27_115#_c_148_n 0.00729726f $X=0.95 $Y=2.31 $X2=1.43
+ $Y2=1.755
cc_91 B N_A_27_115#_c_148_n 0.00785353f $X=0.95 $Y=2.48 $X2=1.43 $Y2=1.755
cc_92 N_B_M1001_g N_A_27_115#_c_150_n 0.00906251f $X=0.835 $Y=0.755 $X2=0.65
+ $Y2=3.025
cc_93 N_B_M1004_g N_A_27_115#_c_150_n 0.0103379f $X=0.905 $Y=3.445 $X2=0.65
+ $Y2=3.025
cc_94 N_B_c_102_n N_A_27_115#_c_150_n 0.0281763f $X=0.95 $Y=2.31 $X2=0.65
+ $Y2=3.025
cc_95 B N_A_27_115#_c_150_n 0.0027933f $X=0.95 $Y=2.48 $X2=0.65 $Y2=3.025
cc_96 N_B_c_101_n N_A_27_115#_c_160_n 4.41582e-19 $X=0.95 $Y=2.31 $X2=0.65
+ $Y2=3.195
cc_97 N_B_c_102_n N_Y_c_210_n 0.00431037f $X=0.95 $Y=2.31 $X2=1.55 $Y2=2.48
cc_98 B N_Y_c_210_n 9.40757e-19 $X=0.95 $Y=2.48 $X2=1.55 $Y2=2.48
cc_99 N_B_M1001_g Y 9.65944e-19 $X=0.835 $Y=0.755 $X2=1.555 $Y2=2.11
cc_100 N_B_c_102_n Y 0.00711983f $X=0.95 $Y=2.31 $X2=1.555 $Y2=2.11
cc_101 N_B_M1001_g N_Y_c_212_n 0.00101796f $X=0.835 $Y=0.755 $X2=1.55 $Y2=1.37
cc_102 N_B_c_102_n N_Y_c_213_n 9.85288e-19 $X=0.95 $Y=2.31 $X2=1.55 $Y2=2.48
cc_103 B N_Y_c_213_n 0.019951f $X=0.95 $Y=2.48 $X2=1.55 $Y2=2.48
cc_104 N_A_27_115#_M1000_g N_Y_c_208_n 0.0190376f $X=1.335 $Y=0.755 $X2=1.55
+ $Y2=0.74
cc_105 N_A_27_115#_c_140_n N_Y_c_208_n 0.0018791f $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=0.74
cc_106 N_A_27_115#_c_148_n N_Y_c_208_n 0.00712153f $X=1.43 $Y=1.755 $X2=1.55
+ $Y2=0.74
cc_107 N_A_27_115#_M1005_g N_Y_c_210_n 0.0088603f $X=1.335 $Y=3.445 $X2=1.55
+ $Y2=2.48
cc_108 N_A_27_115#_c_140_n N_Y_c_210_n 0.00131535f $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=2.48
cc_109 N_A_27_115#_c_141_n N_Y_c_210_n 0.0154438f $X=1.352 $Y=2.7 $X2=1.55
+ $Y2=2.48
cc_110 N_A_27_115#_c_148_n N_Y_c_210_n 0.00222212f $X=1.43 $Y=1.755 $X2=1.55
+ $Y2=2.48
cc_111 N_A_27_115#_M1000_g Y 0.00243059f $X=1.335 $Y=0.755 $X2=1.555 $Y2=2.11
cc_112 N_A_27_115#_c_140_n Y 0.00917711f $X=1.37 $Y=1.99 $X2=1.555 $Y2=2.11
cc_113 N_A_27_115#_c_141_n Y 0.00892438f $X=1.352 $Y=2.7 $X2=1.555 $Y2=2.11
cc_114 N_A_27_115#_c_148_n Y 0.0150696f $X=1.43 $Y=1.755 $X2=1.555 $Y2=2.11
cc_115 N_A_27_115#_M1000_g N_Y_c_212_n 0.00724699f $X=1.335 $Y=0.755 $X2=1.55
+ $Y2=1.37
cc_116 N_A_27_115#_c_140_n N_Y_c_212_n 0.00163148f $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=1.37
cc_117 N_A_27_115#_c_148_n N_Y_c_212_n 0.00257483f $X=1.43 $Y=1.755 $X2=1.55
+ $Y2=1.37
cc_118 N_A_27_115#_c_140_n N_Y_c_213_n 4.73507e-19 $X=1.37 $Y=1.99 $X2=1.55
+ $Y2=2.48
cc_119 N_A_27_115#_c_141_n N_Y_c_213_n 0.00583635f $X=1.352 $Y=2.7 $X2=1.55
+ $Y2=2.48
cc_120 N_A_27_115#_c_148_n N_Y_c_213_n 0.00169031f $X=1.43 $Y=1.755 $X2=1.55
+ $Y2=2.48
