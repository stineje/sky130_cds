* File: sky130_osu_sc_12T_ls__or2_4.spice
* Created: Fri Nov 12 15:39:49 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__or2_4.pex.spice"
.subckt sky130_osu_sc_12T_ls__or2_4  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1006 N_A_27_521#_M1006_d N_B_M1006_g N_GND_M1006_s N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75002.3 A=0.078 P=1.34 MULT=1
MM1000 N_GND_M1000_d N_A_M1000_g N_A_27_521#_M1006_d N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1001 N_Y_M1001_d N_A_27_521#_M1001_g N_GND_M1000_d N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75001.5 A=0.078 P=1.34 MULT=1
MM1008 N_Y_M1001_d N_A_27_521#_M1008_g N_GND_M1008_s N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.5
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1009 N_Y_M1009_d N_A_27_521#_M1009_g N_GND_M1008_s N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.9
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1011 N_Y_M1009_d N_A_27_521#_M1011_g N_GND_M1011_s N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75002.3
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1004 A_110_521# N_B_M1004_g N_A_27_521#_M1004_s N_VDD_M1004_b PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1010 N_VDD_M1010_d N_A_M1010_g A_110_521# N_VDD_M1004_b PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1002 N_VDD_M1010_d N_A_27_521#_M1002_g N_Y_M1002_s N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_27_521#_M1003_g N_Y_M1002_s N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1003_d N_A_27_521#_M1005_g N_Y_M1005_s N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_VDD_M1007_d N_A_27_521#_M1007_g N_Y_M1005_s N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1006_b N_VDD_M1004_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_8 B B PROBETYPE=1
pX14_noxref noxref_9 A A PROBETYPE=1
pX15_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__or2_4.pxi.spice"
*
.ends
*
*
