magic
tech sky130A
magscale 1 2
timestamp 1638894743
<< nwell >>
rect 78 529 1020 1119
<< nmoslvt >>
rect 171 115 201 263
rect 257 115 287 263
rect 329 115 359 263
rect 449 115 479 263
rect 521 115 551 263
rect 607 115 637 263
rect 815 115 845 218
rect 901 115 931 218
<< pmos >>
rect 171 595 201 995
rect 257 595 287 995
rect 329 595 359 995
rect 449 595 479 995
rect 521 595 551 995
rect 607 595 637 995
rect 815 743 845 995
rect 901 743 931 995
<< ndiff >>
rect 118 215 171 263
rect 118 131 126 215
rect 160 131 171 215
rect 118 115 171 131
rect 201 215 257 263
rect 201 131 212 215
rect 246 131 257 215
rect 201 115 257 131
rect 287 115 329 263
rect 359 215 449 263
rect 359 131 370 215
rect 438 131 449 215
rect 359 115 449 131
rect 479 115 521 263
rect 551 215 607 263
rect 551 131 562 215
rect 596 131 607 215
rect 551 115 607 131
rect 637 215 690 263
rect 637 131 648 215
rect 682 131 690 215
rect 637 115 690 131
rect 762 170 815 218
rect 762 131 770 170
rect 804 131 815 170
rect 762 115 815 131
rect 845 170 901 218
rect 845 131 856 170
rect 890 131 901 170
rect 845 115 901 131
rect 931 170 984 218
rect 931 131 942 170
rect 976 131 984 170
rect 931 115 984 131
<< pdiff >>
rect 118 979 171 995
rect 118 703 126 979
rect 160 703 171 979
rect 118 595 171 703
rect 201 979 257 995
rect 201 703 212 979
rect 246 703 257 979
rect 201 595 257 703
rect 287 595 329 995
rect 359 979 449 995
rect 359 635 370 979
rect 438 635 449 979
rect 359 595 449 635
rect 479 595 521 995
rect 551 979 607 995
rect 551 635 562 979
rect 596 635 607 979
rect 551 595 607 635
rect 637 979 690 995
rect 637 635 648 979
rect 682 635 690 979
rect 762 979 815 995
rect 762 783 770 979
rect 804 783 815 979
rect 762 743 815 783
rect 845 979 901 995
rect 845 783 856 979
rect 890 783 901 979
rect 845 743 901 783
rect 931 979 984 995
rect 931 783 942 979
rect 976 783 984 979
rect 931 743 984 783
rect 637 595 690 635
<< ndiffc >>
rect 126 131 160 215
rect 212 131 246 215
rect 370 131 438 215
rect 562 131 596 215
rect 648 131 682 215
rect 770 131 804 170
rect 856 131 890 170
rect 942 131 976 170
<< pdiffc >>
rect 126 703 160 979
rect 212 703 246 979
rect 370 635 438 979
rect 562 635 596 979
rect 648 635 682 979
rect 770 783 804 979
rect 856 783 890 979
rect 942 783 976 979
<< psubdiff >>
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
<< nsubdiff >>
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
rect 571 1049 595 1083
rect 629 1049 653 1083
rect 707 1049 731 1083
rect 765 1049 789 1083
rect 843 1049 867 1083
rect 901 1049 925 1083
<< psubdiffcont >>
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
<< nsubdiffcont >>
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
rect 595 1049 629 1083
rect 731 1049 765 1083
rect 867 1049 901 1083
<< poly >>
rect 171 995 201 1021
rect 257 995 287 1021
rect 329 995 359 1021
rect 449 995 479 1021
rect 521 995 551 1021
rect 607 995 637 1021
rect 815 995 845 1021
rect 901 995 931 1021
rect 815 727 845 743
rect 805 697 845 727
rect 171 543 201 595
rect 161 509 201 543
rect 161 351 191 509
rect 257 466 287 595
rect 329 534 359 595
rect 449 534 479 595
rect 329 518 383 534
rect 329 484 339 518
rect 373 484 383 518
rect 329 468 383 484
rect 425 518 479 534
rect 425 484 435 518
rect 469 484 479 518
rect 425 468 479 484
rect 233 450 287 466
rect 233 416 243 450
rect 277 416 287 450
rect 425 423 455 468
rect 233 400 287 416
rect 161 335 215 351
rect 161 301 171 335
rect 205 301 215 335
rect 161 285 215 301
rect 171 263 201 285
rect 257 263 287 400
rect 329 393 455 423
rect 521 425 551 595
rect 607 534 637 595
rect 607 518 678 534
rect 607 504 634 518
rect 618 484 634 504
rect 668 484 678 518
rect 618 468 678 484
rect 521 409 575 425
rect 329 263 359 393
rect 521 375 531 409
rect 565 375 575 409
rect 521 359 575 375
rect 425 335 479 351
rect 425 301 435 335
rect 469 301 479 335
rect 425 285 479 301
rect 449 263 479 285
rect 521 263 551 359
rect 618 311 648 468
rect 805 425 835 697
rect 901 425 931 743
rect 780 409 835 425
rect 780 375 790 409
rect 824 375 835 409
rect 780 359 835 375
rect 877 409 931 425
rect 877 375 887 409
rect 921 375 931 409
rect 877 359 931 375
rect 607 281 648 311
rect 805 308 835 359
rect 607 263 637 281
rect 805 278 845 308
rect 815 218 845 278
rect 901 218 931 359
rect 171 89 201 115
rect 257 89 287 115
rect 329 89 359 115
rect 449 89 479 115
rect 521 89 551 115
rect 607 89 637 115
rect 815 89 845 115
rect 901 89 931 115
<< polycont >>
rect 339 484 373 518
rect 435 484 469 518
rect 243 416 277 450
rect 171 301 205 335
rect 634 484 668 518
rect 531 375 565 409
rect 435 301 469 335
rect 790 375 824 409
rect 887 375 921 409
<< locali >>
rect 86 1089 1017 1110
rect 86 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 595 1089
rect 629 1049 731 1089
rect 765 1049 867 1089
rect 901 1049 1017 1089
rect 126 979 160 995
rect 103 703 126 769
rect 103 686 160 703
rect 212 979 246 1049
rect 212 687 246 703
rect 370 979 438 995
rect 103 409 137 686
rect 370 632 438 635
rect 103 244 137 375
rect 171 598 438 632
rect 562 979 596 1049
rect 562 619 596 635
rect 648 979 682 995
rect 770 979 804 995
rect 770 735 804 783
rect 856 979 890 1049
rect 856 767 890 783
rect 942 979 976 995
rect 976 775 989 792
rect 942 758 989 775
rect 770 696 804 701
rect 770 662 921 696
rect 648 632 682 635
rect 648 598 736 632
rect 171 335 205 598
rect 435 518 469 534
rect 323 484 339 518
rect 373 484 389 518
rect 243 400 277 416
rect 355 335 389 484
rect 435 483 469 484
rect 634 518 668 534
rect 634 483 668 484
rect 702 409 736 598
rect 887 409 921 662
rect 515 375 531 409
rect 565 375 581 409
rect 648 375 736 409
rect 774 375 790 409
rect 824 375 840 409
rect 648 335 682 375
rect 887 335 921 375
rect 205 301 314 335
rect 355 301 435 335
rect 469 301 682 335
rect 171 285 205 301
rect 280 251 314 301
rect 103 215 160 244
rect 103 210 126 215
rect 126 115 160 131
rect 212 215 246 231
rect 280 217 438 251
rect 212 61 246 131
rect 370 215 438 217
rect 370 115 438 131
rect 562 215 596 231
rect 562 61 596 131
rect 648 215 682 301
rect 648 115 682 131
rect 770 301 921 335
rect 770 170 804 301
rect 955 222 989 758
rect 942 188 989 222
rect 770 115 804 131
rect 856 170 890 186
rect 856 61 890 131
rect 942 170 976 188
rect 942 115 976 131
rect 71 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1017 61
rect 71 0 1017 21
<< viali >>
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 595 1083 629 1089
rect 595 1055 629 1083
rect 731 1083 765 1089
rect 731 1055 765 1083
rect 867 1083 901 1089
rect 867 1055 901 1083
rect 103 375 137 409
rect 942 783 976 809
rect 942 775 976 783
rect 770 701 804 735
rect 243 450 277 484
rect 435 449 469 483
rect 634 449 668 483
rect 531 375 565 409
rect 790 375 824 409
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
<< metal1 >>
rect 86 1089 1017 1110
rect 86 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 595 1089
rect 629 1055 731 1089
rect 765 1055 867 1089
rect 901 1055 1017 1089
rect 86 1049 1017 1055
rect 930 809 988 815
rect 907 775 942 809
rect 976 775 988 809
rect 930 769 988 775
rect 758 735 816 741
rect 751 734 770 735
rect 736 702 770 734
rect 751 701 770 702
rect 804 701 816 735
rect 758 695 816 701
rect 231 484 290 490
rect 231 450 243 484
rect 277 450 310 484
rect 423 483 481 489
rect 622 483 680 489
rect 231 444 290 450
rect 423 449 435 483
rect 469 449 634 483
rect 668 449 680 483
rect 423 443 481 449
rect 622 443 680 449
rect 90 409 149 415
rect 90 375 103 409
rect 137 402 149 409
rect 519 409 578 415
rect 519 402 531 409
rect 137 375 531 402
rect 565 406 578 409
rect 778 409 836 415
rect 778 406 790 409
rect 565 378 790 406
rect 565 375 578 378
rect 90 374 578 375
rect 90 369 149 374
rect 519 369 578 374
rect 778 375 790 378
rect 824 375 836 409
rect 778 369 836 375
rect 71 55 1017 61
rect 71 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1017 55
rect 71 0 1017 21
<< labels >>
rlabel metal1 651 466 651 466 1 CK
port 1 n
rlabel metal1 260 466 260 466 1 D
port 2 n
rlabel viali 959 792 959 792 1 Q
port 3 n
rlabel viali 788 718 788 718 1 QN
port 4 n
<< end >>
