* File: sky130_osu_sc_18T_ls__addh_l.pex.spice
* Created: Fri Nov 12 14:13:11 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%GND 1 2 45 47 55 57 70 86 88
r96 86 88 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r97 72 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.152
+ $X2=2.56 $Y2=0.152
r98 68 82 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.152
r99 68 70 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.56 $Y=0.305
+ $X2=2.56 $Y2=0.825
r100 58 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.152
+ $X2=0.75 $Y2=0.152
r101 57 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.152
+ $X2=2.56 $Y2=0.152
r102 53 81 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.152
r103 53 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=0.305
+ $X2=0.75 $Y2=0.825
r104 47 81 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.152
+ $X2=0.75 $Y2=0.152
r105 45 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.19
+ $X2=3.74 $Y2=0.19
r106 45 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r107 45 72 15.6808 $w=3.03e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.645 $Y2=0.152
r108 45 57 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.475 $Y2=0.152
r109 45 58 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.835 $Y2=0.152
r110 45 47 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.665 $Y2=0.152
r111 2 70 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.575 $X2=2.56 $Y2=0.825
r112 1 55 91 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.75 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%VDD 1 2 3 37 39 46 50 56 60 68 74 82 86
r58 82 86 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.74 $Y2=6.507
r59 74 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=6.47
+ $X2=3.74 $Y2=6.47
r60 72 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.05 $Y2=6.507
r61 72 74 22.8599 $w=3.03e-07 $l=6.05e-07 $layer=LI1_cond $X=3.135 $Y=6.507
+ $X2=3.74 $Y2=6.507
r62 68 71 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.05 $Y=3.455
+ $X2=3.05 $Y2=5.835
r63 66 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=6.507
r64 66 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.05 $Y=6.355
+ $X2=3.05 $Y2=5.835
r65 63 65 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=6.507
+ $X2=2.38 $Y2=6.507
r66 61 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.61 $Y2=6.507
r67 61 63 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=1.695 $Y=6.507
+ $X2=1.7 $Y2=6.507
r68 60 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=3.05 $Y2=6.507
r69 60 65 22.1042 $w=3.03e-07 $l=5.85e-07 $layer=LI1_cond $X=2.965 $Y=6.507
+ $X2=2.38 $Y2=6.507
r70 56 59 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.61 $Y=3.795
+ $X2=1.61 $Y2=5.835
r71 54 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=6.507
r72 54 59 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.61 $Y=6.355
+ $X2=1.61 $Y2=5.835
r73 51 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=0.75 $Y2=6.507
r74 51 53 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=0.835 $Y=6.507
+ $X2=1.02 $Y2=6.507
r75 50 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.61 $Y2=6.507
r76 50 53 19.0814 $w=3.03e-07 $l=5.05e-07 $layer=LI1_cond $X=1.525 $Y=6.507
+ $X2=1.02 $Y2=6.507
r77 46 49 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.75 $Y=3.455
+ $X2=0.75 $Y2=5.835
r78 44 77 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=6.507
r79 44 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.75 $Y=6.355
+ $X2=0.75 $Y2=5.835
r80 41 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r81 39 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.75 $Y2=6.507
r82 39 41 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=0.665 $Y=6.507
+ $X2=0.34 $Y2=6.507
r83 37 74 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r84 37 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r85 37 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r86 37 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r87 37 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r88 37 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r89 3 59 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=5.835
r90 3 56 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.47
+ $Y=3.085 $X2=1.61 $Y2=3.795
r91 2 49 150 $w=1.7e-07 $l=1.49666e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=4.435 $X2=0.75 $Y2=5.835
r92 2 46 150 $w=1.7e-07 $l=1.07536e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=4.435 $X2=0.75 $Y2=3.455
r93 1 71 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=5.835
r94 1 68 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=3.085 $X2=3.05 $Y2=3.455
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%CON 1 3 4 15 19 22 29 31 32 35 39 41 43
+ 45 49 55 58 59 64 67
c128 67 0 2.7119e-19 $X=3.42 $Y=1.85
c129 59 0 1.57622e-19 $X=0.78 $Y=1.85
c130 43 0 1.92558e-19 $X=3.42 $Y=1.765
r131 59 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.78 $Y=1.85
+ $X2=0.635 $Y2=1.85
r132 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=2.62 $Y2=1.85
r133 58 59 1.63209 $w=1.7e-07 $l=1.695e-06 $layer=MET1_cond $X=2.475 $Y=1.85
+ $X2=0.78 $Y2=1.85
r134 57 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=1.85
+ $X2=3.42 $Y2=1.85
r135 54 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.62 $Y=1.85
+ $X2=2.62 $Y2=1.85
r136 49 51 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.84 $Y=3.455
+ $X2=3.84 $Y2=5.835
r137 47 49 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.84 $Y=3.035
+ $X2=3.84 $Y2=3.455
r138 43 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.85
r139 43 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.42 $Y=1.765
+ $X2=3.42 $Y2=1.165
r140 42 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.95
+ $X2=2.62 $Y2=2.95
r141 41 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=3.84 $Y2=3.035
r142 41 42 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.755 $Y=2.95
+ $X2=2.705 $Y2=2.95
r143 40 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.85
+ $X2=2.62 $Y2=1.85
r144 39 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=3.42 $Y2=1.85
r145 39 40 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.335 $Y=1.85
+ $X2=2.705 $Y2=1.85
r146 35 37 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.62 $Y=3.455
+ $X2=2.62 $Y2=5.835
r147 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=2.95
r148 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.62 $Y=3.035
+ $X2=2.62 $Y2=3.455
r149 32 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.865
+ $X2=2.62 $Y2=2.95
r150 31 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=1.85
r151 31 32 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.62 $Y=1.935
+ $X2=2.62 $Y2=2.865
r152 29 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=1.85
+ $X2=0.635 $Y2=1.85
r153 26 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.35 $Y=1.85
+ $X2=0.635 $Y2=1.85
r154 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.85 $X2=0.35 $Y2=1.85
r155 22 24 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=2.015
r156 22 23 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.85
+ $X2=0.382 $Y2=1.685
r157 19 24 1663.93 $w=1.5e-07 $l=3.245e-06 $layer=POLY_cond $X=0.475 $Y=5.26
+ $X2=0.475 $Y2=2.015
r158 15 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=1.685
r159 4 51 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=5.835
r160 4 49 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.7
+ $Y=3.085 $X2=3.84 $Y2=3.455
r161 3 37 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=5.835
r162 3 35 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=2.495
+ $Y=3.085 $X2=2.62 $Y2=3.455
r163 1 45 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.575 $X2=3.42 $Y2=1.165
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%B 3 7 11 15 18 22 25 30 39 42 44
c101 44 0 4.99902e-20 $X=3.21 $Y=2.22
c102 22 0 1.42567e-19 $X=3.205 $Y=2.22
c103 18 0 1.57622e-19 $X=0.905 $Y=2.22
r104 41 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=3.205 $Y=2.22
+ $X2=3.21 $Y2=2.22
r105 41 42 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.205 $Y=2.22
+ $X2=3.06 $Y2=2.22
r106 39 42 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.05 $Y=2.222
+ $X2=3.06 $Y2=2.222
r107 37 39 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.905 $Y=2.22
+ $X2=1.05 $Y2=2.22
r108 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.22
r109 25 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.22
r110 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=2.22 $X2=3.205 $Y2=2.22
r111 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.22
+ $X2=3.205 $Y2=2.385
r112 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=2.22 $X2=0.905 $Y2=2.22
r113 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.385
r114 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.22
+ $X2=0.905 $Y2=2.055
r115 15 23 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=3.265 $Y=4.585
+ $X2=3.265 $Y2=2.385
r116 9 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=2.22
r117 9 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.205 $Y=2.055
+ $X2=3.205 $Y2=1.075
r118 7 20 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=0.965 $Y=4.585
+ $X2=0.965 $Y2=2.385
r119 3 19 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.965 $Y=1.075
+ $X2=0.965 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%A 3 7 11 15 18 22 26 31 40 42 43
c87 22 0 1.74252e-19 $X=3.685 $Y=2.59
r88 42 43 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.685 $Y=2.59
+ $X2=3.54 $Y2=2.59
r89 40 43 1.81922 $w=1.75e-07 $l=2.01e-06 $layer=MET1_cond $X=1.53 $Y=2.587
+ $X2=3.54 $Y2=2.587
r90 38 40 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.385 $Y=2.59
+ $X2=1.53 $Y2=2.59
r91 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.59
r92 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.59
r93 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=2.59 $X2=3.685 $Y2=2.59
r94 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.755
r95 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=2.59
+ $X2=3.685 $Y2=2.425
r96 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=2.59 $X2=1.385 $Y2=2.59
r97 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.755
r98 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.59
+ $X2=1.385 $Y2=2.425
r99 15 23 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=3.635 $Y=1.075
+ $X2=3.635 $Y2=2.425
r100 11 24 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.625 $Y=4.585
+ $X2=3.625 $Y2=2.755
r101 7 20 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=1.395 $Y=4.585
+ $X2=1.395 $Y2=2.755
r102 3 19 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=1.325 $Y=1.075
+ $X2=1.325 $Y2=2.425
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%A_208_617# 1 3 10 13 15 17 21 23 27 31
+ 33 38 39 42 46 47 50 53 55
c114 31 0 2.52869e-20 $X=2.835 $Y=4.585
c115 23 0 9.69384e-20 $X=2.7 $Y=1.8
r116 55 57 4.62121 $w=2.64e-07 $l=1e-07 $layer=LI1_cond $X=1.725 $Y=1.955
+ $X2=1.825 $Y2=1.955
r117 54 55 8.54924 $w=2.64e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.955
+ $X2=1.725 $Y2=1.955
r118 52 55 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=1.955
r119 52 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.725 $Y=2.12
+ $X2=1.725 $Y2=2.925
r120 48 54 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=1.955
r121 48 50 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.54 $Y=1.79
+ $X2=1.54 $Y2=0.825
r122 46 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.725 $Y2=2.925
r123 46 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.64 $Y=3.01
+ $X2=1.265 $Y2=3.01
r124 42 44 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.18 $Y=3.795
+ $X2=1.18 $Y2=5.835
r125 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.265 $Y2=3.01
r126 40 42 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.18 $Y=3.095
+ $X2=1.18 $Y2=3.795
r127 36 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.955 $X2=1.825 $Y2=1.955
r128 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.955
+ $X2=1.825 $Y2=2.12
r129 33 36 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.8
+ $X2=1.825 $Y2=1.955
r130 29 31 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=2.835 $Y=2.745
+ $X2=2.835 $Y2=4.585
r131 25 27 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=1.075
r132 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.8
+ $X2=2.285 $Y2=1.8
r133 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=1.8
+ $X2=2.775 $Y2=1.725
r134 23 24 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.8 $X2=2.36
+ $Y2=1.8
r135 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=1.8
r136 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.285 $Y=1.725
+ $X2=2.285 $Y2=0.895
r137 18 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=2.67
+ $X2=1.885 $Y2=2.67
r138 17 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=2.67
+ $X2=2.835 $Y2=2.745
r139 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.76 $Y=2.67 $X2=1.96
+ $Y2=2.67
r140 16 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.8
+ $X2=1.825 $Y2=1.8
r141 15 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=2.285 $Y2=1.8
r142 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.21 $Y=1.8
+ $X2=1.96 $Y2=1.8
r143 11 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=2.67
r144 11 13 1289.61 $w=1.5e-07 $l=2.515e-06 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=5.26
r145 10 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.67
r146 10 37 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.885 $Y=2.595
+ $X2=1.885 $Y2=2.12
r147 3 44 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=5.835
r148 3 42 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.04
+ $Y=3.085 $X2=1.18 $Y2=3.795
r149 1 50 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.575 $X2=1.54 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%S 1 3 10 16 26 29 32
r32 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=3.33
r33 24 26 0.799192 $w=1.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=2.385
r34 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=1.475
r35 23 26 0.765491 $w=1.7e-07 $l=7.95e-07 $layer=MET1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=2.385
r36 19 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=4.815
+ $X2=0.26 $Y2=5.835
r37 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=3.33
r38 16 19 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=0.26 $Y=3.33
+ $X2=0.26 $Y2=4.815
r39 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=1.475
+ $X2=0.26 $Y2=1.475
r40 10 13 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.26 $Y=0.825
+ $X2=0.26 $Y2=1.475
r41 3 21 300 $w=1.7e-07 $l=1.46116e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.435 $X2=0.26 $Y2=5.835
r42 3 19 300 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.435 $X2=0.26 $Y2=4.815
r43 1 10 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%CO 1 3 11 15 23 26 27 30
c55 26 0 2.52869e-20 $X=2.175 $Y=2.96
r56 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.175 $Y=2.96
+ $X2=2.175 $Y2=2.96
r57 26 28 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=3.045
r58 26 27 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.96
+ $X2=2.137 $Y2=2.875
r59 21 23 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.472
+ $X2=2.175 $Y2=1.472
r60 19 23 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=1.472
r61 19 27 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.175 $Y=1.56
+ $X2=2.175 $Y2=2.875
r62 15 17 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.1 $Y=4.815
+ $X2=2.1 $Y2=5.835
r63 15 28 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=2.1 $Y=4.815
+ $X2=2.1 $Y2=3.045
r64 9 21 0.89264 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.07 $Y=1.385 $X2=2.07
+ $Y2=1.472
r65 9 11 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.07 $Y=1.385
+ $X2=2.07 $Y2=0.825
r66 3 17 300 $w=1.7e-07 $l=1.46833e-06 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=4.435 $X2=2.1 $Y2=5.835
r67 3 15 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=4.435 $X2=2.1 $Y2=4.815
r68 1 11 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.575 $X2=2.07 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDH_L%A_570_115# 1 2 11 13 14
r11 15 17 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.85 $Y=0.72
+ $X2=3.85 $Y2=0.825
r12 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.85 $Y2=0.72
r13 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.635
+ $X2=3.075 $Y2=0.635
r14 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.72
+ $X2=3.075 $Y2=0.635
r15 9 11 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.72
+ $X2=2.99 $Y2=0.825
r16 2 17 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.575 $X2=3.85 $Y2=0.825
r17 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.575 $X2=2.99 $Y2=0.825
.ends

