* File: sky130_osu_sc_12T_hs__xor2_l.pex.spice
* Created: Fri Nov 12 15:14:16 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%GND 1 2 33 35 43 45 55 67 69
r66 67 69 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r67 53 55 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.755
r68 46 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r69 41 59 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r70 41 43 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.755
r71 35 59 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r72 33 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r73 33 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r74 33 53 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r75 33 45 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r76 33 45 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r77 33 46 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r78 33 35 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r79 2 55 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.3 $Y=0.575
+ $X2=2.44 $Y2=0.755
r80 1 43 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.575
+ $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%VDD 1 2 25 27 34 36 44 50 53 57
r45 53 57 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=2.38 $Y2=4.287
r46 50 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=4.25
+ $X2=2.38 $Y2=4.25
r47 42 50 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=4.135
+ $X2=2.44 $Y2=4.287
r48 42 44 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.44 $Y=4.135 $X2=2.44
+ $Y2=3.635
r49 39 41 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=4.287
+ $X2=1.7 $Y2=4.287
r50 37 48 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=0.69 $Y2=4.287
r51 37 39 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=4.287
+ $X2=1.02 $Y2=4.287
r52 36 50 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=4.287
+ $X2=2.44 $Y2=4.287
r53 36 41 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=4.287
+ $X2=1.7 $Y2=4.287
r54 32 48 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=4.287
r55 32 34 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=4.135 $X2=0.69
+ $Y2=3.635
r56 29 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r57 27 48 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.69 $Y2=4.287
r58 27 29 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=4.287
+ $X2=0.34 $Y2=4.287
r59 25 50 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r60 25 41 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r61 25 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r62 25 29 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r63 2 44 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.605 $X2=2.44 $Y2=3.635
r64 1 34 600 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%A_27_115# 1 3 11 15 18 22 27 31 35 41 43
c76 41 0 6.74854e-20 $X=1.805 $Y=2.285
c77 35 0 1.52002e-20 $X=1.72 $Y=1.745
r78 39 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.805 $Y=1.83
+ $X2=1.805 $Y2=2.285
r79 36 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.745
+ $X2=0.26 $Y2=1.745
r80 36 38 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=1.745
+ $X2=0.845 $Y2=1.745
r81 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=1.745
+ $X2=1.805 $Y2=1.83
r82 35 38 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.72 $Y=1.745
+ $X2=0.845 $Y2=1.745
r83 31 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.955
+ $X2=0.26 $Y2=3.635
r84 29 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.83 $X2=0.26
+ $Y2=1.745
r85 29 31 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=0.26 $Y=1.83
+ $X2=0.26 $Y2=2.955
r86 25 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.66 $X2=0.26
+ $Y2=1.745
r87 25 27 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=0.755
r88 22 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=2.285 $X2=1.805 $Y2=2.285
r89 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=2.285
+ $X2=1.805 $Y2=2.45
r90 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=1.745 $X2=0.845 $Y2=1.745
r91 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=1.745
+ $X2=0.845 $Y2=1.58
r92 15 24 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.865 $Y=3.235
+ $X2=1.865 $Y2=2.45
r93 11 19 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.905 $Y=0.85
+ $X2=0.905 $Y2=1.58
r94 3 33 400 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
r95 3 31 400 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=2.955
r96 1 27 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%A 2 5 6 8 9 13 16 18 19 20 21 22 24 27
+ 28 34 37 40 45 50 52 53 58 61
c122 50 0 3.33037e-19 $X=2.235 $Y=1.74
r123 55 58 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=1.085 $Y=2.85
+ $X2=1.09 $Y2=2.85
r124 53 58 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=1.23 $Y=2.85
+ $X2=1.09 $Y2=2.85
r125 52 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2 $Y=2.85
+ $X2=2.145 $Y2=2.85
r126 52 53 0.741419 $w=1.7e-07 $l=7.7e-07 $layer=MET1_cond $X=2 $Y=2.85 $X2=1.23
+ $Y2=2.85
r127 47 50 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.145 $Y=1.74
+ $X2=2.235 $Y2=1.74
r128 45 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=2.85
+ $X2=1.085 $Y2=2.85
r129 42 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.845 $Y=2.85
+ $X2=1.085 $Y2=2.85
r130 37 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=2.85
+ $X2=2.145 $Y2=2.85
r131 35 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.825
+ $X2=2.145 $Y2=1.74
r132 35 37 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.145 $Y=1.825
+ $X2=2.145 $Y2=2.85
r133 34 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=2.765
+ $X2=0.845 $Y2=2.85
r134 33 40 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=2.37
+ $X2=0.845 $Y2=2.285
r135 33 34 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.845 $Y=2.37
+ $X2=0.845 $Y2=2.765
r136 31 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.74 $X2=2.235 $Y2=1.74
r137 28 31 23.3282 $w=2.7e-07 $l=1.05e-07 $layer=POLY_cond $X=2.235 $Y=1.635
+ $X2=2.235 $Y2=1.74
r138 26 27 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=2.455
+ $X2=0.845 $Y2=2.53
r139 24 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.285 $X2=0.845 $Y2=2.285
r140 24 26 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=0.845 $Y=2.285
+ $X2=0.845 $Y2=2.455
r141 20 21 41.4471 $w=2e-07 $l=1.25e-07 $layer=POLY_cond $X=0.45 $Y=1.2 $X2=0.45
+ $Y2=1.325
r142 18 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.1 $Y=1.635
+ $X2=2.235 $Y2=1.635
r143 18 19 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.1 $Y=1.635
+ $X2=1.94 $Y2=1.635
r144 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.865 $Y=1.56
+ $X2=1.94 $Y2=1.635
r145 14 16 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.865 $Y=1.56
+ $X2=1.865 $Y2=0.85
r146 13 27 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=3.235
+ $X2=0.905 $Y2=2.53
r147 10 22 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=2.455
+ $X2=0.45 $Y2=2.455
r148 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=2.455
+ $X2=0.845 $Y2=2.455
r149 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=2.455
+ $X2=0.55 $Y2=2.455
r150 6 22 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=2.53
+ $X2=0.45 $Y2=2.455
r151 6 8 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.475 $Y=2.53
+ $X2=0.475 $Y2=3.235
r152 5 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.475 $Y=0.85
+ $X2=0.475 $Y2=1.2
r153 2 22 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=2.38
+ $X2=0.45 $Y2=2.455
r154 2 21 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.425 $Y=2.38
+ $X2=0.425 $Y2=1.325
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%A_238_89# 1 3 11 14 17 18 20 26 30 34
r64 30 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.87 $Y=2.955
+ $X2=2.87 $Y2=3.635
r65 28 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.485
+ $X2=2.87 $Y2=1.4
r66 28 30 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=2.87 $Y=1.485
+ $X2=2.87 $Y2=2.955
r67 24 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.315
+ $X2=2.87 $Y2=1.4
r68 24 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.87 $Y=1.315
+ $X2=2.87 $Y2=0.755
r69 20 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.4 $X2=2.87
+ $Y2=1.4
r70 20 22 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=1.4
+ $X2=1.325 $Y2=1.4
r71 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.4 $X2=1.325 $Y2=1.4
r72 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.4
+ $X2=1.325 $Y2=1.565
r73 17 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.4
+ $X2=1.325 $Y2=1.235
r74 14 19 856.319 $w=1.5e-07 $l=1.67e-06 $layer=POLY_cond $X=1.265 $Y=3.235
+ $X2=1.265 $Y2=1.565
r75 11 18 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.265 $Y=0.85
+ $X2=1.265 $Y2=1.235
r76 3 32 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.605 $X2=2.87 $Y2=3.635
r77 3 30 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.605 $X2=2.87 $Y2=2.955
r78 1 26 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.73 $Y=0.575
+ $X2=2.87 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 20 21 23 29
c56 20 0 6.74854e-20 $X=2.655 $Y=2.325
c57 13 0 1.52002e-20 $X=2.655 $Y=2.12
c58 8 0 1.82321e-19 $X=2.3 $Y=1.275
c59 7 0 1.50716e-19 $X=2.58 $Y=1.275
r60 26 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.48
+ $X2=2.53 $Y2=2.48
r61 23 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.53 $Y=2.285
+ $X2=2.53 $Y2=2.48
r62 19 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=2.285 $X2=2.53 $Y2=2.285
r63 19 20 20.0833 $w=3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=2.325
+ $X2=2.655 $Y2=2.325
r64 14 20 18.9685 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.655 $Y=2.53
+ $X2=2.655 $Y2=2.325
r65 14 16 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.655 $Y=2.53
+ $X2=2.655 $Y2=3.235
r66 13 20 18.9685 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.655 $Y=2.12
+ $X2=2.655 $Y2=2.325
r67 12 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.35
+ $X2=2.655 $Y2=1.275
r68 12 13 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.655 $Y=1.35
+ $X2=2.655 $Y2=2.12
r69 9 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.2
+ $X2=2.655 $Y2=1.275
r70 9 11 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.655 $Y=1.2
+ $X2=2.655 $Y2=0.85
r71 7 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.275
+ $X2=2.655 $Y2=1.275
r72 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=1.275 $X2=2.3
+ $Y2=1.275
r73 4 19 49.0033 $w=3e-07 $l=3.94398e-07 $layer=POLY_cond $X=2.225 $Y=2.53
+ $X2=2.53 $Y2=2.325
r74 4 6 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.225 $Y=2.53
+ $X2=2.225 $Y2=3.235
r75 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=1.2
+ $X2=2.3 $Y2=1.275
r76 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.225 $Y=1.2 $X2=2.225
+ $Y2=0.85
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__XOR2_L%Y 1 3 11 15 20 22 28 31 33
r58 33 35 0.0784753 $w=2.23e-07 $l=1.4e-07 $layer=MET1_cond $X=1.425 $Y=1
+ $X2=1.565 $Y2=1
r59 26 31 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.995
+ $X2=1.425 $Y2=2.11
r60 26 28 0.0433297 $w=1.7e-07 $l=4.5e-08 $layer=MET1_cond $X=1.425 $Y=1.995
+ $X2=1.425 $Y2=1.95
r61 25 33 0.0238602 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.115
+ $X2=1.425 $Y2=1
r62 25 28 0.804007 $w=1.7e-07 $l=8.35e-07 $layer=MET1_cond $X=1.425 $Y=1.115
+ $X2=1.425 $Y2=1.95
r63 24 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.565 $Y=1 $X2=1.565
+ $Y2=1
r64 22 24 10.3069 $w=2.9e-07 $l=2.45e-07 $layer=LI1_cond $X=1.565 $Y=0.755
+ $X2=1.565 $Y2=1
r65 19 20 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.537 $Y=2.725
+ $X2=1.537 $Y2=2.895
r66 15 17 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=1.565 $Y=2.955
+ $X2=1.565 $Y2=3.635
r67 15 20 2.03372 $w=3.38e-07 $l=6e-08 $layer=LI1_cond $X=1.565 $Y=2.955
+ $X2=1.565 $Y2=2.895
r68 11 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=2.11
+ $X2=1.425 $Y2=2.11
r69 11 19 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.425 $Y=2.11
+ $X2=1.425 $Y2=2.725
r70 3 17 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.565 $Y2=3.635
r71 3 15 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.605 $X2=1.565 $Y2=2.955
r72 1 22 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.755
.ends

