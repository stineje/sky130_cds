* File: sky130_osu_sc_18T_ls__buf_6.pex.spice
* Created: Thu Oct 29 17:35:01 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_1 1 2 3 4 33 35 42 44 51 53 60 62
+ 69 71 72
r86 67 69 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.825
r87 62 67 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=3.185 $Y=0.152
+ $X2=3.27 $Y2=0.305
r88 58 60 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.825
r89 54 72 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0.152
+ $X2=1.55 $Y2=0.152
r90 49 72 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.152
r91 49 51 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.825
r92 45 71 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r93 44 72 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.152
r94 40 71 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r95 40 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r96 35 71 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r97 33 58 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.41 $Y2=0.305
r98 33 53 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.325 $Y2=0.152
r99 33 63 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.495 $Y2=0.152
r100 33 62 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.185 $Y2=0.152
r101 33 63 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.495 $Y2=0.152
r102 33 53 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r103 33 54 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r104 33 44 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r105 33 45 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r106 33 35 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r107 4 69 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.825
r108 3 60 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r109 2 51 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r110 1 42 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%noxref_2 1 2 3 4 28 30 36 40 46 50 56 60
+ 66 70 71 73
r60 66 69 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.27 $Y=3.455
+ $X2=3.27 $Y2=5.835
r61 64 69 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=6.355
+ $X2=3.27 $Y2=5.835
r62 61 73 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=2.41 $Y2=6.507
r63 61 63 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=3.06 $Y2=6.507
r64 60 64 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.27 $Y2=6.355
r65 60 63 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.06 $Y2=6.507
r66 56 59 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r67 54 73 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=6.507
r68 54 59 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=5.835
r69 51 71 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.55 $Y2=6.507
r70 51 53 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.7 $Y2=6.507
r71 50 73 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=2.41 $Y2=6.507
r72 50 53 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=1.7 $Y2=6.507
r73 46 49 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r74 44 71 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=6.507
r75 44 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=5.835
r76 41 70 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r77 41 43 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r78 40 71 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.55 $Y2=6.507
r79 40 43 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.02 $Y2=6.507
r80 36 39 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r81 34 70 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r82 34 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r83 30 70 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r84 30 32 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r85 28 73 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r86 28 63 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r87 28 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r88 28 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r89 28 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r90 4 69 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=5.835
r91 4 66 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=3.455
r92 3 59 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r93 3 56 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r94 2 49 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r95 2 46 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r96 1 39 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r97 1 36 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%A 3 7 10 15 16
r40 16 18 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.645
r41 16 17 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.315
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.48 $X2=0.635 $Y2=2.48
r43 12 15 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=2.48
r44 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=3.33
r45 7 18 994.766 $w=1.5e-07 $l=1.94e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.645
r46 3 17 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.315
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%A_27_115# 1 2 9 11 13 15 18 20 22 23 24
+ 25 26 29 31 33 34 36 40 42 44 45 47 51 54 55 57 58 60 64 66 68 73 74 75 76 77
+ 78 81 85 89 91 94
c177 55 0 1.33323e-19 $X=2.625 $Y=3.01
c178 51 0 1.33323e-19 $X=2.625 $Y=1.075
c179 42 0 1.33323e-19 $X=2.195 $Y=3.01
c180 40 0 1.33323e-19 $X=2.195 $Y=1.075
c181 31 0 1.33323e-19 $X=1.765 $Y=3.01
c182 29 0 1.33323e-19 $X=1.765 $Y=1.075
c183 20 0 1.33323e-19 $X=1.335 $Y=3.01
c184 18 0 1.33323e-19 $X=1.335 $Y=1.075
r185 95 99 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=1.18 $Y2=1.935
r186 95 97 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=0.905 $Y2=1.935
r187 94 95 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.935 $X2=0.965 $Y2=1.935
r188 90 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.935
+ $X2=0.26 $Y2=1.935
r189 89 94 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.965 $Y2=1.935
r190 89 90 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.345 $Y2=1.935
r191 85 87 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r192 83 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=1.935
r193 83 85 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=3.455
r194 79 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=1.935
r195 79 81 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r196 71 72 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.935
+ $X2=1.335 $Y2=2.935
r197 69 71 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.935
+ $X2=1.18 $Y2=2.935
r198 66 68 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.055 $Y=3.01
+ $X2=3.055 $Y2=4.585
r199 62 64 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.075
r200 61 78 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.935 $X2=2.625
+ $Y2=2.935
r201 60 66 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=3.055 $Y2=3.01
r202 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=2.7 $Y2=2.935
r203 59 77 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.845 $X2=2.625
+ $Y2=1.845
r204 58 62 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=3.055 $Y2=1.77
r205 58 59 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=2.7 $Y2=1.845
r206 55 78 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=2.935
r207 55 57 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=4.585
r208 54 78 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.86
+ $X2=2.625 $Y2=2.935
r209 53 77 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.92
+ $X2=2.625 $Y2=1.845
r210 53 54 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.625 $Y=1.92 $X2=2.625
+ $Y2=2.86
r211 49 77 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.845
r212 49 51 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.075
r213 48 76 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.935
+ $X2=2.195 $Y2=2.935
r214 47 78 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.625 $Y2=2.935
r215 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.27 $Y2=2.935
r216 46 75 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.195 $Y2=1.845
r217 45 77 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.625 $Y2=1.845
r218 45 46 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.27 $Y2=1.845
r219 42 76 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=2.935
r220 42 44 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=4.585
r221 38 75 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.845
r222 38 40 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r223 37 74 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.935
+ $X2=1.765 $Y2=2.935
r224 36 76 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=2.195 $Y2=2.935
r225 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=1.84 $Y2=2.935
r226 35 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.765 $Y2=1.845
r227 34 75 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.845
r228 34 35 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r229 31 74 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=2.935
r230 31 33 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=4.585
r231 27 73 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.845
r232 27 29 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r233 26 72 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.935
+ $X2=1.335 $Y2=2.935
r234 25 74 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.765 $Y2=2.935
r235 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.41 $Y2=2.935
r236 23 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.765 $Y2=1.845
r237 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.41 $Y2=1.845
r238 20 72 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=2.935
r239 20 22 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=4.585
r240 16 24 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.41 $Y2=1.845
r241 16 99 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.18 $Y2=1.935
r242 16 18 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r243 15 71 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.86
+ $X2=1.18 $Y2=2.935
r244 14 99 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=1.935
r245 14 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=2.86
r246 11 69 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=2.935
r247 11 13 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=4.585
r248 7 97 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.935
r249 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.075
r250 2 87 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r251 2 85 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r252 1 81 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_6%Y 1 2 3 4 5 6 19 20 22 24 26 29 30 31 32
+ 33 34 35 41 47 53 55 67 79
c124 35 0 1.33323e-19 $X=2.84 $Y=2.845
c125 34 0 1.33323e-19 $X=2.84 $Y=1.595
c126 33 0 2.66647e-19 $X=2.125 $Y=2.96
c127 31 0 2.66647e-19 $X=2.125 $Y=1.48
c128 20 0 1.33323e-19 $X=1.12 $Y=2.845
c129 19 0 1.33323e-19 $X=1.12 $Y=1.595
r130 86 88 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r131 74 76 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r132 62 64 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r133 53 86 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=3.455
r134 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=2.96
r135 50 79 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.84 $Y=1.48
+ $X2=2.84 $Y2=0.825
r136 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=1.48
+ $X2=2.84 $Y2=1.48
r137 47 74 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=3.455
r138 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=2.96
r139 44 67 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=0.825
r140 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=1.48
r141 41 62 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=3.455
r142 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=2.96
r143 38 55 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=0.825
r144 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=1.48
r145 35 52 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=2.845
+ $X2=2.84 $Y2=2.96
r146 34 49 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=1.48
r147 34 35 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=2.845
r148 33 46 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=2.96
+ $X2=1.98 $Y2=2.96
r149 32 52 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.84 $Y2=2.96
r150 32 33 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.125 $Y2=2.96
r151 31 43 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=1.48
+ $X2=1.98 $Y2=1.48
r152 30 49 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.84 $Y2=1.48
r153 30 31 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.125 $Y2=1.48
r154 29 46 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.845
+ $X2=1.98 $Y2=2.96
r155 28 43 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=1.48
r156 28 29 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=2.845
r157 27 40 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.96
+ $X2=1.12 $Y2=2.96
r158 26 46 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.98 $Y2=2.96
r159 26 27 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.265 $Y2=2.96
r160 25 37 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1.48
+ $X2=1.12 $Y2=1.48
r161 24 43 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.98 $Y2=1.48
r162 24 25 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.265 $Y2=1.48
r163 20 40 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.96
r164 20 22 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.27
r165 19 37 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=1.48
r166 19 22 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=2.27
r167 6 88 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r168 6 86 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r169 5 76 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r170 5 74 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r171 4 64 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r172 4 62 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r173 3 79 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r174 2 67 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r175 1 55 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
.ends

