* File: sky130_osu_sc_12T_ls__inv_6.pex.spice
* Created: Fri Nov 12 15:38:05 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_LS__INV_6%GND 1 2 3 4 41 45 47 54 56 63 65 73 84 86
r89 84 86 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r90 71 73 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.755
r91 66 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r92 65 71 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.305
r93 61 80 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r94 61 63 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.755
r95 57 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r96 56 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r97 52 79 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r98 52 54 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.755
r99 47 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r100 43 45 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r101 41 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r102 41 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r103 41 43 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r104 41 48 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r105 41 65 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r106 41 66 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r107 41 56 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r108 41 57 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r109 41 47 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r110 41 48 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r111 4 73 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.7 $Y=0.575
+ $X2=2.84 $Y2=0.755
r112 3 63 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.755
r113 2 54 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.755
r114 1 45 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_6%VDD 1 2 3 4 33 37 39 45 49 55 59 66 76 80
r58 76 80 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=2.38 $Y2=4.287
r59 71 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=4.25
+ $X2=0.34 $Y2=4.25
r60 66 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=2.955
+ $X2=2.84 $Y2=3.635
r61 64 69 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.84 $Y=4.135 $X2=2.84
+ $Y2=3.635
r62 62 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=4.25
+ $X2=2.38 $Y2=4.25
r63 60 74 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=1.98 $Y2=4.287
r64 60 62 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=4.287
+ $X2=2.38 $Y2=4.287
r65 59 64 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.84 $Y2=4.135
r66 59 62 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=4.287
+ $X2=2.38 $Y2=4.287
r67 55 58 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=2.955
+ $X2=1.98 $Y2=3.635
r68 53 74 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=4.287
r69 53 58 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.98 $Y=4.135 $X2=1.98
+ $Y2=3.635
r70 50 73 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.12 $Y2=4.287
r71 50 52 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=4.287
+ $X2=1.7 $Y2=4.287
r72 49 74 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.98 $Y2=4.287
r73 49 52 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=4.287
+ $X2=1.7 $Y2=4.287
r74 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=2.955
+ $X2=1.12 $Y2=3.635
r75 43 73 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=4.287
r76 43 48 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.12 $Y=4.135 $X2=1.12
+ $Y2=3.635
r77 40 71 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r78 40 42 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.02 $Y2=4.287
r79 39 73 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.12 $Y2=4.287
r80 39 42 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=4.287
+ $X2=1.02 $Y2=4.287
r81 35 71 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r82 35 37 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135 $X2=0.26
+ $Y2=3.635
r83 33 62 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=4.135 $X2=2.38 $Y2=4.22
r84 33 52 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=4.135 $X2=1.7 $Y2=4.22
r85 33 42 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r86 33 71 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r87 4 69 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=3.635
r88 4 66 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.605 $X2=2.84 $Y2=2.955
r89 3 58 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=3.635
r90 3 55 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.605 $X2=1.98 $Y2=2.955
r91 2 48 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=3.635
r92 2 45 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.605 $X2=1.12 $Y2=2.955
r93 1 37 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_6%A 1 3 7 8 10 11 13 15 17 18 20 21 23 25
+ 27 28 30 31 33 35 37 38 40 41 43 45 47 49 50 52 53 55 57 59 60 62 63 65 66 68
+ 69 70 71 72 73 74 75 76 79 81 83 86
c179 50 0 1.33323e-19 $X=2.195 $Y=2.48
c180 45 0 1.33323e-19 $X=2.195 $Y=1.22
c181 38 0 1.33323e-19 $X=1.765 $Y=2.48
c182 35 0 1.33323e-19 $X=1.765 $Y=1.22
c183 28 0 1.33323e-19 $X=1.335 $Y=2.48
c184 25 0 1.33323e-19 $X=1.335 $Y=1.22
c185 18 0 1.33323e-19 $X=0.905 $Y=2.48
c186 15 0 1.33323e-19 $X=0.905 $Y=1.22
r187 86 89 0.00150602 $w=4.15e-07 $l=5e-09 $layer=MET1_cond $X=0.405 $Y=2.845
+ $X2=0.405 $Y2=2.85
r188 81 83 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.405 $Y=1.825
+ $X2=0.535 $Y2=1.825
r189 79 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r190 77 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.405 $Y2=1.825
r191 77 79 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.32 $Y=1.91
+ $X2=0.32 $Y2=2.85
r192 65 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.825 $X2=0.535 $Y2=1.825
r193 65 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.99
r194 65 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.825
+ $X2=0.535 $Y2=1.66
r195 60 62 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.625 $Y=2.48
+ $X2=2.625 $Y2=3.235
r196 57 59 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.625 $Y=1.22
+ $X2=2.625 $Y2=0.835
r197 56 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.405
+ $X2=2.195 $Y2=2.405
r198 55 60 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.625 $Y2=2.48
r199 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.405
+ $X2=2.27 $Y2=2.405
r200 54 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.295
+ $X2=2.195 $Y2=1.295
r201 53 57 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=1.295
+ $X2=2.625 $Y2=1.22
r202 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.295
+ $X2=2.27 $Y2=1.295
r203 50 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=2.405
r204 50 52 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.195 $Y=2.48
+ $X2=2.195 $Y2=3.235
r205 49 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.33
+ $X2=2.195 $Y2=2.405
r206 48 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.37
+ $X2=2.195 $Y2=1.295
r207 48 49 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.195 $Y=1.37
+ $X2=2.195 $Y2=2.33
r208 45 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.22
+ $X2=2.195 $Y2=1.295
r209 45 47 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.195 $Y=1.22
+ $X2=2.195 $Y2=0.835
r210 44 74 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.405
+ $X2=1.765 $Y2=2.405
r211 43 76 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=2.195 $Y2=2.405
r212 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.405
+ $X2=1.84 $Y2=2.405
r213 42 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.295
+ $X2=1.765 $Y2=1.295
r214 41 75 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.295
+ $X2=2.195 $Y2=1.295
r215 41 42 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.295
+ $X2=1.84 $Y2=1.295
r216 38 74 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=2.405
r217 38 40 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.765 $Y=2.48
+ $X2=1.765 $Y2=3.235
r218 35 73 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.22
+ $X2=1.765 $Y2=1.295
r219 35 37 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.765 $Y=1.22
+ $X2=1.765 $Y2=0.835
r220 34 72 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.405
+ $X2=1.335 $Y2=2.405
r221 33 74 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.765 $Y2=2.405
r222 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.405
+ $X2=1.41 $Y2=2.405
r223 32 71 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.335 $Y2=1.295
r224 31 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.295
+ $X2=1.765 $Y2=1.295
r225 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.295
+ $X2=1.41 $Y2=1.295
r226 28 72 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=2.405
r227 28 30 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.335 $Y=2.48
+ $X2=1.335 $Y2=3.235
r228 25 71 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=1.295
r229 25 27 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.335 $Y=1.22
+ $X2=1.335 $Y2=0.835
r230 24 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=2.405
+ $X2=0.905 $Y2=2.405
r231 23 72 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=1.335 $Y2=2.405
r232 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=2.405
+ $X2=0.98 $Y2=2.405
r233 22 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.295
+ $X2=0.905 $Y2=1.295
r234 21 71 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=1.335 $Y2=1.295
r235 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.26 $Y=1.295
+ $X2=0.98 $Y2=1.295
r236 18 70 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=2.405
r237 18 20 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.905 $Y=2.48
+ $X2=0.905 $Y2=3.235
r238 15 69 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=1.295
r239 15 17 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.905 $Y=1.22
+ $X2=0.905 $Y2=0.835
r240 14 68 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=2.405
+ $X2=0.475 $Y2=2.405
r241 13 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.905 $Y2=2.405
r242 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=2.405
+ $X2=0.55 $Y2=2.405
r243 12 63 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.475 $Y2=1.295
r244 11 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.905 $Y2=1.295
r245 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.83 $Y=1.295
+ $X2=0.55 $Y2=1.295
r246 8 68 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=2.405
r247 8 10 242.607 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.475 $Y=2.48
+ $X2=0.475 $Y2=3.235
r248 7 68 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=2.405
r249 7 67 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.475 $Y=2.33
+ $X2=0.475 $Y2=1.99
r250 4 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.295
r251 4 66 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=1.37
+ $X2=0.475 $Y2=1.66
r252 1 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=1.295
r253 1 3 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=1.22
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_12T_LS__INV_6%Y 1 2 3 7 8 9 26 32 40 46 54 60 67 68 70
+ 72 74 77 78 79 80 81 82 83
c136 83 0 1.33323e-19 $X=2.41 $Y=2.365
c137 82 0 1.33323e-19 $X=2.41 $Y=1.115
c138 81 0 2.66647e-19 $X=1.695 $Y=2.48
c139 79 0 2.66647e-19 $X=1.695 $Y=1
c140 68 0 1.33323e-19 $X=0.69 $Y=2.365
c141 67 0 1.33323e-19 $X=0.69 $Y=1.115
r142 83 95 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.365
+ $X2=2.41 $Y2=2.48
r143 82 93 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=1
r144 82 83 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.41 $Y=1.115
+ $X2=2.41 $Y2=2.365
r145 81 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.48
+ $X2=1.55 $Y2=2.48
r146 80 95 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.48
+ $X2=2.41 $Y2=2.48
r147 80 81 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.48
+ $X2=1.695 $Y2=2.48
r148 79 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1
+ $X2=1.55 $Y2=1
r149 78 93 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=2.41 $Y2=1
r150 78 79 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1
+ $X2=1.695 $Y2=1
r151 77 91 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.365
+ $X2=1.55 $Y2=2.48
r152 76 89 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=1
r153 76 77 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.55 $Y=1.115
+ $X2=1.55 $Y2=2.365
r154 75 87 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=2.48
+ $X2=0.69 $Y2=2.48
r155 74 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=1.55 $Y2=2.48
r156 74 75 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=2.48
+ $X2=0.835 $Y2=2.48
r157 73 85 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1
+ $X2=0.69 $Y2=1
r158 72 89 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=1.55 $Y2=1
r159 72 73 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.405 $Y=1
+ $X2=0.835 $Y2=1
r160 68 87 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=2.48
r161 68 70 0.621059 $w=1.7e-07 $l=6.45e-07 $layer=MET1_cond $X=0.69 $Y=2.365
+ $X2=0.69 $Y2=1.72
r162 67 85 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1
r163 67 70 0.582544 $w=1.7e-07 $l=6.05e-07 $layer=MET1_cond $X=0.69 $Y=1.115
+ $X2=0.69 $Y2=1.72
r164 63 65 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.41 $Y=2.955
+ $X2=2.41 $Y2=3.635
r165 60 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.48
+ $X2=2.41 $Y2=2.48
r166 60 63 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.41 $Y=2.48
+ $X2=2.41 $Y2=2.955
r167 57 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1 $X2=2.41
+ $Y2=1
r168 54 57 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.41 $Y=0.755
+ $X2=2.41 $Y2=1
r169 49 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=2.955
+ $X2=1.55 $Y2=3.635
r170 46 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.48
r171 46 49 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.55 $Y=2.48
+ $X2=1.55 $Y2=2.955
r172 43 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1 $X2=1.55
+ $Y2=1
r173 40 43 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.755
+ $X2=1.55 $Y2=1
r174 35 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.955
+ $X2=0.69 $Y2=3.635
r175 32 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.48
r176 32 35 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.69 $Y=2.48
+ $X2=0.69 $Y2=2.955
r177 29 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1 $X2=0.69
+ $Y2=1
r178 26 29 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0.755
+ $X2=0.69 $Y2=1
r179 9 65 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=3.635
r180 9 63 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.605 $X2=2.41 $Y2=2.955
r181 8 51 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=3.635
r182 8 49 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.605 $X2=1.55 $Y2=2.955
r183 7 37 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.635
r184 7 35 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.955
r185 3 54 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.755
r186 2 40 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.755
r187 1 26 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

