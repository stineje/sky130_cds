* File: sky130_osu_sc_15T_hs__and2_8.pxi.spice
* Created: Fri Nov 12 14:27:15 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__AND2_8%GND N_GND_M1004_d N_GND_M1008_s N_GND_M1013_s
+ N_GND_M1015_s N_GND_M1017_s N_GND_M1007_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p
+ N_GND_c_22_p N_GND_c_30_p N_GND_c_36_p N_GND_c_43_p N_GND_c_50_p N_GND_c_57_p
+ N_GND_c_63_p GND N_GND_c_3_p PM_SKY130_OSU_SC_15T_HS__AND2_8%GND
x_PM_SKY130_OSU_SC_15T_HS__AND2_8%VDD N_VDD_M1010_s N_VDD_M1005_d N_VDD_M1001_d
+ N_VDD_M1006_d N_VDD_M1012_d N_VDD_M1019_d N_VDD_M1010_b N_VDD_c_143_p
+ N_VDD_c_144_p N_VDD_c_155_p N_VDD_c_162_p N_VDD_c_168_p N_VDD_c_174_p
+ N_VDD_c_179_p N_VDD_c_185_p N_VDD_c_190_p N_VDD_c_196_p N_VDD_c_201_p VDD
+ N_VDD_c_145_p PM_SKY130_OSU_SC_15T_HS__AND2_8%VDD
x_PM_SKY130_OSU_SC_15T_HS__AND2_8%A N_A_M1007_g N_A_M1010_g N_A_c_232_n
+ N_A_c_233_n A PM_SKY130_OSU_SC_15T_HS__AND2_8%A
x_PM_SKY130_OSU_SC_15T_HS__AND2_8%B N_B_M1004_g N_B_M1005_g N_B_c_266_n
+ N_B_c_267_n B PM_SKY130_OSU_SC_15T_HS__AND2_8%B
x_PM_SKY130_OSU_SC_15T_HS__AND2_8%A_27_115# N_A_27_115#_M1007_s
+ N_A_27_115#_M1010_d N_A_27_115#_M1003_g N_A_27_115#_c_375_n
+ N_A_27_115#_M1000_g N_A_27_115#_c_306_n N_A_27_115#_c_307_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_380_n N_A_27_115#_M1001_g
+ N_A_27_115#_c_312_n N_A_27_115#_c_314_n N_A_27_115#_c_315_n
+ N_A_27_115#_M1009_g N_A_27_115#_c_387_n N_A_27_115#_M1002_g
+ N_A_27_115#_c_320_n N_A_27_115#_c_321_n N_A_27_115#_M1013_g
+ N_A_27_115#_c_392_n N_A_27_115#_M1006_g N_A_27_115#_c_326_n
+ N_A_27_115#_c_328_n N_A_27_115#_M1014_g N_A_27_115#_c_333_n
+ N_A_27_115#_c_398_n N_A_27_115#_M1011_g N_A_27_115#_c_334_n
+ N_A_27_115#_c_335_n N_A_27_115#_M1015_g N_A_27_115#_c_403_n
+ N_A_27_115#_M1012_g N_A_27_115#_c_340_n N_A_27_115#_c_342_n
+ N_A_27_115#_M1016_g N_A_27_115#_c_409_n N_A_27_115#_M1018_g
+ N_A_27_115#_c_347_n N_A_27_115#_c_348_n N_A_27_115#_M1017_g
+ N_A_27_115#_c_414_n N_A_27_115#_M1019_g N_A_27_115#_c_353_n
+ N_A_27_115#_c_354_n N_A_27_115#_c_355_n N_A_27_115#_c_356_n
+ N_A_27_115#_c_357_n N_A_27_115#_c_358_n N_A_27_115#_c_359_n
+ N_A_27_115#_c_360_n N_A_27_115#_c_361_n N_A_27_115#_c_362_n
+ N_A_27_115#_c_363_n N_A_27_115#_c_364_n N_A_27_115#_c_365_n
+ N_A_27_115#_c_369_n N_A_27_115#_c_370_n N_A_27_115#_c_425_n
+ N_A_27_115#_c_371_n N_A_27_115#_c_373_n N_A_27_115#_c_374_n
+ N_A_27_115#_c_441_n PM_SKY130_OSU_SC_15T_HS__AND2_8%A_27_115#
x_PM_SKY130_OSU_SC_15T_HS__AND2_8%Y N_Y_M1003_d N_Y_M1009_d N_Y_M1014_d
+ N_Y_M1016_d N_Y_M1000_s N_Y_M1002_s N_Y_M1011_s N_Y_M1018_s N_Y_c_545_n
+ N_Y_c_550_n N_Y_c_551_n N_Y_c_556_n N_Y_c_557_n N_Y_c_562_n N_Y_c_563_n
+ N_Y_c_568_n N_Y_c_569_n N_Y_c_572_n Y N_Y_c_574_n N_Y_c_577_n N_Y_c_578_n
+ N_Y_c_579_n N_Y_c_582_n N_Y_c_585_n N_Y_c_586_n N_Y_c_587_n N_Y_c_590_n
+ N_Y_c_591_n N_Y_c_592_n N_Y_c_593_n N_Y_c_596_n N_Y_c_597_n
+ PM_SKY130_OSU_SC_15T_HS__AND2_8%Y
cc_1 N_GND_M1007_b N_A_M1007_g 0.0859626f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.895
cc_2 N_GND_c_2_p N_A_M1007_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.895
cc_3 N_GND_c_3_p N_A_M1007_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.475 $Y2=0.895
cc_4 N_GND_M1007_b N_A_c_232_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.505
cc_5 N_GND_M1007_b N_A_c_233_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.505
cc_6 N_GND_M1007_b N_B_M1004_g 0.0514444f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.895
cc_7 N_GND_c_2_p N_B_M1004_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.895
cc_8 N_GND_c_8_p N_B_M1004_g 0.00487132f $X=1.05 $Y=0.9 $X2=0.835 $Y2=0.895
cc_9 N_GND_c_3_p N_B_M1004_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.835 $Y2=0.895
cc_10 N_GND_M1007_b N_B_M1005_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.825
cc_11 N_GND_M1007_b N_B_c_266_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.165
cc_12 N_GND_M1007_b N_B_c_267_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.165
cc_13 N_GND_M1007_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.7
cc_14 N_GND_M1007_b N_A_27_115#_M1003_g 0.0266646f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.895
cc_15 N_GND_c_8_p N_A_27_115#_M1003_g 0.00883341f $X=1.05 $Y=0.9 $X2=1.335
+ $Y2=0.895
cc_16 N_GND_c_16_p N_A_27_115#_M1003_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.895
cc_17 N_GND_c_3_p N_A_27_115#_M1003_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.335
+ $Y2=0.895
cc_18 N_GND_M1007_b N_A_27_115#_c_306_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.55
cc_19 N_GND_M1007_b N_A_27_115#_c_307_n 0.00727817f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.625
cc_20 N_GND_M1007_b N_A_27_115#_M1008_g 0.0245311f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.895
cc_21 N_GND_c_16_p N_A_27_115#_M1008_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.895
cc_22 N_GND_c_22_p N_A_27_115#_M1008_g 0.00443715f $X=1.98 $Y=0.9 $X2=1.765
+ $Y2=0.895
cc_23 N_GND_c_3_p N_A_27_115#_M1008_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.765
+ $Y2=0.895
cc_24 N_GND_M1007_b N_A_27_115#_c_312_n 0.0179436f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.585
cc_25 N_GND_c_22_p N_A_27_115#_c_312_n 0.00291042f $X=1.98 $Y=0.9 $X2=2.12
+ $Y2=1.585
cc_26 N_GND_M1007_b N_A_27_115#_c_314_n 0.0456099f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.585
cc_27 N_GND_M1007_b N_A_27_115#_c_315_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.625
cc_28 N_GND_M1007_b N_A_27_115#_M1009_g 0.0245289f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.895
cc_29 N_GND_c_22_p N_A_27_115#_M1009_g 0.00443715f $X=1.98 $Y=0.9 $X2=2.195
+ $Y2=0.895
cc_30 N_GND_c_30_p N_A_27_115#_M1009_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.895
cc_31 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=4.42 $Y=0.19 $X2=2.195
+ $Y2=0.895
cc_32 N_GND_M1007_b N_A_27_115#_c_320_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.585
cc_33 N_GND_M1007_b N_A_27_115#_c_321_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.625
cc_34 N_GND_M1007_b N_A_27_115#_M1013_g 0.0245289f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.895
cc_35 N_GND_c_30_p N_A_27_115#_M1013_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.895
cc_36 N_GND_c_36_p N_A_27_115#_M1013_g 0.00443715f $X=2.84 $Y=0.9 $X2=2.625
+ $Y2=0.895
cc_37 N_GND_c_3_p N_A_27_115#_M1013_g 0.00468827f $X=4.42 $Y=0.19 $X2=2.625
+ $Y2=0.895
cc_38 N_GND_M1007_b N_A_27_115#_c_326_n 0.0179436f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.585
cc_39 N_GND_c_36_p N_A_27_115#_c_326_n 0.00291042f $X=2.84 $Y=0.9 $X2=2.98
+ $Y2=1.585
cc_40 N_GND_M1007_b N_A_27_115#_c_328_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.625
cc_41 N_GND_M1007_b N_A_27_115#_M1014_g 0.0245289f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=0.895
cc_42 N_GND_c_36_p N_A_27_115#_M1014_g 0.00443715f $X=2.84 $Y=0.9 $X2=3.055
+ $Y2=0.895
cc_43 N_GND_c_43_p N_A_27_115#_M1014_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.055
+ $Y2=0.895
cc_44 N_GND_c_3_p N_A_27_115#_M1014_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.055
+ $Y2=0.895
cc_45 N_GND_M1007_b N_A_27_115#_c_333_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.55
cc_46 N_GND_M1007_b N_A_27_115#_c_334_n 0.0180386f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.585
cc_47 N_GND_M1007_b N_A_27_115#_c_335_n 0.0118833f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.625
cc_48 N_GND_M1007_b N_A_27_115#_M1015_g 0.0245289f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=0.895
cc_49 N_GND_c_43_p N_A_27_115#_M1015_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.485
+ $Y2=0.895
cc_50 N_GND_c_50_p N_A_27_115#_M1015_g 0.00443715f $X=3.7 $Y=0.9 $X2=3.485
+ $Y2=0.895
cc_51 N_GND_c_3_p N_A_27_115#_M1015_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.485
+ $Y2=0.895
cc_52 N_GND_M1007_b N_A_27_115#_c_340_n 0.0179436f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.585
cc_53 N_GND_c_50_p N_A_27_115#_c_340_n 0.00291042f $X=3.7 $Y=0.9 $X2=3.84
+ $Y2=1.585
cc_54 N_GND_M1007_b N_A_27_115#_c_342_n 0.013058f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.625
cc_55 N_GND_M1007_b N_A_27_115#_M1016_g 0.0245289f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=0.895
cc_56 N_GND_c_50_p N_A_27_115#_M1016_g 0.00443715f $X=3.7 $Y=0.9 $X2=3.915
+ $Y2=0.895
cc_57 N_GND_c_57_p N_A_27_115#_M1016_g 0.00606474f $X=4.475 $Y=0.152 $X2=3.915
+ $Y2=0.895
cc_58 N_GND_c_3_p N_A_27_115#_M1016_g 0.00468827f $X=4.42 $Y=0.19 $X2=3.915
+ $Y2=0.895
cc_59 N_GND_M1007_b N_A_27_115#_c_347_n 0.0369419f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=1.585
cc_60 N_GND_M1007_b N_A_27_115#_c_348_n 0.0268552f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=2.625
cc_61 N_GND_M1007_b N_A_27_115#_M1017_g 0.0333625f $X=-0.045 $Y=0 $X2=4.345
+ $Y2=0.895
cc_62 N_GND_c_57_p N_A_27_115#_M1017_g 0.00606474f $X=4.475 $Y=0.152 $X2=4.345
+ $Y2=0.895
cc_63 N_GND_c_63_p N_A_27_115#_M1017_g 0.0105074f $X=4.56 $Y=0.9 $X2=4.345
+ $Y2=0.895
cc_64 N_GND_c_3_p N_A_27_115#_M1017_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.345
+ $Y2=0.895
cc_65 N_GND_M1007_b N_A_27_115#_c_353_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.625
cc_66 N_GND_M1007_b N_A_27_115#_c_354_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.625
cc_67 N_GND_M1007_b N_A_27_115#_c_355_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.585
cc_68 N_GND_M1007_b N_A_27_115#_c_356_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.625
cc_69 N_GND_M1007_b N_A_27_115#_c_357_n 0.00873941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.585
cc_70 N_GND_M1007_b N_A_27_115#_c_358_n 0.00735657f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.625
cc_71 N_GND_M1007_b N_A_27_115#_c_359_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.585
cc_72 N_GND_M1007_b N_A_27_115#_c_360_n 0.00151234f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.625
cc_73 N_GND_M1007_b N_A_27_115#_c_361_n 0.00873941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.585
cc_74 N_GND_M1007_b N_A_27_115#_c_362_n 0.00735657f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.625
cc_75 N_GND_M1007_b N_A_27_115#_c_363_n 0.00873941f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=1.585
cc_76 N_GND_M1007_b N_A_27_115#_c_364_n 0.00735657f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=2.625
cc_77 N_GND_M1007_b N_A_27_115#_c_365_n 0.0193081f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.9
cc_78 N_GND_c_2_p N_A_27_115#_c_365_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.9
cc_79 N_GND_c_8_p N_A_27_115#_c_365_n 8.71428e-19 $X=1.05 $Y=0.9 $X2=0.26
+ $Y2=0.9
cc_80 N_GND_c_3_p N_A_27_115#_c_365_n 0.00476261f $X=4.42 $Y=0.19 $X2=0.26
+ $Y2=0.9
cc_81 N_GND_M1007_b N_A_27_115#_c_369_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.675
cc_82 N_GND_M1007_b N_A_27_115#_c_370_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.675
cc_83 N_GND_M1007_b N_A_27_115#_c_371_n 0.0227928f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.675
cc_84 N_GND_c_8_p N_A_27_115#_c_371_n 0.00867832f $X=1.05 $Y=0.9 $X2=1.43
+ $Y2=1.675
cc_85 N_GND_M1007_b N_A_27_115#_c_373_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.675
cc_86 N_GND_M1007_b N_A_27_115#_c_374_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.305
cc_87 N_GND_M1007_b N_Y_c_545_n 0.00515424f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.9
cc_88 N_GND_c_8_p N_Y_c_545_n 0.0153376f $X=1.05 $Y=0.9 $X2=1.55 $Y2=0.9
cc_89 N_GND_c_16_p N_Y_c_545_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.9
cc_90 N_GND_c_22_p N_Y_c_545_n 0.00358291f $X=1.98 $Y=0.9 $X2=1.55 $Y2=0.9
cc_91 N_GND_c_3_p N_Y_c_545_n 0.00475776f $X=4.42 $Y=0.19 $X2=1.55 $Y2=0.9
cc_92 N_GND_M1007_b N_Y_c_550_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.33
cc_93 N_GND_M1007_b N_Y_c_551_n 0.00610793f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.9
cc_94 N_GND_c_22_p N_Y_c_551_n 0.00358291f $X=1.98 $Y=0.9 $X2=2.41 $Y2=0.9
cc_95 N_GND_c_30_p N_Y_c_551_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.9
cc_96 N_GND_c_36_p N_Y_c_551_n 0.00358291f $X=2.84 $Y=0.9 $X2=2.41 $Y2=0.9
cc_97 N_GND_c_3_p N_Y_c_551_n 0.00475776f $X=4.42 $Y=0.19 $X2=2.41 $Y2=0.9
cc_98 N_GND_M1007_b N_Y_c_556_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.33
cc_99 N_GND_M1007_b N_Y_c_557_n 0.00610793f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.9
cc_100 N_GND_c_36_p N_Y_c_557_n 0.00358291f $X=2.84 $Y=0.9 $X2=3.27 $Y2=0.9
cc_101 N_GND_c_43_p N_Y_c_557_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.9
cc_102 N_GND_c_50_p N_Y_c_557_n 0.00358291f $X=3.7 $Y=0.9 $X2=3.27 $Y2=0.9
cc_103 N_GND_c_3_p N_Y_c_557_n 0.00475776f $X=4.42 $Y=0.19 $X2=3.27 $Y2=0.9
cc_104 N_GND_M1007_b N_Y_c_562_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.33
cc_105 N_GND_M1007_b N_Y_c_563_n 0.00610793f $X=-0.045 $Y=0 $X2=4.13 $Y2=0.9
cc_106 N_GND_c_50_p N_Y_c_563_n 0.00358291f $X=3.7 $Y=0.9 $X2=4.13 $Y2=0.9
cc_107 N_GND_c_57_p N_Y_c_563_n 0.0075556f $X=4.475 $Y=0.152 $X2=4.13 $Y2=0.9
cc_108 N_GND_c_63_p N_Y_c_563_n 0.00251593f $X=4.56 $Y=0.9 $X2=4.13 $Y2=0.9
cc_109 N_GND_c_3_p N_Y_c_563_n 0.00475776f $X=4.42 $Y=0.19 $X2=4.13 $Y2=0.9
cc_110 N_GND_M1007_b N_Y_c_568_n 0.0152877f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.33
cc_111 N_GND_M1007_b N_Y_c_569_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.335
cc_112 N_GND_c_8_p N_Y_c_569_n 0.00377613f $X=1.05 $Y=0.9 $X2=1.55 $Y2=1.335
cc_113 N_GND_c_22_p N_Y_c_569_n 7.53951e-19 $X=1.98 $Y=0.9 $X2=1.55 $Y2=1.335
cc_114 N_GND_M1007_b N_Y_c_572_n 0.00509006f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.215
cc_115 N_GND_M1007_b Y 0.0306813f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.96
cc_116 N_GND_M1008_s N_Y_c_574_n 0.00418405f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.22
cc_117 N_GND_M1007_b N_Y_c_574_n 0.00793787f $X=-0.045 $Y=0 $X2=2.265 $Y2=1.22
cc_118 N_GND_c_22_p N_Y_c_574_n 0.0179014f $X=1.98 $Y=0.9 $X2=2.265 $Y2=1.22
cc_119 N_GND_M1007_b N_Y_c_577_n 0.0188475f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.33
cc_120 N_GND_M1007_b N_Y_c_578_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.215
cc_121 N_GND_M1013_s N_Y_c_579_n 0.00418405f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.22
cc_122 N_GND_M1007_b N_Y_c_579_n 0.00793787f $X=-0.045 $Y=0 $X2=3.125 $Y2=1.22
cc_123 N_GND_c_36_p N_Y_c_579_n 0.0179014f $X=2.84 $Y=0.9 $X2=3.125 $Y2=1.22
cc_124 N_GND_M1007_b N_Y_c_582_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.22
cc_125 N_GND_c_22_p N_Y_c_582_n 7.53951e-19 $X=1.98 $Y=0.9 $X2=2.555 $Y2=1.22
cc_126 N_GND_c_36_p N_Y_c_582_n 7.53951e-19 $X=2.84 $Y=0.9 $X2=2.555 $Y2=1.22
cc_127 N_GND_M1007_b N_Y_c_585_n 0.0144616f $X=-0.045 $Y=0 $X2=3.125 $Y2=2.33
cc_128 N_GND_M1007_b N_Y_c_586_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.33
cc_129 N_GND_M1007_b N_Y_c_587_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.335
cc_130 N_GND_c_36_p N_Y_c_587_n 7.53951e-19 $X=2.84 $Y=0.9 $X2=3.27 $Y2=1.335
cc_131 N_GND_c_50_p N_Y_c_587_n 0.00113348f $X=3.7 $Y=0.9 $X2=3.27 $Y2=1.335
cc_132 N_GND_M1007_b N_Y_c_590_n 0.0358528f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.215
cc_133 N_GND_M1007_b N_Y_c_591_n 0.0188475f $X=-0.045 $Y=0 $X2=3.985 $Y2=2.33
cc_134 N_GND_M1007_b N_Y_c_592_n 0.00584404f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.33
cc_135 N_GND_M1007_b N_Y_c_593_n 0.00409378f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.335
cc_136 N_GND_c_50_p N_Y_c_593_n 7.53951e-19 $X=3.7 $Y=0.9 $X2=4.13 $Y2=1.335
cc_137 N_GND_c_63_p N_Y_c_593_n 0.00402079f $X=4.56 $Y=0.9 $X2=4.13 $Y2=1.335
cc_138 N_GND_M1007_b N_Y_c_596_n 0.06145f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.215
cc_139 N_GND_M1015_s N_Y_c_597_n 0.00418405f $X=3.56 $Y=0.575 $X2=4.13 $Y2=1.22
cc_140 N_GND_M1007_b N_Y_c_597_n 0.00793787f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.22
cc_141 N_GND_c_50_p N_Y_c_597_n 0.0169856f $X=3.7 $Y=0.9 $X2=4.13 $Y2=1.22
cc_142 N_VDD_M1010_b N_A_M1010_g 0.0193382f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_143 N_VDD_c_143_p N_A_M1010_g 0.00713292f $X=0.26 $Y=3.895 $X2=0.475
+ $Y2=3.825
cc_144 N_VDD_c_144_p N_A_M1010_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_145 N_VDD_c_145_p N_A_M1010_g 0.00429146f $X=4.42 $Y=5.36 $X2=0.475 $Y2=3.825
cc_146 N_VDD_M1010_b N_A_c_232_n 0.0111025f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=2.505
cc_147 N_VDD_M1010_s N_A_c_233_n 0.0127742f $X=0.135 $Y=2.825 $X2=0.27 $Y2=2.505
cc_148 N_VDD_M1010_b N_A_c_233_n 0.00612103f $X=-0.045 $Y=2.645 $X2=0.27
+ $Y2=2.505
cc_149 N_VDD_c_143_p N_A_c_233_n 0.00352433f $X=0.26 $Y=3.895 $X2=0.27 $Y2=2.505
cc_150 N_VDD_M1010_s A 0.00746694f $X=0.135 $Y=2.825 $X2=0.275 $Y2=3.07
cc_151 N_VDD_M1010_b A 0.00970321f $X=-0.045 $Y=2.645 $X2=0.275 $Y2=3.07
cc_152 N_VDD_c_143_p A 0.00428937f $X=0.26 $Y=3.895 $X2=0.275 $Y2=3.07
cc_153 N_VDD_M1010_b N_B_M1005_g 0.0191387f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=3.825
cc_154 N_VDD_c_144_p N_B_M1005_g 0.00496961f $X=1.035 $Y=5.397 $X2=0.905
+ $Y2=3.825
cc_155 N_VDD_c_155_p N_B_M1005_g 0.00354579f $X=1.12 $Y=3.555 $X2=0.905
+ $Y2=3.825
cc_156 N_VDD_c_145_p N_B_M1005_g 0.00429146f $X=4.42 $Y=5.36 $X2=0.905 $Y2=3.825
cc_157 N_VDD_M1010_b N_B_c_267_n 0.00170274f $X=-0.045 $Y=2.645 $X2=0.95
+ $Y2=2.165
cc_158 N_VDD_M1010_b B 0.00860092f $X=-0.045 $Y=2.645 $X2=0.955 $Y2=2.7
cc_159 N_VDD_c_155_p B 0.00236322f $X=1.12 $Y=3.555 $X2=0.955 $Y2=2.7
cc_160 N_VDD_M1010_b N_A_27_115#_c_375_n 0.0174951f $X=-0.045 $Y=2.645 $X2=1.335
+ $Y2=2.7
cc_161 N_VDD_c_155_p N_A_27_115#_c_375_n 0.00354579f $X=1.12 $Y=3.555 $X2=1.335
+ $Y2=2.7
cc_162 N_VDD_c_162_p N_A_27_115#_c_375_n 0.00496961f $X=1.895 $Y=5.397 $X2=1.335
+ $Y2=2.7
cc_163 N_VDD_c_145_p N_A_27_115#_c_375_n 0.00429146f $X=4.42 $Y=5.36 $X2=1.335
+ $Y2=2.7
cc_164 N_VDD_M1010_b N_A_27_115#_c_307_n 0.00427883f $X=-0.045 $Y=2.645 $X2=1.69
+ $Y2=2.625
cc_165 N_VDD_M1010_b N_A_27_115#_c_380_n 0.0173909f $X=-0.045 $Y=2.645 $X2=1.765
+ $Y2=2.7
cc_166 N_VDD_c_155_p N_A_27_115#_c_380_n 3.67508e-19 $X=1.12 $Y=3.555 $X2=1.765
+ $Y2=2.7
cc_167 N_VDD_c_162_p N_A_27_115#_c_380_n 0.00500229f $X=1.895 $Y=5.397 $X2=1.765
+ $Y2=2.7
cc_168 N_VDD_c_168_p N_A_27_115#_c_380_n 0.00373985f $X=1.98 $Y=3.215 $X2=1.765
+ $Y2=2.7
cc_169 N_VDD_c_145_p N_A_27_115#_c_380_n 0.00430409f $X=4.42 $Y=5.36 $X2=1.765
+ $Y2=2.7
cc_170 N_VDD_M1010_b N_A_27_115#_c_315_n 0.00399373f $X=-0.045 $Y=2.645 $X2=2.12
+ $Y2=2.625
cc_171 N_VDD_c_168_p N_A_27_115#_c_315_n 0.0037128f $X=1.98 $Y=3.215 $X2=2.12
+ $Y2=2.625
cc_172 N_VDD_M1010_b N_A_27_115#_c_387_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.195
+ $Y2=2.7
cc_173 N_VDD_c_168_p N_A_27_115#_c_387_n 0.00354579f $X=1.98 $Y=3.215 $X2=2.195
+ $Y2=2.7
cc_174 N_VDD_c_174_p N_A_27_115#_c_387_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.195
+ $Y2=2.7
cc_175 N_VDD_c_145_p N_A_27_115#_c_387_n 0.00429146f $X=4.42 $Y=5.36 $X2=2.195
+ $Y2=2.7
cc_176 N_VDD_M1010_b N_A_27_115#_c_321_n 0.00448664f $X=-0.045 $Y=2.645 $X2=2.55
+ $Y2=2.625
cc_177 N_VDD_M1010_b N_A_27_115#_c_392_n 0.0170809f $X=-0.045 $Y=2.645 $X2=2.625
+ $Y2=2.7
cc_178 N_VDD_c_174_p N_A_27_115#_c_392_n 0.00496961f $X=2.755 $Y=5.397 $X2=2.625
+ $Y2=2.7
cc_179 N_VDD_c_179_p N_A_27_115#_c_392_n 0.00354579f $X=2.84 $Y=3.215 $X2=2.625
+ $Y2=2.7
cc_180 N_VDD_c_145_p N_A_27_115#_c_392_n 0.00429146f $X=4.42 $Y=5.36 $X2=2.625
+ $Y2=2.7
cc_181 N_VDD_M1010_b N_A_27_115#_c_328_n 0.00399373f $X=-0.045 $Y=2.645 $X2=2.98
+ $Y2=2.625
cc_182 N_VDD_c_179_p N_A_27_115#_c_328_n 0.0037128f $X=2.84 $Y=3.215 $X2=2.98
+ $Y2=2.625
cc_183 N_VDD_M1010_b N_A_27_115#_c_398_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.055
+ $Y2=2.7
cc_184 N_VDD_c_179_p N_A_27_115#_c_398_n 0.00354579f $X=2.84 $Y=3.215 $X2=3.055
+ $Y2=2.7
cc_185 N_VDD_c_185_p N_A_27_115#_c_398_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.055
+ $Y2=2.7
cc_186 N_VDD_c_145_p N_A_27_115#_c_398_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.055
+ $Y2=2.7
cc_187 N_VDD_M1010_b N_A_27_115#_c_335_n 0.00448664f $X=-0.045 $Y=2.645 $X2=3.41
+ $Y2=2.625
cc_188 N_VDD_M1010_b N_A_27_115#_c_403_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.485
+ $Y2=2.7
cc_189 N_VDD_c_185_p N_A_27_115#_c_403_n 0.00496961f $X=3.615 $Y=5.397 $X2=3.485
+ $Y2=2.7
cc_190 N_VDD_c_190_p N_A_27_115#_c_403_n 0.00354579f $X=3.7 $Y=3.215 $X2=3.485
+ $Y2=2.7
cc_191 N_VDD_c_145_p N_A_27_115#_c_403_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.485
+ $Y2=2.7
cc_192 N_VDD_M1010_b N_A_27_115#_c_342_n 0.00399373f $X=-0.045 $Y=2.645 $X2=3.84
+ $Y2=2.625
cc_193 N_VDD_c_190_p N_A_27_115#_c_342_n 0.0037128f $X=3.7 $Y=3.215 $X2=3.84
+ $Y2=2.625
cc_194 N_VDD_M1010_b N_A_27_115#_c_409_n 0.0170809f $X=-0.045 $Y=2.645 $X2=3.915
+ $Y2=2.7
cc_195 N_VDD_c_190_p N_A_27_115#_c_409_n 0.00354579f $X=3.7 $Y=3.215 $X2=3.915
+ $Y2=2.7
cc_196 N_VDD_c_196_p N_A_27_115#_c_409_n 0.00496961f $X=4.475 $Y=5.397 $X2=3.915
+ $Y2=2.7
cc_197 N_VDD_c_145_p N_A_27_115#_c_409_n 0.00429146f $X=4.42 $Y=5.36 $X2=3.915
+ $Y2=2.7
cc_198 N_VDD_M1010_b N_A_27_115#_c_348_n 0.00840215f $X=-0.045 $Y=2.645 $X2=4.27
+ $Y2=2.625
cc_199 N_VDD_M1010_b N_A_27_115#_c_414_n 0.0212947f $X=-0.045 $Y=2.645 $X2=4.345
+ $Y2=2.7
cc_200 N_VDD_c_196_p N_A_27_115#_c_414_n 0.00496961f $X=4.475 $Y=5.397 $X2=4.345
+ $Y2=2.7
cc_201 N_VDD_c_201_p N_A_27_115#_c_414_n 0.00713292f $X=4.56 $Y=3.215 $X2=4.345
+ $Y2=2.7
cc_202 N_VDD_c_145_p N_A_27_115#_c_414_n 0.00429146f $X=4.42 $Y=5.36 $X2=4.345
+ $Y2=2.7
cc_203 N_VDD_M1010_b N_A_27_115#_c_353_n 0.0021704f $X=-0.045 $Y=2.645 $X2=1.352
+ $Y2=2.625
cc_204 N_VDD_M1010_b N_A_27_115#_c_354_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=1.765 $Y2=2.625
cc_205 N_VDD_M1010_b N_A_27_115#_c_356_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.195 $Y2=2.625
cc_206 N_VDD_M1010_b N_A_27_115#_c_358_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=2.625 $Y2=2.625
cc_207 N_VDD_M1010_b N_A_27_115#_c_360_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.055 $Y2=2.625
cc_208 N_VDD_M1010_b N_A_27_115#_c_362_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.485 $Y2=2.625
cc_209 N_VDD_M1010_b N_A_27_115#_c_364_n 8.75564e-19 $X=-0.045 $Y=2.645
+ $X2=3.915 $Y2=2.625
cc_210 N_VDD_M1010_b N_A_27_115#_c_425_n 0.00198641f $X=-0.045 $Y=2.645 $X2=0.69
+ $Y2=3.555
cc_211 N_VDD_c_144_p N_A_27_115#_c_425_n 0.00475585f $X=1.035 $Y=5.397 $X2=0.69
+ $Y2=3.555
cc_212 N_VDD_c_145_p N_A_27_115#_c_425_n 0.00434939f $X=4.42 $Y=5.36 $X2=0.69
+ $Y2=3.555
cc_213 N_VDD_M1010_b N_A_27_115#_c_374_n 8.22047e-19 $X=-0.045 $Y=2.645 $X2=0.65
+ $Y2=3.305
cc_214 N_VDD_M1010_b N_Y_c_550_n 0.00388477f $X=-0.045 $Y=2.645 $X2=1.55
+ $Y2=2.33
cc_215 N_VDD_c_162_p N_Y_c_550_n 0.00455459f $X=1.895 $Y=5.397 $X2=1.55 $Y2=2.33
cc_216 N_VDD_c_145_p N_Y_c_550_n 0.00434939f $X=4.42 $Y=5.36 $X2=1.55 $Y2=2.33
cc_217 N_VDD_M1010_b N_Y_c_556_n 0.0042387f $X=-0.045 $Y=2.645 $X2=2.41 $Y2=2.33
cc_218 N_VDD_c_174_p N_Y_c_556_n 0.0045126f $X=2.755 $Y=5.397 $X2=2.41 $Y2=2.33
cc_219 N_VDD_c_145_p N_Y_c_556_n 0.00434939f $X=4.42 $Y=5.36 $X2=2.41 $Y2=2.33
cc_220 N_VDD_M1010_b N_Y_c_562_n 0.0042387f $X=-0.045 $Y=2.645 $X2=3.27 $Y2=2.33
cc_221 N_VDD_c_185_p N_Y_c_562_n 0.00464147f $X=3.615 $Y=5.397 $X2=3.27 $Y2=2.33
cc_222 N_VDD_c_145_p N_Y_c_562_n 0.00434939f $X=4.42 $Y=5.36 $X2=3.27 $Y2=2.33
cc_223 N_VDD_M1010_b N_Y_c_568_n 0.0042387f $X=-0.045 $Y=2.645 $X2=4.13 $Y2=2.33
cc_224 N_VDD_c_196_p N_Y_c_568_n 0.00475585f $X=4.475 $Y=5.397 $X2=4.13 $Y2=2.33
cc_225 N_VDD_c_145_p N_Y_c_568_n 0.00434939f $X=4.42 $Y=5.36 $X2=4.13 $Y2=2.33
cc_226 N_VDD_c_168_p N_Y_c_577_n 0.00622932f $X=1.98 $Y=3.215 $X2=2.265 $Y2=2.33
cc_227 N_VDD_c_179_p N_Y_c_585_n 0.00622932f $X=2.84 $Y=3.215 $X2=3.125 $Y2=2.33
cc_228 N_VDD_c_190_p N_Y_c_591_n 0.00622932f $X=3.7 $Y=3.215 $X2=3.985 $Y2=2.33
cc_229 N_A_M1007_g N_B_M1004_g 0.113664f $X=0.475 $Y=0.895 $X2=0.835 $Y2=0.895
cc_230 N_A_M1007_g N_B_M1005_g 0.0506107f $X=0.475 $Y=0.895 $X2=0.905 $Y2=3.825
cc_231 N_A_M1007_g N_B_c_267_n 7.8234e-19 $X=0.475 $Y=0.895 $X2=0.95 $Y2=2.165
cc_232 N_A_M1007_g N_A_27_115#_c_365_n 0.0189753f $X=0.475 $Y=0.895 $X2=0.26
+ $Y2=0.9
cc_233 N_A_M1007_g N_A_27_115#_c_369_n 0.0160984f $X=0.475 $Y=0.895 $X2=0.525
+ $Y2=1.675
cc_234 N_A_c_232_n N_A_27_115#_c_369_n 0.00117122f $X=0.475 $Y=2.505 $X2=0.525
+ $Y2=1.675
cc_235 N_A_c_233_n N_A_27_115#_c_369_n 2.65873e-19 $X=0.27 $Y=2.505 $X2=0.525
+ $Y2=1.675
cc_236 N_A_c_232_n N_A_27_115#_c_370_n 0.00133457f $X=0.475 $Y=2.505 $X2=0.345
+ $Y2=1.675
cc_237 N_A_c_233_n N_A_27_115#_c_370_n 0.0055861f $X=0.27 $Y=2.505 $X2=0.345
+ $Y2=1.675
cc_238 N_A_M1007_g N_A_27_115#_c_373_n 0.00322084f $X=0.475 $Y=0.895 $X2=0.61
+ $Y2=1.675
cc_239 N_A_M1007_g N_A_27_115#_c_374_n 0.0265302f $X=0.475 $Y=0.895 $X2=0.65
+ $Y2=3.305
cc_240 N_A_M1010_g N_A_27_115#_c_374_n 0.0149699f $X=0.475 $Y=3.825 $X2=0.65
+ $Y2=3.305
cc_241 N_A_c_232_n N_A_27_115#_c_374_n 0.00766302f $X=0.475 $Y=2.505 $X2=0.65
+ $Y2=3.305
cc_242 N_A_c_233_n N_A_27_115#_c_374_n 0.0456533f $X=0.27 $Y=2.505 $X2=0.65
+ $Y2=3.305
cc_243 A N_A_27_115#_c_374_n 0.00758489f $X=0.275 $Y=3.07 $X2=0.65 $Y2=3.305
cc_244 N_A_M1010_g N_A_27_115#_c_441_n 0.00884152f $X=0.475 $Y=3.825 $X2=0.65
+ $Y2=3.475
cc_245 N_B_M1004_g N_A_27_115#_M1003_g 0.0316307f $X=0.835 $Y=0.895 $X2=1.335
+ $Y2=0.895
cc_246 N_B_M1005_g N_A_27_115#_c_306_n 0.00773101f $X=0.905 $Y=3.825 $X2=1.37
+ $Y2=2.55
cc_247 N_B_c_266_n N_A_27_115#_c_306_n 0.0206104f $X=0.95 $Y=2.165 $X2=1.37
+ $Y2=2.55
cc_248 N_B_c_267_n N_A_27_115#_c_306_n 0.0033451f $X=0.95 $Y=2.165 $X2=1.37
+ $Y2=2.55
cc_249 N_B_M1004_g N_A_27_115#_c_314_n 0.0104742f $X=0.835 $Y=0.895 $X2=1.84
+ $Y2=1.585
cc_250 N_B_M1005_g N_A_27_115#_c_353_n 0.0410292f $X=0.905 $Y=3.825 $X2=1.352
+ $Y2=2.625
cc_251 N_B_c_267_n N_A_27_115#_c_353_n 0.00173699f $X=0.95 $Y=2.165 $X2=1.352
+ $Y2=2.625
cc_252 B N_A_27_115#_c_353_n 0.00389258f $X=0.955 $Y=2.7 $X2=1.352 $Y2=2.625
cc_253 N_B_M1004_g N_A_27_115#_c_371_n 0.0182215f $X=0.835 $Y=0.895 $X2=1.43
+ $Y2=1.675
cc_254 N_B_c_266_n N_A_27_115#_c_371_n 0.00258465f $X=0.95 $Y=2.165 $X2=1.43
+ $Y2=1.675
cc_255 N_B_c_267_n N_A_27_115#_c_371_n 0.0101796f $X=0.95 $Y=2.165 $X2=1.43
+ $Y2=1.675
cc_256 N_B_M1004_g N_A_27_115#_c_374_n 0.00755919f $X=0.835 $Y=0.895 $X2=0.65
+ $Y2=3.305
cc_257 N_B_M1005_g N_A_27_115#_c_374_n 0.0137515f $X=0.905 $Y=3.825 $X2=0.65
+ $Y2=3.305
cc_258 N_B_c_267_n N_A_27_115#_c_374_n 0.0541375f $X=0.95 $Y=2.165 $X2=0.65
+ $Y2=3.305
cc_259 B N_A_27_115#_c_374_n 0.00866797f $X=0.955 $Y=2.7 $X2=0.65 $Y2=3.305
cc_260 B N_A_27_115#_c_441_n 0.00281588f $X=0.955 $Y=2.7 $X2=0.65 $Y2=3.475
cc_261 N_B_c_267_n N_Y_c_550_n 0.0149875f $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.33
cc_262 B N_Y_c_550_n 0.00649253f $X=0.955 $Y=2.7 $X2=1.55 $Y2=2.33
cc_263 N_B_M1004_g N_Y_c_569_n 4.07255e-19 $X=0.835 $Y=0.895 $X2=1.55 $Y2=1.335
cc_264 N_B_c_266_n N_Y_c_572_n 5.85867e-19 $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.215
cc_265 N_B_c_267_n N_Y_c_572_n 0.00592261f $X=0.95 $Y=2.165 $X2=1.55 $Y2=2.215
cc_266 N_B_M1004_g Y 6.71108e-19 $X=0.835 $Y=0.895 $X2=1.555 $Y2=1.96
cc_267 N_B_c_267_n Y 0.00695761f $X=0.95 $Y=2.165 $X2=1.555 $Y2=1.96
cc_268 N_A_27_115#_M1003_g N_Y_c_545_n 0.00267571f $X=1.335 $Y=0.895 $X2=1.55
+ $Y2=0.9
cc_269 N_A_27_115#_M1008_g N_Y_c_545_n 0.00260839f $X=1.765 $Y=0.895 $X2=1.55
+ $Y2=0.9
cc_270 N_A_27_115#_c_314_n N_Y_c_545_n 0.00171364f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=0.9
cc_271 N_A_27_115#_c_371_n N_Y_c_545_n 0.00520269f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=0.9
cc_272 N_A_27_115#_c_375_n N_Y_c_550_n 0.00287202f $X=1.335 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_273 N_A_27_115#_c_306_n N_Y_c_550_n 0.00744772f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.33
cc_274 N_A_27_115#_c_307_n N_Y_c_550_n 0.0156184f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.33
cc_275 N_A_27_115#_c_380_n N_Y_c_550_n 0.00401146f $X=1.765 $Y=2.7 $X2=1.55
+ $Y2=2.33
cc_276 N_A_27_115#_c_314_n N_Y_c_550_n 0.00182797f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.33
cc_277 N_A_27_115#_c_371_n N_Y_c_550_n 0.00273485f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.33
cc_278 N_A_27_115#_M1009_g N_Y_c_551_n 0.00260839f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=0.9
cc_279 N_A_27_115#_c_320_n N_Y_c_551_n 0.00280419f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=0.9
cc_280 N_A_27_115#_M1013_g N_Y_c_551_n 0.00260839f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=0.9
cc_281 N_A_27_115#_c_387_n N_Y_c_556_n 0.00401146f $X=2.195 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_282 N_A_27_115#_c_320_n N_Y_c_556_n 0.00250559f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.33
cc_283 N_A_27_115#_c_321_n N_Y_c_556_n 0.021445f $X=2.55 $Y=2.625 $X2=2.41
+ $Y2=2.33
cc_284 N_A_27_115#_c_392_n N_Y_c_556_n 0.00401146f $X=2.625 $Y=2.7 $X2=2.41
+ $Y2=2.33
cc_285 N_A_27_115#_c_333_n N_Y_c_556_n 0.00361281f $X=3.055 $Y=2.55 $X2=2.41
+ $Y2=2.33
cc_286 N_A_27_115#_M1014_g N_Y_c_557_n 0.00260839f $X=3.055 $Y=0.895 $X2=3.27
+ $Y2=0.9
cc_287 N_A_27_115#_c_334_n N_Y_c_557_n 0.00280419f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=0.9
cc_288 N_A_27_115#_M1015_g N_Y_c_557_n 0.00260839f $X=3.485 $Y=0.895 $X2=3.27
+ $Y2=0.9
cc_289 N_A_27_115#_c_333_n N_Y_c_562_n 0.00721971f $X=3.055 $Y=2.55 $X2=3.27
+ $Y2=2.33
cc_290 N_A_27_115#_c_398_n N_Y_c_562_n 0.00401146f $X=3.055 $Y=2.7 $X2=3.27
+ $Y2=2.33
cc_291 N_A_27_115#_c_334_n N_Y_c_562_n 0.00250559f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=2.33
cc_292 N_A_27_115#_c_335_n N_Y_c_562_n 0.021445f $X=3.41 $Y=2.625 $X2=3.27
+ $Y2=2.33
cc_293 N_A_27_115#_c_403_n N_Y_c_562_n 0.00401146f $X=3.485 $Y=2.7 $X2=3.27
+ $Y2=2.33
cc_294 N_A_27_115#_M1016_g N_Y_c_563_n 0.00260839f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=0.9
cc_295 N_A_27_115#_c_347_n N_Y_c_563_n 0.00280419f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=0.9
cc_296 N_A_27_115#_M1017_g N_Y_c_563_n 0.00260839f $X=4.345 $Y=0.895 $X2=4.13
+ $Y2=0.9
cc_297 N_A_27_115#_c_409_n N_Y_c_568_n 0.00401146f $X=3.915 $Y=2.7 $X2=4.13
+ $Y2=2.33
cc_298 N_A_27_115#_c_347_n N_Y_c_568_n 0.00250559f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=2.33
cc_299 N_A_27_115#_c_348_n N_Y_c_568_n 0.0206674f $X=4.27 $Y=2.625 $X2=4.13
+ $Y2=2.33
cc_300 N_A_27_115#_c_414_n N_Y_c_568_n 0.00401146f $X=4.345 $Y=2.7 $X2=4.13
+ $Y2=2.33
cc_301 N_A_27_115#_M1003_g N_Y_c_569_n 0.00471447f $X=1.335 $Y=0.895 $X2=1.55
+ $Y2=1.335
cc_302 N_A_27_115#_M1008_g N_Y_c_569_n 0.00259902f $X=1.765 $Y=0.895 $X2=1.55
+ $Y2=1.335
cc_303 N_A_27_115#_c_371_n N_Y_c_569_n 0.00238892f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=1.335
cc_304 N_A_27_115#_c_306_n N_Y_c_572_n 0.00821104f $X=1.37 $Y=2.55 $X2=1.55
+ $Y2=2.215
cc_305 N_A_27_115#_c_307_n N_Y_c_572_n 0.00186325f $X=1.69 $Y=2.625 $X2=1.55
+ $Y2=2.215
cc_306 N_A_27_115#_c_314_n N_Y_c_572_n 0.00194187f $X=1.84 $Y=1.585 $X2=1.55
+ $Y2=2.215
cc_307 N_A_27_115#_c_371_n N_Y_c_572_n 0.00181779f $X=1.43 $Y=1.675 $X2=1.55
+ $Y2=2.215
cc_308 N_A_27_115#_M1003_g Y 0.00251111f $X=1.335 $Y=0.895 $X2=1.555 $Y2=1.96
cc_309 N_A_27_115#_c_306_n Y 0.00892438f $X=1.37 $Y=2.55 $X2=1.555 $Y2=1.96
cc_310 N_A_27_115#_M1008_g Y 0.00251111f $X=1.765 $Y=0.895 $X2=1.555 $Y2=1.96
cc_311 N_A_27_115#_c_314_n Y 0.0131748f $X=1.84 $Y=1.585 $X2=1.555 $Y2=1.96
cc_312 N_A_27_115#_c_371_n Y 0.0148238f $X=1.43 $Y=1.675 $X2=1.555 $Y2=1.96
cc_313 N_A_27_115#_M1008_g N_Y_c_574_n 0.0129109f $X=1.765 $Y=0.895 $X2=2.265
+ $Y2=1.22
cc_314 N_A_27_115#_c_312_n N_Y_c_574_n 0.00213861f $X=2.12 $Y=1.585 $X2=2.265
+ $Y2=1.22
cc_315 N_A_27_115#_M1009_g N_Y_c_574_n 0.0129109f $X=2.195 $Y=0.895 $X2=2.265
+ $Y2=1.22
cc_316 N_A_27_115#_c_314_n N_Y_c_577_n 0.0121767f $X=1.84 $Y=1.585 $X2=2.265
+ $Y2=2.33
cc_317 N_A_27_115#_c_354_n N_Y_c_577_n 0.0158479f $X=1.765 $Y=2.625 $X2=2.265
+ $Y2=2.33
cc_318 N_A_27_115#_M1009_g N_Y_c_578_n 0.00251111f $X=2.195 $Y=0.895 $X2=2.41
+ $Y2=2.215
cc_319 N_A_27_115#_c_320_n N_Y_c_578_n 0.0177725f $X=2.55 $Y=1.585 $X2=2.41
+ $Y2=2.215
cc_320 N_A_27_115#_M1013_g N_Y_c_578_n 0.00251111f $X=2.625 $Y=0.895 $X2=2.41
+ $Y2=2.215
cc_321 N_A_27_115#_c_333_n N_Y_c_578_n 0.00843025f $X=3.055 $Y=2.55 $X2=2.41
+ $Y2=2.215
cc_322 N_A_27_115#_M1013_g N_Y_c_579_n 0.0129109f $X=2.625 $Y=0.895 $X2=3.125
+ $Y2=1.22
cc_323 N_A_27_115#_c_326_n N_Y_c_579_n 0.00213861f $X=2.98 $Y=1.585 $X2=3.125
+ $Y2=1.22
cc_324 N_A_27_115#_M1014_g N_Y_c_579_n 0.0135609f $X=3.055 $Y=0.895 $X2=3.125
+ $Y2=1.22
cc_325 N_A_27_115#_M1009_g N_Y_c_582_n 0.00259902f $X=2.195 $Y=0.895 $X2=2.555
+ $Y2=1.22
cc_326 N_A_27_115#_M1013_g N_Y_c_582_n 0.00259902f $X=2.625 $Y=0.895 $X2=2.555
+ $Y2=1.22
cc_327 N_A_27_115#_c_333_n N_Y_c_585_n 0.0155956f $X=3.055 $Y=2.55 $X2=3.125
+ $Y2=2.33
cc_328 N_A_27_115#_c_357_n N_Y_c_585_n 0.00894336f $X=2.625 $Y=1.585 $X2=3.125
+ $Y2=2.33
cc_329 N_A_27_115#_c_358_n N_Y_c_585_n 0.00903839f $X=2.625 $Y=2.625 $X2=3.125
+ $Y2=2.33
cc_330 N_A_27_115#_c_320_n N_Y_c_586_n 0.00140336f $X=2.55 $Y=1.585 $X2=2.555
+ $Y2=2.33
cc_331 N_A_27_115#_c_333_n N_Y_c_586_n 0.0012308f $X=3.055 $Y=2.55 $X2=2.555
+ $Y2=2.33
cc_332 N_A_27_115#_c_355_n N_Y_c_586_n 0.00140336f $X=2.195 $Y=1.585 $X2=2.555
+ $Y2=2.33
cc_333 N_A_27_115#_c_356_n N_Y_c_586_n 0.00372651f $X=2.195 $Y=2.625 $X2=2.555
+ $Y2=2.33
cc_334 N_A_27_115#_M1014_g N_Y_c_587_n 0.00262362f $X=3.055 $Y=0.895 $X2=3.27
+ $Y2=1.335
cc_335 N_A_27_115#_M1015_g N_Y_c_587_n 0.00371302f $X=3.485 $Y=0.895 $X2=3.27
+ $Y2=1.335
cc_336 N_A_27_115#_M1014_g N_Y_c_590_n 0.00251111f $X=3.055 $Y=0.895 $X2=3.27
+ $Y2=2.215
cc_337 N_A_27_115#_c_333_n N_Y_c_590_n 0.0108556f $X=3.055 $Y=2.55 $X2=3.27
+ $Y2=2.215
cc_338 N_A_27_115#_c_334_n N_Y_c_590_n 0.0177725f $X=3.41 $Y=1.585 $X2=3.27
+ $Y2=2.215
cc_339 N_A_27_115#_M1015_g N_Y_c_590_n 0.00251111f $X=3.485 $Y=0.895 $X2=3.27
+ $Y2=2.215
cc_340 N_A_27_115#_c_361_n N_Y_c_591_n 0.0121767f $X=3.485 $Y=1.585 $X2=3.985
+ $Y2=2.33
cc_341 N_A_27_115#_c_362_n N_Y_c_591_n 0.0158479f $X=3.485 $Y=2.625 $X2=3.985
+ $Y2=2.33
cc_342 N_A_27_115#_c_333_n N_Y_c_592_n 0.00618817f $X=3.055 $Y=2.55 $X2=3.415
+ $Y2=2.33
cc_343 N_A_27_115#_c_334_n N_Y_c_592_n 0.00268861f $X=3.41 $Y=1.585 $X2=3.415
+ $Y2=2.33
cc_344 N_A_27_115#_c_335_n N_Y_c_592_n 0.00357274f $X=3.41 $Y=2.625 $X2=3.415
+ $Y2=2.33
cc_345 N_A_27_115#_M1016_g N_Y_c_593_n 0.00259902f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=1.335
cc_346 N_A_27_115#_M1017_g N_Y_c_593_n 0.00670165f $X=4.345 $Y=0.895 $X2=4.13
+ $Y2=1.335
cc_347 N_A_27_115#_M1016_g N_Y_c_596_n 0.00251111f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=2.215
cc_348 N_A_27_115#_c_347_n N_Y_c_596_n 0.0184054f $X=4.27 $Y=1.585 $X2=4.13
+ $Y2=2.215
cc_349 N_A_27_115#_M1017_g N_Y_c_596_n 0.00251111f $X=4.345 $Y=0.895 $X2=4.13
+ $Y2=2.215
cc_350 N_A_27_115#_c_363_n N_Y_c_596_n 0.00140336f $X=3.915 $Y=1.585 $X2=4.13
+ $Y2=2.215
cc_351 N_A_27_115#_c_364_n N_Y_c_596_n 0.00372651f $X=3.915 $Y=2.625 $X2=4.13
+ $Y2=2.215
cc_352 N_A_27_115#_M1015_g N_Y_c_597_n 8.84842e-19 $X=3.485 $Y=0.895 $X2=4.13
+ $Y2=1.22
cc_353 N_A_27_115#_c_340_n N_Y_c_597_n 0.00213861f $X=3.84 $Y=1.585 $X2=4.13
+ $Y2=1.22
cc_354 N_A_27_115#_M1016_g N_Y_c_597_n 0.0129441f $X=3.915 $Y=0.895 $X2=4.13
+ $Y2=1.22
