* File: sky130_osu_sc_18T_ls__xor2_l.pex.spice
* Created: Thu Oct 29 17:39:01 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%GND 1 2 23 27 29 39 43 49 51
r66 49 51 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r67 43 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r68 37 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.44 $Y=0.305
+ $X2=2.44 $Y2=0.825
r69 30 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r70 25 44 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r71 25 27 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r72 23 37 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.44 $Y2=0.305
r73 23 29 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.152
+ $X2=2.355 $Y2=0.152
r74 23 43 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r75 23 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.17
+ $X2=2.38 $Y2=0.17
r76 23 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r77 23 29 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.355 $Y2=0.152
r78 23 30 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r79 2 39 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.575 $X2=2.44 $Y2=0.825
r80 1 27 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%VDD 1 2 19 23 27 35 41 44 49 50
r45 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=6.49
+ $X2=2.38 $Y2=6.49
r46 44 49 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=2.38 $Y2=6.507
r47 44 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r48 41 53 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r49 41 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r50 35 38 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.44 $Y=4.135
+ $X2=2.44 $Y2=5.835
r51 33 50 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.44 $Y=6.355
+ $X2=2.44 $Y2=6.507
r52 33 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.44 $Y=6.355
+ $X2=2.44 $Y2=5.835
r53 30 32 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r54 28 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r55 28 30 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r56 27 50 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=6.507
+ $X2=2.44 $Y2=6.507
r57 27 32 24.7492 $w=3.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.355 $Y=6.507
+ $X2=1.7 $Y2=6.507
r58 23 26 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r59 21 42 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r60 21 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r61 19 50 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r62 19 53 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r63 19 32 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r64 19 30 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r65 2 38 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.3
+ $Y=3.085 $X2=2.44 $Y2=5.835
r66 2 35 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=2.3
+ $Y=3.085 $X2=2.44 $Y2=4.135
r67 1 26 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r68 1 23 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%A_27_115# 1 2 9 13 17 21 25 29 32 33 35
c76 32 0 6.74854e-20 $X=1.805 $Y=2.765
c77 25 0 1.52002e-20 $X=1.72 $Y=2.225
r78 33 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=2.765
+ $X2=1.805 $Y2=2.93
r79 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=2.765 $X2=1.805 $Y2=2.765
r80 30 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.805 $Y=2.31
+ $X2=1.805 $Y2=2.765
r81 29 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=2.225
+ $X2=0.845 $Y2=2.06
r82 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.225 $X2=0.845 $Y2=2.225
r83 26 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.225
+ $X2=0.26 $Y2=2.225
r84 26 28 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.345 $Y=2.225
+ $X2=0.845 $Y2=2.225
r85 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=2.225
+ $X2=1.805 $Y2=2.31
r86 25 28 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.72 $Y=2.225
+ $X2=0.845 $Y2=2.225
r87 21 23 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r88 19 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.31 $X2=0.26
+ $Y2=2.225
r89 19 21 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=0.26 $Y=2.31
+ $X2=0.26 $Y2=3.455
r90 15 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.14 $X2=0.26
+ $Y2=2.225
r91 15 17 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=0.26 $Y=2.14
+ $X2=0.26 $Y2=0.825
r92 13 41 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.865 $Y=4.585
+ $X2=1.865 $Y2=2.93
r93 9 37 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.06
r94 2 23 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r95 2 21 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r96 1 17 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%A 2 5 6 8 9 13 16 18 19 20 21 22 24 26
+ 27 33 36 37 40 42 45 46 51 52
c122 33 0 3.28297e-19 $X=2.235 $Y=2.22
r123 50 51 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=2.935
+ $X2=0.845 $Y2=3.01
r124 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.145 $Y=3.33
+ $X2=2.145 $Y2=3.33
r125 40 58 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.845 $Y2=3.33
r126 40 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=3.33
+ $X2=1.085 $Y2=3.33
r127 37 42 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.23 $Y=3.33
+ $X2=1.085 $Y2=3.33
r128 36 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2 $Y=3.33
+ $X2=2.145 $Y2=3.33
r129 36 37 0.741419 $w=1.7e-07 $l=7.7e-07 $layer=MET1_cond $X=2 $Y=3.33 $X2=1.23
+ $Y2=3.33
r130 34 52 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=2.22
+ $X2=2.235 $Y2=2.085
r131 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=2.22 $X2=2.235 $Y2=2.22
r132 30 46 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.145 $Y=2.305
+ $X2=2.145 $Y2=3.33
r133 29 33 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.145 $Y=2.22
+ $X2=2.235 $Y2=2.22
r134 29 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.22
+ $X2=2.145 $Y2=2.305
r135 27 50 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=0.845 $Y=2.765
+ $X2=0.845 $Y2=2.935
r136 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.845
+ $Y=2.765 $X2=0.845 $Y2=2.765
r137 24 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=3.245
+ $X2=0.845 $Y2=3.33
r138 23 26 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=2.85
+ $X2=0.845 $Y2=2.765
r139 23 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.845 $Y=2.85
+ $X2=0.845 $Y2=3.245
r140 20 21 41.4471 $w=2e-07 $l=1.25e-07 $layer=POLY_cond $X=0.45 $Y=1.65
+ $X2=0.45 $Y2=1.775
r141 18 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.1 $Y=2.085
+ $X2=2.235 $Y2=2.085
r142 18 19 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.1 $Y=2.085
+ $X2=1.94 $Y2=2.085
r143 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.865 $Y=2.01
+ $X2=1.94 $Y2=2.085
r144 14 16 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.865 $Y=2.01
+ $X2=1.865 $Y2=1.075
r145 13 51 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=3.01
r146 10 22 5.30422 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.55 $Y=2.935
+ $X2=0.45 $Y2=2.935
r147 9 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.71 $Y=2.935
+ $X2=0.845 $Y2=2.935
r148 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=2.935
+ $X2=0.55 $Y2=2.935
r149 6 22 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.45 $Y2=2.935
r150 6 8 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.475 $Y=3.01
+ $X2=0.475 $Y2=4.585
r151 5 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=1.65
r152 2 22 20.4101 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.425 $Y=2.86
+ $X2=0.45 $Y2=2.935
r153 2 21 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=0.425 $Y=2.86
+ $X2=0.425 $Y2=1.775
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%A_238_89# 1 2 9 12 14 17 21 25 29 31
r64 25 27 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.87 $Y=3.455
+ $X2=2.87 $Y2=5.835
r65 23 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.935
+ $X2=2.87 $Y2=1.85
r66 23 25 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=2.87 $Y=1.935
+ $X2=2.87 $Y2=3.455
r67 19 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.765
+ $X2=2.87 $Y2=1.85
r68 19 21 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.87 $Y=1.765
+ $X2=2.87 $Y2=0.825
r69 17 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.85
+ $X2=1.325 $Y2=2.015
r70 17 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.85
+ $X2=1.325 $Y2=1.685
r71 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.85 $X2=1.325 $Y2=1.85
r72 14 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.85
+ $X2=2.87 $Y2=1.85
r73 14 16 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.785 $Y=1.85
+ $X2=1.325 $Y2=1.85
r74 12 32 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=1.265 $Y=4.585
+ $X2=1.265 $Y2=2.015
r75 9 31 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.265 $Y=1.075
+ $X2=1.265 $Y2=1.685
r76 2 27 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.73
+ $Y=3.085 $X2=2.87 $Y2=5.835
r77 2 25 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.73
+ $Y=3.085 $X2=2.87 $Y2=3.455
r78 1 21 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.73
+ $Y=0.575 $X2=2.87 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%B 1 3 4 6 7 8 9 11 13 14 16 17 19 25 27
c56 27 0 6.74854e-20 $X=2.655 $Y=2.805
c57 13 0 1.52002e-20 $X=2.655 $Y=2.6
c58 8 0 1.7901e-19 $X=2.3 $Y=1.725
c59 7 0 1.49287e-19 $X=2.58 $Y=1.725
r60 26 27 20.0833 $w=3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.53 $Y=2.805
+ $X2=2.655 $Y2=2.805
r61 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=2.765 $X2=2.53 $Y2=2.765
r62 21 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.53 $Y=2.96
+ $X2=2.53 $Y2=2.765
r63 19 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.96
+ $X2=2.53 $Y2=2.96
r64 14 27 18.9685 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.655 $Y=3.01
+ $X2=2.655 $Y2=2.805
r65 14 16 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.655 $Y=3.01
+ $X2=2.655 $Y2=4.585
r66 13 27 18.9685 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.655 $Y=2.6
+ $X2=2.655 $Y2=2.805
r67 12 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.8
+ $X2=2.655 $Y2=1.725
r68 12 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.655 $Y=1.8 $X2=2.655
+ $Y2=2.6
r69 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.725
r70 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.075
r71 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.725
+ $X2=2.655 $Y2=1.725
r72 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.58 $Y=1.725 $X2=2.3
+ $Y2=1.725
r73 4 26 49.0033 $w=3e-07 $l=3.94398e-07 $layer=POLY_cond $X=2.225 $Y=3.01
+ $X2=2.53 $Y2=2.805
r74 4 6 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.225 $Y=3.01
+ $X2=2.225 $Y2=4.585
r75 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=1.65
+ $X2=2.3 $Y2=1.725
r76 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.225 $Y=1.65
+ $X2=2.225 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__XOR2_L%Y 1 2 7 9 13 19 23 26 27 29
r58 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.565 $Y=1.48
+ $X2=1.565 $Y2=1.48
r59 29 31 0.0784753 $w=2.23e-07 $l=1.4e-07 $layer=MET1_cond $X=1.425 $Y=1.48
+ $X2=1.565 $Y2=1.48
r60 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.425 $Y=2.59
+ $X2=1.425 $Y2=2.59
r61 21 26 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=2.475
+ $X2=1.425 $Y2=2.59
r62 21 23 0.0433297 $w=1.7e-07 $l=4.5e-08 $layer=MET1_cond $X=1.425 $Y=2.475
+ $X2=1.425 $Y2=2.43
r63 20 29 0.0238602 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.425 $Y=1.595
+ $X2=1.425 $Y2=1.48
r64 20 23 0.804007 $w=1.7e-07 $l=8.35e-07 $layer=MET1_cond $X=1.425 $Y=1.595
+ $X2=1.425 $Y2=2.43
r65 18 27 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.425 $Y=3.205
+ $X2=1.425 $Y2=2.59
r66 18 19 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.537 $Y=3.205
+ $X2=1.537 $Y2=3.375
r67 13 15 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.565 $Y=3.455
+ $X2=1.565 $Y2=5.835
r68 13 19 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=1.565 $Y=3.455
+ $X2=1.565 $Y2=3.375
r69 7 32 9.13816 $w=3.4e-07 $l=2.35e-07 $layer=LI1_cond $X=1.565 $Y=1.245
+ $X2=1.565 $Y2=1.48
r70 7 9 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.565 $Y=1.245
+ $X2=1.565 $Y2=0.825
r71 2 15 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.565 $Y2=5.835
r72 2 13 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.34
+ $Y=3.085 $X2=1.565 $Y2=3.455
r73 1 9 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.34
+ $Y=0.575 $X2=1.565 $Y2=0.825
.ends

