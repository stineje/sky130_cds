* File: sky130_osu_sc_12T_ls__dlat_1.pxi.spice
* Created: Fri Nov 12 15:36:56 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%GND N_GND_M1002_s N_GND_M1003_d N_GND_M1006_s
+ N_GND_M1007_d N_GND_M1002_b N_GND_c_2_p N_GND_c_3_p N_GND_c_26_p N_GND_c_41_p
+ N_GND_c_7_p N_GND_c_8_p N_GND_c_78_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_LS__DLAT_1%GND
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%VDD N_VDD_M1013_s N_VDD_M1015_d N_VDD_M1000_s
+ N_VDD_M1004_d N_VDD_M1013_b N_VDD_c_123_p N_VDD_c_124_p N_VDD_c_139_p
+ N_VDD_c_140_p N_VDD_c_127_p N_VDD_c_128_p N_VDD_c_161_p N_VDD_c_174_p VDD
+ N_VDD_c_125_p PM_SKY130_OSU_SC_12T_LS__DLAT_1%VDD
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%D N_D_M1012_d N_D_M1011_d N_D_M1002_g
+ N_D_M1013_g N_D_c_189_n N_D_M1006_g N_D_M1000_g N_D_c_194_n N_D_c_196_n
+ N_D_c_198_n N_D_c_199_n N_D_c_237_p N_D_c_310_p N_D_c_224_n N_D_c_200_n
+ N_D_c_201_n N_D_c_203_n N_D_c_205_n N_D_c_207_n N_D_c_208_n D N_D_c_211_n
+ N_D_c_212_n N_D_c_213_n PM_SKY130_OSU_SC_12T_LS__DLAT_1%D
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%CK N_CK_M1012_g N_CK_M1014_g N_CK_M1005_g
+ N_CK_c_311_n N_CK_M1008_g N_CK_c_312_n N_CK_c_313_n N_CK_c_314_n N_CK_c_317_n
+ N_CK_c_318_n N_CK_c_323_n N_CK_c_324_n N_CK_c_325_n N_CK_c_326_n N_CK_c_327_n
+ N_CK_c_328_n N_CK_c_329_n N_CK_c_330_n CK PM_SKY130_OSU_SC_12T_LS__DLAT_1%CK
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%A_157_349# N_A_157_349#_M1005_d
+ N_A_157_349#_M1008_d N_A_157_349#_M1011_g N_A_157_349#_c_458_n
+ N_A_157_349#_c_459_n N_A_157_349#_M1010_g N_A_157_349#_c_463_n
+ N_A_157_349#_c_464_n N_A_157_349#_c_465_n N_A_157_349#_c_477_n
+ N_A_157_349#_c_469_n N_A_157_349#_c_470_n N_A_157_349#_c_482_n
+ N_A_157_349#_c_471_n N_A_157_349#_c_472_n N_A_157_349#_c_473_n
+ PM_SKY130_OSU_SC_12T_LS__DLAT_1%A_157_349#
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%A_349_89# N_A_349_89#_M1006_d
+ N_A_349_89#_M1000_d N_A_349_89#_M1003_g N_A_349_89#_M1015_g
+ N_A_349_89#_c_598_n N_A_349_89#_M1007_g N_A_349_89#_M1004_g
+ N_A_349_89#_c_603_n N_A_349_89#_c_605_n N_A_349_89#_c_606_n
+ N_A_349_89#_c_607_n N_A_349_89#_c_608_n N_A_349_89#_c_609_n
+ N_A_349_89#_c_612_n N_A_349_89#_c_613_n N_A_349_89#_c_614_n
+ N_A_349_89#_c_615_n N_A_349_89#_c_616_n N_A_349_89#_c_617_n
+ N_A_349_89#_c_618_n N_A_349_89#_c_619_n N_A_349_89#_c_620_n
+ PM_SKY130_OSU_SC_12T_LS__DLAT_1%A_349_89#
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%ON N_ON_M1007_s N_ON_M1004_s N_ON_M1009_g
+ N_ON_M1001_g N_ON_c_763_n N_ON_c_764_n N_ON_c_767_n N_ON_c_768_n N_ON_c_769_n
+ N_ON_c_771_n N_ON_c_772_n N_ON_c_773_n N_ON_c_774_n N_ON_c_775_n ON
+ PM_SKY130_OSU_SC_12T_LS__DLAT_1%ON
x_PM_SKY130_OSU_SC_12T_LS__DLAT_1%Q N_Q_M1009_d N_Q_M1001_d N_Q_c_837_n
+ N_Q_c_843_n N_Q_c_839_n N_Q_c_840_n N_Q_c_841_n Q
+ PM_SKY130_OSU_SC_12T_LS__DLAT_1%Q
cc_1 N_GND_M1002_b N_D_M1002_g 0.0476101f $X=-0.045 $Y=0 $X2=0.5 $Y2=0.835
cc_2 N_GND_c_2_p N_D_M1002_g 0.00502587f $X=0.285 $Y=0.74 $X2=0.5 $Y2=0.835
cc_3 N_GND_c_3_p N_D_M1002_g 0.00606474f $X=1.95 $Y=0.152 $X2=0.5 $Y2=0.835
cc_4 N_GND_c_4_p N_D_M1002_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.5 $Y2=0.835
cc_5 N_GND_M1002_b N_D_M1013_g 0.0379931f $X=-0.045 $Y=0 $X2=0.5 $Y2=3.235
cc_6 N_GND_M1002_b N_D_c_189_n 0.0221119f $X=-0.045 $Y=0 $X2=3.2 $Y2=1.205
cc_7 N_GND_c_7_p N_D_c_189_n 0.00502587f $X=2.985 $Y=0.74 $X2=3.2 $Y2=1.205
cc_8 N_GND_c_8_p N_D_c_189_n 0.00606474f $X=4.28 $Y=0.152 $X2=3.2 $Y2=1.205
cc_9 N_GND_c_4_p N_D_c_189_n 0.00468827f $X=4.42 $Y=0.19 $X2=3.2 $Y2=1.205
cc_10 N_GND_M1002_b N_D_M1000_g 0.0594603f $X=-0.045 $Y=0 $X2=3.2 $Y2=3.235
cc_11 N_GND_M1002_b N_D_c_194_n 0.0361824f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.74
cc_12 N_GND_c_2_p N_D_c_194_n 0.00142801f $X=0.285 $Y=0.74 $X2=0.44 $Y2=1.74
cc_13 N_GND_M1002_b N_D_c_196_n 0.0483832f $X=-0.045 $Y=0 $X2=3.2 $Y2=1.37
cc_14 N_GND_c_7_p N_D_c_196_n 0.00378206f $X=2.985 $Y=0.74 $X2=3.2 $Y2=1.37
cc_15 N_GND_M1002_b N_D_c_198_n 0.00248795f $X=-0.045 $Y=0 $X2=0.58 $Y2=1.37
cc_16 N_GND_M1002_b N_D_c_199_n 0.00380459f $X=-0.045 $Y=0 $X2=0.58 $Y2=2.62
cc_17 N_GND_M1002_b N_D_c_200_n 0.00919218f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.34
cc_18 N_GND_M1002_b N_D_c_201_n 0.00162209f $X=-0.045 $Y=0 $X2=2.995 $Y2=1.37
cc_19 N_GND_c_7_p N_D_c_201_n 0.00461497f $X=2.985 $Y=0.74 $X2=2.995 $Y2=1.37
cc_20 N_GND_M1002_b N_D_c_203_n 0.00652056f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.74
cc_21 N_GND_c_2_p N_D_c_203_n 3.46856e-19 $X=0.285 $Y=0.74 $X2=0.44 $Y2=1.74
cc_22 N_GND_c_3_p N_D_c_205_n 0.0145094f $X=1.95 $Y=0.152 $X2=1.26 $Y2=0.74
cc_23 N_GND_c_4_p N_D_c_205_n 0.00983195f $X=4.42 $Y=0.19 $X2=1.26 $Y2=0.74
cc_24 N_GND_M1002_b N_D_c_207_n 0.00716398f $X=-0.045 $Y=0 $X2=0.725 $Y2=1.37
cc_25 N_GND_M1002_b N_D_c_208_n 0.0300537f $X=-0.045 $Y=0 $X2=2.85 $Y2=1.37
cc_26 N_GND_c_26_p N_D_c_208_n 0.00707192f $X=2.035 $Y=0.74 $X2=2.85 $Y2=1.37
cc_27 N_GND_M1002_b D 0.011851f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.74
cc_28 N_GND_M1002_b N_D_c_211_n 0.00546614f $X=-0.045 $Y=0 $X2=1.115 $Y2=1.34
cc_29 N_GND_M1002_b N_D_c_212_n 0.00431866f $X=-0.045 $Y=0 $X2=1.405 $Y2=1.34
cc_30 N_GND_M1002_b N_D_c_213_n 9.68419e-19 $X=-0.045 $Y=0 $X2=2.995 $Y2=1.37
cc_31 N_GND_c_7_p N_D_c_213_n 0.00379624f $X=2.985 $Y=0.74 $X2=2.995 $Y2=1.37
cc_32 N_GND_M1002_b N_CK_c_311_n 0.0307453f $X=-0.045 $Y=0 $X2=2.25 $Y2=2.45
cc_33 N_GND_M1002_b N_CK_c_312_n 0.0445582f $X=-0.045 $Y=0 $X2=2.305 $Y2=2.12
cc_34 N_GND_M1002_b N_CK_c_313_n 0.0267362f $X=-0.045 $Y=0 $X2=0.92 $Y2=1.37
cc_35 N_GND_M1002_b N_CK_c_314_n 0.0174883f $X=-0.045 $Y=0 $X2=0.92 $Y2=1.205
cc_36 N_GND_c_3_p N_CK_c_314_n 0.00606474f $X=1.95 $Y=0.152 $X2=0.92 $Y2=1.205
cc_37 N_GND_c_4_p N_CK_c_314_n 0.00468827f $X=4.42 $Y=0.19 $X2=0.92 $Y2=1.205
cc_38 N_GND_M1002_b N_CK_c_317_n 0.0219022f $X=-0.045 $Y=0 $X2=1.4 $Y2=2.285
cc_39 N_GND_M1002_b N_CK_c_318_n 0.0183851f $X=-0.045 $Y=0 $X2=2.277 $Y2=1.205
cc_40 N_GND_c_26_p N_CK_c_318_n 0.00308284f $X=2.035 $Y=0.74 $X2=2.277 $Y2=1.205
cc_41 N_GND_c_41_p N_CK_c_318_n 0.00606474f $X=2.9 $Y=0.152 $X2=2.277 $Y2=1.205
cc_42 N_GND_c_7_p N_CK_c_318_n 0.00359543f $X=2.985 $Y=0.74 $X2=2.277 $Y2=1.205
cc_43 N_GND_c_4_p N_CK_c_318_n 0.00468827f $X=4.42 $Y=0.19 $X2=2.277 $Y2=1.205
cc_44 N_GND_M1002_b N_CK_c_323_n 0.0141068f $X=-0.045 $Y=0 $X2=2.277 $Y2=1.355
cc_45 N_GND_M1002_b N_CK_c_324_n 0.00861118f $X=-0.045 $Y=0 $X2=0.92 $Y2=1.37
cc_46 N_GND_M1002_b N_CK_c_325_n 0.00500343f $X=-0.045 $Y=0 $X2=1.315 $Y2=2.11
cc_47 N_GND_M1002_b N_CK_c_326_n 9.63154e-19 $X=-0.045 $Y=0 $X2=1.005 $Y2=2.11
cc_48 N_GND_M1002_b N_CK_c_327_n 7.11312e-19 $X=-0.045 $Y=0 $X2=2.395 $Y2=2.11
cc_49 N_GND_M1002_b N_CK_c_328_n 0.00120157f $X=-0.045 $Y=0 $X2=1.4 $Y2=2.11
cc_50 N_GND_M1002_b N_CK_c_329_n 0.0139101f $X=-0.045 $Y=0 $X2=2.25 $Y2=2.11
cc_51 N_GND_M1002_b N_CK_c_330_n 0.00256396f $X=-0.045 $Y=0 $X2=1.545 $Y2=2.11
cc_52 N_GND_M1002_b CK 0.00144547f $X=-0.045 $Y=0 $X2=2.395 $Y2=2.11
cc_53 N_GND_M1002_b N_A_157_349#_M1011_g 0.0286835f $X=-0.045 $Y=0 $X2=0.86
+ $Y2=3.235
cc_54 N_GND_M1002_b N_A_157_349#_c_458_n 0.0211051f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=1.825
cc_55 N_GND_M1002_b N_A_157_349#_c_459_n 0.00713103f $X=-0.045 $Y=0 $X2=0.935
+ $Y2=1.825
cc_56 N_GND_M1002_b N_A_157_349#_M1010_g 0.0351889f $X=-0.045 $Y=0 $X2=1.46
+ $Y2=0.835
cc_57 N_GND_c_3_p N_A_157_349#_M1010_g 0.00606474f $X=1.95 $Y=0.152 $X2=1.46
+ $Y2=0.835
cc_58 N_GND_c_4_p N_A_157_349#_M1010_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.46
+ $Y2=0.835
cc_59 N_GND_M1002_b N_A_157_349#_c_463_n 0.0257525f $X=-0.045 $Y=0 $X2=1.4
+ $Y2=1.74
cc_60 N_GND_M1002_b N_A_157_349#_c_464_n 0.00205129f $X=-0.045 $Y=0 $X2=1.4
+ $Y2=1.74
cc_61 N_GND_M1002_b N_A_157_349#_c_465_n 0.0151485f $X=-0.045 $Y=0 $X2=2.465
+ $Y2=0.74
cc_62 N_GND_c_41_p N_A_157_349#_c_465_n 0.00736239f $X=2.9 $Y=0.152 $X2=2.465
+ $Y2=0.74
cc_63 N_GND_c_7_p N_A_157_349#_c_465_n 0.0140971f $X=2.985 $Y=0.74 $X2=2.465
+ $Y2=0.74
cc_64 N_GND_c_4_p N_A_157_349#_c_465_n 0.00476261f $X=4.42 $Y=0.19 $X2=2.465
+ $Y2=0.74
cc_65 N_GND_M1002_b N_A_157_349#_c_469_n 0.0123446f $X=-0.045 $Y=0 $X2=2.735
+ $Y2=2.62
cc_66 N_GND_M1002_b N_A_157_349#_c_470_n 0.011016f $X=-0.045 $Y=0 $X2=2.735
+ $Y2=1.725
cc_67 N_GND_M1002_b N_A_157_349#_c_471_n 0.00149882f $X=-0.045 $Y=0 $X2=1.545
+ $Y2=1.725
cc_68 N_GND_M1002_b N_A_157_349#_c_472_n 0.00217465f $X=-0.045 $Y=0 $X2=2.465
+ $Y2=1.74
cc_69 N_GND_M1002_b N_A_157_349#_c_473_n 0.00682657f $X=-0.045 $Y=0 $X2=2.32
+ $Y2=1.74
cc_70 N_GND_M1002_b N_A_349_89#_M1003_g 0.0337299f $X=-0.045 $Y=0 $X2=1.82
+ $Y2=0.835
cc_71 N_GND_c_3_p N_A_349_89#_M1003_g 0.00606474f $X=1.95 $Y=0.152 $X2=1.82
+ $Y2=0.835
cc_72 N_GND_c_26_p N_A_349_89#_M1003_g 0.00308284f $X=2.035 $Y=0.74 $X2=1.82
+ $Y2=0.835
cc_73 N_GND_c_4_p N_A_349_89#_M1003_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.82
+ $Y2=0.835
cc_74 N_GND_M1002_b N_A_349_89#_M1015_g 0.0286123f $X=-0.045 $Y=0 $X2=1.82
+ $Y2=3.235
cc_75 N_GND_M1002_b N_A_349_89#_c_598_n 0.0524785f $X=-0.045 $Y=0 $X2=4.1
+ $Y2=1.905
cc_76 N_GND_M1002_b N_A_349_89#_M1007_g 0.024302f $X=-0.045 $Y=0 $X2=4.15
+ $Y2=0.835
cc_77 N_GND_c_8_p N_A_349_89#_M1007_g 0.00606474f $X=4.28 $Y=0.152 $X2=4.15
+ $Y2=0.835
cc_78 N_GND_c_78_p N_A_349_89#_M1007_g 0.00308284f $X=4.365 $Y=0.74 $X2=4.15
+ $Y2=0.835
cc_79 N_GND_c_4_p N_A_349_89#_M1007_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.15
+ $Y2=0.835
cc_80 N_GND_M1002_b N_A_349_89#_c_603_n 0.0263018f $X=-0.045 $Y=0 $X2=1.88
+ $Y2=1.74
cc_81 N_GND_c_26_p N_A_349_89#_c_603_n 0.0014075f $X=2.035 $Y=0.74 $X2=1.88
+ $Y2=1.74
cc_82 N_GND_M1002_b N_A_349_89#_c_605_n 0.0266574f $X=-0.045 $Y=0 $X2=4.125
+ $Y2=2.36
cc_83 N_GND_M1002_b N_A_349_89#_c_606_n 0.00535389f $X=-0.045 $Y=0 $X2=4.125
+ $Y2=2.49
cc_84 N_GND_M1002_b N_A_349_89#_c_607_n 8.70944e-19 $X=-0.045 $Y=0 $X2=1.882
+ $Y2=1.812
cc_85 N_GND_M1002_b N_A_349_89#_c_608_n 0.00374026f $X=-0.045 $Y=0 $X2=1.88
+ $Y2=2.48
cc_86 N_GND_M1002_b N_A_349_89#_c_609_n 0.0143842f $X=-0.045 $Y=0 $X2=3.415
+ $Y2=0.74
cc_87 N_GND_c_8_p N_A_349_89#_c_609_n 0.00757793f $X=4.28 $Y=0.152 $X2=3.415
+ $Y2=0.74
cc_88 N_GND_c_4_p N_A_349_89#_c_609_n 0.00476261f $X=4.42 $Y=0.19 $X2=3.415
+ $Y2=0.74
cc_89 N_GND_M1002_b N_A_349_89#_c_612_n 0.013534f $X=-0.045 $Y=0 $X2=3.415
+ $Y2=2.935
cc_90 N_GND_M1002_b N_A_349_89#_c_613_n 0.0121972f $X=-0.045 $Y=0 $X2=4.035
+ $Y2=1.74
cc_91 N_GND_M1002_b N_A_349_89#_c_614_n 0.00242672f $X=-0.045 $Y=0 $X2=3.415
+ $Y2=1.74
cc_92 N_GND_M1002_b N_A_349_89#_c_615_n 0.00262889f $X=-0.045 $Y=0 $X2=2.755
+ $Y2=2.48
cc_93 N_GND_M1002_b N_A_349_89#_c_616_n 0.00120404f $X=-0.045 $Y=0 $X2=2.025
+ $Y2=2.48
cc_94 N_GND_M1002_b N_A_349_89#_c_617_n 0.0053881f $X=-0.045 $Y=0 $X2=2.827
+ $Y2=2.395
cc_95 N_GND_M1002_b N_A_349_89#_c_618_n 0.0342266f $X=-0.045 $Y=0 $X2=3.9
+ $Y2=1.74
cc_96 N_GND_M1002_b N_A_349_89#_c_619_n 3.47949e-19 $X=-0.045 $Y=0 $X2=2.9
+ $Y2=1.74
cc_97 N_GND_M1002_b N_A_349_89#_c_620_n 0.00114019f $X=-0.045 $Y=0 $X2=4.035
+ $Y2=1.74
cc_98 N_GND_M1002_b N_ON_M1009_g 0.061038f $X=-0.045 $Y=0 $X2=4.58 $Y2=0.835
cc_99 N_GND_c_78_p N_ON_M1009_g 0.00308284f $X=4.365 $Y=0.74 $X2=4.58 $Y2=0.835
cc_100 N_GND_c_4_p N_ON_M1009_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.58 $Y2=0.835
cc_101 N_GND_M1002_b N_ON_M1001_g 0.0148247f $X=-0.045 $Y=0 $X2=4.58 $Y2=3.235
cc_102 N_GND_M1002_b N_ON_c_763_n 0.0284977f $X=-0.045 $Y=0 $X2=4.52 $Y2=2.015
cc_103 N_GND_M1002_b N_ON_c_764_n 0.00589726f $X=-0.045 $Y=0 $X2=3.935 $Y2=0.74
cc_104 N_GND_c_8_p N_ON_c_764_n 0.00745733f $X=4.28 $Y=0.152 $X2=3.935 $Y2=0.74
cc_105 N_GND_c_4_p N_ON_c_764_n 0.00476261f $X=4.42 $Y=0.19 $X2=3.935 $Y2=0.74
cc_106 N_GND_M1002_b N_ON_c_767_n 0.00173247f $X=-0.045 $Y=0 $X2=3.935 $Y2=2.195
cc_107 N_GND_M1002_b N_ON_c_768_n 0.00445082f $X=-0.045 $Y=0 $X2=3.935 $Y2=3.615
cc_108 N_GND_M1002_b N_ON_c_769_n 0.00947205f $X=-0.045 $Y=0 $X2=4.43 $Y2=1.4
cc_109 N_GND_c_78_p N_ON_c_769_n 0.00740779f $X=4.365 $Y=0.74 $X2=4.43 $Y2=1.4
cc_110 N_GND_M1002_b N_ON_c_771_n 0.0026304f $X=-0.045 $Y=0 $X2=4.02 $Y2=1.4
cc_111 N_GND_M1002_b N_ON_c_772_n 0.0130744f $X=-0.045 $Y=0 $X2=4.435 $Y2=2.11
cc_112 N_GND_M1002_b N_ON_c_773_n 0.00154106f $X=-0.045 $Y=0 $X2=4.517 $Y2=1.658
cc_113 N_GND_M1002_b N_ON_c_774_n 5.47532e-19 $X=-0.045 $Y=0 $X2=4.52 $Y2=2.015
cc_114 N_GND_M1002_b N_ON_c_775_n 5.00369e-19 $X=-0.045 $Y=0 $X2=4.517 $Y2=1.745
cc_115 N_GND_M1002_b ON 0.00962953f $X=-0.045 $Y=0 $X2=3.935 $Y2=2.11
cc_116 N_GND_M1002_b N_Q_c_837_n 0.00910394f $X=-0.045 $Y=0 $X2=4.795 $Y2=0.74
cc_117 N_GND_c_4_p N_Q_c_837_n 0.00475329f $X=4.42 $Y=0.19 $X2=4.795 $Y2=0.74
cc_118 N_GND_M1002_b N_Q_c_839_n 0.0107289f $X=-0.045 $Y=0 $X2=4.827 $Y2=1.155
cc_119 N_GND_M1002_b N_Q_c_840_n 0.00185739f $X=-0.045 $Y=0 $X2=4.795 $Y2=2.48
cc_120 N_GND_M1002_b N_Q_c_841_n 0.0577223f $X=-0.045 $Y=0 $X2=4.827 $Y2=2.395
cc_121 N_GND_M1002_b Q 0.00682487f $X=-0.045 $Y=0 $X2=4.795 $Y2=2.48
cc_122 N_VDD_M1013_b N_D_M1013_g 0.0239842f $X=-0.045 $Y=2.425 $X2=0.5 $Y2=3.235
cc_123 N_VDD_c_123_p N_D_M1013_g 0.00713292f $X=0.285 $Y=3.275 $X2=0.5 $Y2=3.235
cc_124 N_VDD_c_124_p N_D_M1013_g 0.00606474f $X=1.95 $Y=4.287 $X2=0.5 $Y2=3.235
cc_125 N_VDD_c_125_p N_D_M1013_g 0.00468827f $X=4.42 $Y=4.25 $X2=0.5 $Y2=3.235
cc_126 N_VDD_M1013_b N_D_M1000_g 0.0260072f $X=-0.045 $Y=2.425 $X2=3.2 $Y2=3.235
cc_127 N_VDD_c_127_p N_D_M1000_g 0.00713292f $X=2.985 $Y=3.275 $X2=3.2 $Y2=3.235
cc_128 N_VDD_c_128_p N_D_M1000_g 0.00606474f $X=4.28 $Y=4.287 $X2=3.2 $Y2=3.235
cc_129 N_VDD_c_125_p N_D_M1000_g 0.00468827f $X=4.42 $Y=4.25 $X2=3.2 $Y2=3.235
cc_130 N_VDD_M1013_b N_D_c_199_n 0.00168314f $X=-0.045 $Y=2.425 $X2=0.58
+ $Y2=2.62
cc_131 N_VDD_M1013_b N_D_c_224_n 0.00313975f $X=-0.045 $Y=2.425 $X2=1.16
+ $Y2=3.275
cc_132 N_VDD_c_124_p N_D_c_224_n 0.0149461f $X=1.95 $Y=4.287 $X2=1.16 $Y2=3.275
cc_133 N_VDD_c_125_p N_D_c_224_n 0.00958198f $X=4.42 $Y=4.25 $X2=1.16 $Y2=3.275
cc_134 N_VDD_M1013_b N_CK_M1014_g 0.0201163f $X=-0.045 $Y=2.425 $X2=1.46
+ $Y2=3.235
cc_135 N_VDD_c_124_p N_CK_M1014_g 0.00606474f $X=1.95 $Y=4.287 $X2=1.46
+ $Y2=3.235
cc_136 N_VDD_c_125_p N_CK_M1014_g 0.00468827f $X=4.42 $Y=4.25 $X2=1.46 $Y2=3.235
cc_137 N_VDD_M1013_b N_CK_c_311_n 0.007968f $X=-0.045 $Y=2.425 $X2=2.25 $Y2=2.45
cc_138 N_VDD_M1013_b N_CK_M1008_g 0.0218804f $X=-0.045 $Y=2.425 $X2=2.25
+ $Y2=3.235
cc_139 N_VDD_c_139_p N_CK_M1008_g 0.00354579f $X=2.035 $Y=3.275 $X2=2.25
+ $Y2=3.235
cc_140 N_VDD_c_140_p N_CK_M1008_g 0.00606474f $X=2.9 $Y=4.287 $X2=2.25 $Y2=3.235
cc_141 N_VDD_c_127_p N_CK_M1008_g 0.00463923f $X=2.985 $Y=3.275 $X2=2.25
+ $Y2=3.235
cc_142 N_VDD_c_125_p N_CK_M1008_g 0.00468827f $X=4.42 $Y=4.25 $X2=2.25 $Y2=3.235
cc_143 N_VDD_M1013_b N_CK_c_317_n 0.00486793f $X=-0.045 $Y=2.425 $X2=1.4
+ $Y2=2.285
cc_144 N_VDD_M1013_b N_CK_c_327_n 0.0010436f $X=-0.045 $Y=2.425 $X2=2.395
+ $Y2=2.11
cc_145 N_VDD_M1013_b N_CK_c_328_n 0.0022456f $X=-0.045 $Y=2.425 $X2=1.4 $Y2=2.11
cc_146 N_VDD_M1013_b N_A_157_349#_M1011_g 0.0214821f $X=-0.045 $Y=2.425 $X2=0.86
+ $Y2=3.235
cc_147 N_VDD_c_124_p N_A_157_349#_M1011_g 0.00606474f $X=1.95 $Y=4.287 $X2=0.86
+ $Y2=3.235
cc_148 N_VDD_c_125_p N_A_157_349#_M1011_g 0.00468827f $X=4.42 $Y=4.25 $X2=0.86
+ $Y2=3.235
cc_149 N_VDD_M1013_b N_A_157_349#_c_477_n 0.00156053f $X=-0.045 $Y=2.425
+ $X2=2.465 $Y2=2.935
cc_150 N_VDD_c_140_p N_A_157_349#_c_477_n 0.00736239f $X=2.9 $Y=4.287 $X2=2.465
+ $Y2=2.935
cc_151 N_VDD_c_127_p N_A_157_349#_c_477_n 0.0358835f $X=2.985 $Y=3.275 $X2=2.465
+ $Y2=2.935
cc_152 N_VDD_c_125_p N_A_157_349#_c_477_n 0.00476261f $X=4.42 $Y=4.25 $X2=2.465
+ $Y2=2.935
cc_153 N_VDD_M1013_b N_A_157_349#_c_469_n 0.00543969f $X=-0.045 $Y=2.425
+ $X2=2.735 $Y2=2.62
cc_154 N_VDD_M1013_b N_A_157_349#_c_482_n 0.0119291f $X=-0.045 $Y=2.425
+ $X2=2.735 $Y2=2.705
cc_155 N_VDD_M1013_b N_A_349_89#_M1015_g 0.0178558f $X=-0.045 $Y=2.425 $X2=1.82
+ $Y2=3.235
cc_156 N_VDD_c_124_p N_A_349_89#_M1015_g 0.00606474f $X=1.95 $Y=4.287 $X2=1.82
+ $Y2=3.235
cc_157 N_VDD_c_139_p N_A_349_89#_M1015_g 0.00354579f $X=2.035 $Y=3.275 $X2=1.82
+ $Y2=3.235
cc_158 N_VDD_c_125_p N_A_349_89#_M1015_g 0.00468827f $X=4.42 $Y=4.25 $X2=1.82
+ $Y2=3.235
cc_159 N_VDD_M1013_b N_A_349_89#_c_606_n 0.027733f $X=-0.045 $Y=2.425 $X2=4.125
+ $Y2=2.49
cc_160 N_VDD_c_128_p N_A_349_89#_c_606_n 0.00606474f $X=4.28 $Y=4.287 $X2=4.125
+ $Y2=2.49
cc_161 N_VDD_c_161_p N_A_349_89#_c_606_n 0.00354579f $X=4.365 $Y=3.615 $X2=4.125
+ $Y2=2.49
cc_162 N_VDD_c_125_p N_A_349_89#_c_606_n 0.00468827f $X=4.42 $Y=4.25 $X2=4.125
+ $Y2=2.49
cc_163 N_VDD_M1013_b N_A_349_89#_c_608_n 0.00248522f $X=-0.045 $Y=2.425 $X2=1.88
+ $Y2=2.48
cc_164 N_VDD_c_139_p N_A_349_89#_c_608_n 4.51972e-19 $X=2.035 $Y=3.275 $X2=1.88
+ $Y2=2.48
cc_165 N_VDD_M1013_b N_A_349_89#_c_612_n 0.00576734f $X=-0.045 $Y=2.425
+ $X2=3.415 $Y2=2.935
cc_166 N_VDD_c_128_p N_A_349_89#_c_612_n 0.00757793f $X=4.28 $Y=4.287 $X2=3.415
+ $Y2=2.935
cc_167 N_VDD_c_125_p N_A_349_89#_c_612_n 0.00476261f $X=4.42 $Y=4.25 $X2=3.415
+ $Y2=2.935
cc_168 N_VDD_M1013_b N_A_349_89#_c_615_n 0.0114825f $X=-0.045 $Y=2.425 $X2=2.755
+ $Y2=2.48
cc_169 N_VDD_c_139_p N_A_349_89#_c_615_n 0.003766f $X=2.035 $Y=3.275 $X2=2.755
+ $Y2=2.48
cc_170 N_VDD_M1013_b N_A_349_89#_c_616_n 0.00615199f $X=-0.045 $Y=2.425
+ $X2=2.025 $Y2=2.48
cc_171 N_VDD_c_139_p N_A_349_89#_c_616_n 0.00283724f $X=2.035 $Y=3.275 $X2=2.025
+ $Y2=2.48
cc_172 N_VDD_M1013_b N_ON_M1001_g 0.0267653f $X=-0.045 $Y=2.425 $X2=4.58
+ $Y2=3.235
cc_173 N_VDD_c_161_p N_ON_M1001_g 0.00354579f $X=4.365 $Y=3.615 $X2=4.58
+ $Y2=3.235
cc_174 N_VDD_c_174_p N_ON_M1001_g 0.00606474f $X=4.42 $Y=4.25 $X2=4.58 $Y2=3.235
cc_175 N_VDD_c_125_p N_ON_M1001_g 0.00468827f $X=4.42 $Y=4.25 $X2=4.58 $Y2=3.235
cc_176 N_VDD_M1013_b N_ON_c_768_n 0.00535954f $X=-0.045 $Y=2.425 $X2=3.935
+ $Y2=3.615
cc_177 N_VDD_c_128_p N_ON_c_768_n 0.00745733f $X=4.28 $Y=4.287 $X2=3.935
+ $Y2=3.615
cc_178 N_VDD_c_125_p N_ON_c_768_n 0.00476261f $X=4.42 $Y=4.25 $X2=3.935
+ $Y2=3.615
cc_179 N_VDD_M1013_b N_Q_c_843_n 0.00297074f $X=-0.045 $Y=2.425 $X2=4.795
+ $Y2=3.615
cc_180 N_VDD_c_174_p N_Q_c_843_n 0.00757793f $X=4.42 $Y=4.25 $X2=4.795 $Y2=3.615
cc_181 N_VDD_c_125_p N_Q_c_843_n 0.00476261f $X=4.42 $Y=4.25 $X2=4.795 $Y2=3.615
cc_182 N_VDD_M1013_b N_Q_c_840_n 0.00562959f $X=-0.045 $Y=2.425 $X2=4.795
+ $Y2=2.48
cc_183 N_VDD_M1013_b Q 0.0111813f $X=-0.045 $Y=2.425 $X2=4.795 $Y2=2.48
cc_184 N_D_M1000_g N_CK_c_311_n 0.00468822f $X=3.2 $Y=3.235 $X2=2.25 $Y2=2.45
cc_185 N_D_c_208_n N_CK_c_312_n 0.00321559f $X=2.85 $Y=1.37 $X2=2.305 $Y2=2.12
cc_186 N_D_c_198_n N_CK_c_313_n 0.00120463f $X=0.58 $Y=1.37 $X2=0.92 $Y2=1.37
cc_187 N_D_c_200_n N_CK_c_313_n 0.0015339f $X=1.26 $Y=1.34 $X2=0.92 $Y2=1.37
cc_188 N_D_c_205_n N_CK_c_313_n 0.0018818f $X=1.26 $Y=0.74 $X2=0.92 $Y2=1.37
cc_189 N_D_c_207_n N_CK_c_313_n 6.81488e-19 $X=0.725 $Y=1.37 $X2=0.92 $Y2=1.37
cc_190 N_D_c_211_n N_CK_c_313_n 0.00617909f $X=1.115 $Y=1.34 $X2=0.92 $Y2=1.37
cc_191 N_D_c_212_n N_CK_c_313_n 7.50094e-19 $X=1.405 $Y=1.34 $X2=0.92 $Y2=1.37
cc_192 N_D_M1002_g N_CK_c_314_n 0.0679283f $X=0.5 $Y=0.835 $X2=0.92 $Y2=1.205
cc_193 N_D_c_200_n N_CK_c_314_n 0.00614655f $X=1.26 $Y=1.34 $X2=0.92 $Y2=1.205
cc_194 N_D_c_237_p N_CK_c_317_n 0.00150627f $X=0.99 $Y=2.705 $X2=1.4 $Y2=2.285
cc_195 N_D_c_196_n N_CK_c_323_n 0.00712865f $X=3.2 $Y=1.37 $X2=2.277 $Y2=1.355
cc_196 N_D_c_208_n N_CK_c_323_n 0.0102303f $X=2.85 $Y=1.37 $X2=2.277 $Y2=1.355
cc_197 N_D_M1002_g N_CK_c_324_n 0.00157055f $X=0.5 $Y=0.835 $X2=0.92 $Y2=1.37
cc_198 N_D_c_194_n N_CK_c_324_n 2.72267e-19 $X=0.44 $Y=1.74 $X2=0.92 $Y2=1.37
cc_199 N_D_c_198_n N_CK_c_324_n 0.0511906f $X=0.58 $Y=1.37 $X2=0.92 $Y2=1.37
cc_200 N_D_c_200_n N_CK_c_324_n 0.0166667f $X=1.26 $Y=1.34 $X2=0.92 $Y2=1.37
cc_201 N_D_c_205_n N_CK_c_324_n 6.02726e-19 $X=1.26 $Y=0.74 $X2=0.92 $Y2=1.37
cc_202 N_D_c_207_n N_CK_c_324_n 0.00175437f $X=0.725 $Y=1.37 $X2=0.92 $Y2=1.37
cc_203 D N_CK_c_324_n 0.00254088f $X=0.44 $Y=1.74 $X2=0.92 $Y2=1.37
cc_204 N_D_c_211_n N_CK_c_324_n 0.0178667f $X=1.115 $Y=1.34 $X2=0.92 $Y2=1.37
cc_205 N_D_c_212_n N_CK_c_324_n 0.0012142f $X=1.405 $Y=1.34 $X2=0.92 $Y2=1.37
cc_206 N_D_c_237_p N_CK_c_325_n 0.012157f $X=0.99 $Y=2.705 $X2=1.315 $Y2=2.11
cc_207 N_D_c_200_n N_CK_c_325_n 0.00112328f $X=1.26 $Y=1.34 $X2=1.315 $Y2=2.11
cc_208 N_D_c_211_n N_CK_c_325_n 0.00527669f $X=1.115 $Y=1.34 $X2=1.315 $Y2=2.11
cc_209 N_D_c_212_n N_CK_c_325_n 3.73987e-19 $X=1.405 $Y=1.34 $X2=1.315 $Y2=2.11
cc_210 N_D_c_199_n N_CK_c_326_n 0.0128995f $X=0.58 $Y=2.62 $X2=1.005 $Y2=2.11
cc_211 N_D_c_237_p N_CK_c_326_n 0.0056307f $X=0.99 $Y=2.705 $X2=1.005 $Y2=2.11
cc_212 N_D_c_199_n N_CK_c_328_n 0.00613815f $X=0.58 $Y=2.62 $X2=1.4 $Y2=2.11
cc_213 N_D_c_237_p N_CK_c_328_n 0.00103871f $X=0.99 $Y=2.705 $X2=1.4 $Y2=2.11
cc_214 N_D_c_199_n N_CK_c_330_n 0.00128303f $X=0.58 $Y=2.62 $X2=1.545 $Y2=2.11
cc_215 N_D_c_237_p N_CK_c_330_n 0.00146098f $X=0.99 $Y=2.705 $X2=1.545 $Y2=2.11
cc_216 N_D_M1013_g N_A_157_349#_M1011_g 0.067398f $X=0.5 $Y=3.235 $X2=0.86
+ $Y2=3.235
cc_217 N_D_c_199_n N_A_157_349#_M1011_g 0.00440628f $X=0.58 $Y=2.62 $X2=0.86
+ $Y2=3.235
cc_218 N_D_c_237_p N_A_157_349#_M1011_g 0.0174985f $X=0.99 $Y=2.705 $X2=0.86
+ $Y2=3.235
cc_219 N_D_c_200_n N_A_157_349#_c_458_n 0.00129448f $X=1.26 $Y=1.34 $X2=1.265
+ $Y2=1.825
cc_220 N_D_c_211_n N_A_157_349#_c_458_n 0.00253722f $X=1.115 $Y=1.34 $X2=1.265
+ $Y2=1.825
cc_221 N_D_c_194_n N_A_157_349#_c_459_n 0.067398f $X=0.44 $Y=1.74 $X2=0.935
+ $Y2=1.825
cc_222 N_D_c_203_n N_A_157_349#_c_459_n 0.00440628f $X=0.44 $Y=1.74 $X2=0.935
+ $Y2=1.825
cc_223 D N_A_157_349#_c_459_n 6.88464e-19 $X=0.44 $Y=1.74 $X2=0.935 $Y2=1.825
cc_224 N_D_c_211_n N_A_157_349#_c_459_n 5.21392e-19 $X=1.115 $Y=1.34 $X2=0.935
+ $Y2=1.825
cc_225 N_D_c_200_n N_A_157_349#_M1010_g 0.00957231f $X=1.26 $Y=1.34 $X2=1.46
+ $Y2=0.835
cc_226 N_D_c_208_n N_A_157_349#_M1010_g 0.0076805f $X=2.85 $Y=1.37 $X2=1.46
+ $Y2=0.835
cc_227 N_D_c_212_n N_A_157_349#_M1010_g 0.00345898f $X=1.405 $Y=1.34 $X2=1.46
+ $Y2=0.835
cc_228 N_D_c_194_n N_A_157_349#_c_463_n 0.00179364f $X=0.44 $Y=1.74 $X2=1.4
+ $Y2=1.74
cc_229 N_D_c_200_n N_A_157_349#_c_463_n 0.00189794f $X=1.26 $Y=1.34 $X2=1.4
+ $Y2=1.74
cc_230 N_D_c_212_n N_A_157_349#_c_463_n 6.44446e-19 $X=1.405 $Y=1.34 $X2=1.4
+ $Y2=1.74
cc_231 N_D_c_200_n N_A_157_349#_c_464_n 0.00647247f $X=1.26 $Y=1.34 $X2=1.4
+ $Y2=1.74
cc_232 N_D_c_212_n N_A_157_349#_c_464_n 0.00311227f $X=1.405 $Y=1.34 $X2=1.4
+ $Y2=1.74
cc_233 N_D_c_189_n N_A_157_349#_c_465_n 0.00707028f $X=3.2 $Y=1.205 $X2=2.465
+ $Y2=0.74
cc_234 N_D_M1000_g N_A_157_349#_c_465_n 0.00201047f $X=3.2 $Y=3.235 $X2=2.465
+ $Y2=0.74
cc_235 N_D_c_196_n N_A_157_349#_c_465_n 0.00361086f $X=3.2 $Y=1.37 $X2=2.465
+ $Y2=0.74
cc_236 N_D_c_201_n N_A_157_349#_c_465_n 0.00736723f $X=2.995 $Y=1.37 $X2=2.465
+ $Y2=0.74
cc_237 N_D_c_208_n N_A_157_349#_c_465_n 0.0227582f $X=2.85 $Y=1.37 $X2=2.465
+ $Y2=0.74
cc_238 N_D_c_213_n N_A_157_349#_c_465_n 0.00257549f $X=2.995 $Y=1.37 $X2=2.465
+ $Y2=0.74
cc_239 N_D_M1000_g N_A_157_349#_c_477_n 0.00699772f $X=3.2 $Y=3.235 $X2=2.465
+ $Y2=2.935
cc_240 N_D_M1000_g N_A_157_349#_c_469_n 0.0110692f $X=3.2 $Y=3.235 $X2=2.735
+ $Y2=2.62
cc_241 N_D_M1000_g N_A_157_349#_c_470_n 0.00299487f $X=3.2 $Y=3.235 $X2=2.735
+ $Y2=1.725
cc_242 N_D_c_208_n N_A_157_349#_c_470_n 0.00916047f $X=2.85 $Y=1.37 $X2=2.735
+ $Y2=1.725
cc_243 N_D_M1000_g N_A_157_349#_c_482_n 0.00340068f $X=3.2 $Y=3.235 $X2=2.735
+ $Y2=2.705
cc_244 N_D_c_200_n N_A_157_349#_c_471_n 3.69982e-19 $X=1.26 $Y=1.34 $X2=1.545
+ $Y2=1.725
cc_245 D N_A_157_349#_c_471_n 0.00827339f $X=0.44 $Y=1.74 $X2=1.545 $Y2=1.725
cc_246 N_D_c_212_n N_A_157_349#_c_471_n 0.0279898f $X=1.405 $Y=1.34 $X2=1.545
+ $Y2=1.725
cc_247 N_D_c_208_n N_A_157_349#_c_472_n 0.0251703f $X=2.85 $Y=1.37 $X2=2.465
+ $Y2=1.74
cc_248 N_D_c_208_n N_A_157_349#_c_473_n 0.0641247f $X=2.85 $Y=1.37 $X2=2.32
+ $Y2=1.74
cc_249 N_D_c_208_n N_A_349_89#_M1003_g 0.0105151f $X=2.85 $Y=1.37 $X2=1.82
+ $Y2=0.835
cc_250 N_D_c_212_n N_A_349_89#_M1003_g 2.70194e-19 $X=1.405 $Y=1.34 $X2=1.82
+ $Y2=0.835
cc_251 N_D_M1000_g N_A_349_89#_c_598_n 0.00462538f $X=3.2 $Y=3.235 $X2=4.1
+ $Y2=1.905
cc_252 N_D_c_208_n N_A_349_89#_c_603_n 7.90759e-19 $X=2.85 $Y=1.37 $X2=1.88
+ $Y2=1.74
cc_253 N_D_c_208_n N_A_349_89#_c_607_n 0.00517052f $X=2.85 $Y=1.37 $X2=1.882
+ $Y2=1.812
cc_254 N_D_c_189_n N_A_349_89#_c_609_n 0.0223047f $X=3.2 $Y=1.205 $X2=3.415
+ $Y2=0.74
cc_255 N_D_c_201_n N_A_349_89#_c_609_n 0.0115453f $X=2.995 $Y=1.37 $X2=3.415
+ $Y2=0.74
cc_256 N_D_c_213_n N_A_349_89#_c_609_n 0.00389142f $X=2.995 $Y=1.37 $X2=3.415
+ $Y2=0.74
cc_257 N_D_M1000_g N_A_349_89#_c_612_n 0.023277f $X=3.2 $Y=3.235 $X2=3.415
+ $Y2=2.935
cc_258 N_D_M1000_g N_A_349_89#_c_614_n 0.00244533f $X=3.2 $Y=3.235 $X2=3.415
+ $Y2=1.74
cc_259 N_D_M1000_g N_A_349_89#_c_617_n 0.0141612f $X=3.2 $Y=3.235 $X2=2.827
+ $Y2=2.395
cc_260 N_D_M1000_g N_A_349_89#_c_618_n 0.0162569f $X=3.2 $Y=3.235 $X2=3.9
+ $Y2=1.74
cc_261 N_D_c_201_n N_A_349_89#_c_618_n 7.4919e-19 $X=2.995 $Y=1.37 $X2=3.9
+ $Y2=1.74
cc_262 N_D_c_196_n N_A_349_89#_c_619_n 0.00415861f $X=3.2 $Y=1.37 $X2=2.9
+ $Y2=1.74
cc_263 N_D_c_201_n N_A_349_89#_c_619_n 0.00428868f $X=2.995 $Y=1.37 $X2=2.9
+ $Y2=1.74
cc_264 N_D_c_208_n N_A_349_89#_c_619_n 0.00830534f $X=2.85 $Y=1.37 $X2=2.9
+ $Y2=1.74
cc_265 N_D_c_213_n N_A_349_89#_c_619_n 0.0270542f $X=2.995 $Y=1.37 $X2=2.9
+ $Y2=1.74
cc_266 N_D_c_237_p A_115_521# 0.00473129f $X=0.99 $Y=2.705 $X2=0.575 $Y2=2.605
cc_267 N_D_c_310_p A_115_521# 0.00144354f $X=0.665 $Y=2.705 $X2=0.575 $Y2=2.605
cc_268 N_CK_M1014_g N_A_157_349#_M1011_g 0.0316011f $X=1.46 $Y=3.235 $X2=0.86
+ $Y2=3.235
cc_269 N_CK_c_317_n N_A_157_349#_M1011_g 0.0118393f $X=1.4 $Y=2.285 $X2=0.86
+ $Y2=3.235
cc_270 N_CK_c_324_n N_A_157_349#_M1011_g 0.00360955f $X=0.92 $Y=1.37 $X2=0.86
+ $Y2=3.235
cc_271 N_CK_c_326_n N_A_157_349#_M1011_g 0.0079407f $X=1.005 $Y=2.11 $X2=0.86
+ $Y2=3.235
cc_272 N_CK_c_328_n N_A_157_349#_M1011_g 0.00128351f $X=1.4 $Y=2.11 $X2=0.86
+ $Y2=3.235
cc_273 N_CK_c_330_n N_A_157_349#_M1011_g 4.61617e-19 $X=1.545 $Y=2.11 $X2=0.86
+ $Y2=3.235
cc_274 N_CK_c_324_n N_A_157_349#_c_458_n 0.00679428f $X=0.92 $Y=1.37 $X2=1.265
+ $Y2=1.825
cc_275 N_CK_c_325_n N_A_157_349#_c_458_n 0.00857512f $X=1.315 $Y=2.11 $X2=1.265
+ $Y2=1.825
cc_276 N_CK_c_330_n N_A_157_349#_c_458_n 0.00125393f $X=1.545 $Y=2.11 $X2=1.265
+ $Y2=1.825
cc_277 N_CK_c_313_n N_A_157_349#_c_459_n 0.0184383f $X=0.92 $Y=1.37 $X2=0.935
+ $Y2=1.825
cc_278 N_CK_c_324_n N_A_157_349#_c_459_n 0.00329856f $X=0.92 $Y=1.37 $X2=0.935
+ $Y2=1.825
cc_279 N_CK_c_313_n N_A_157_349#_M1010_g 0.013138f $X=0.92 $Y=1.37 $X2=1.46
+ $Y2=0.835
cc_280 N_CK_c_314_n N_A_157_349#_M1010_g 0.0152516f $X=0.92 $Y=1.205 $X2=1.46
+ $Y2=0.835
cc_281 N_CK_c_324_n N_A_157_349#_M1010_g 0.00166016f $X=0.92 $Y=1.37 $X2=1.46
+ $Y2=0.835
cc_282 N_CK_c_317_n N_A_157_349#_c_463_n 0.017377f $X=1.4 $Y=2.285 $X2=1.4
+ $Y2=1.74
cc_283 N_CK_c_324_n N_A_157_349#_c_463_n 0.00211698f $X=0.92 $Y=1.37 $X2=1.4
+ $Y2=1.74
cc_284 N_CK_c_328_n N_A_157_349#_c_463_n 0.00108353f $X=1.4 $Y=2.11 $X2=1.4
+ $Y2=1.74
cc_285 N_CK_c_317_n N_A_157_349#_c_464_n 7.72371e-19 $X=1.4 $Y=2.285 $X2=1.4
+ $Y2=1.74
cc_286 N_CK_c_324_n N_A_157_349#_c_464_n 0.00780691f $X=0.92 $Y=1.37 $X2=1.4
+ $Y2=1.74
cc_287 N_CK_c_325_n N_A_157_349#_c_464_n 0.00448992f $X=1.315 $Y=2.11 $X2=1.4
+ $Y2=1.74
cc_288 N_CK_c_328_n N_A_157_349#_c_464_n 0.00979766f $X=1.4 $Y=2.11 $X2=1.4
+ $Y2=1.74
cc_289 N_CK_c_329_n N_A_157_349#_c_464_n 5.17303e-19 $X=2.25 $Y=2.11 $X2=1.4
+ $Y2=1.74
cc_290 N_CK_c_330_n N_A_157_349#_c_464_n 0.00182452f $X=1.545 $Y=2.11 $X2=1.4
+ $Y2=1.74
cc_291 N_CK_c_318_n N_A_157_349#_c_465_n 0.00729529f $X=2.277 $Y=1.205 $X2=2.465
+ $Y2=0.74
cc_292 N_CK_c_323_n N_A_157_349#_c_465_n 0.0118432f $X=2.277 $Y=1.355 $X2=2.465
+ $Y2=0.74
cc_293 N_CK_c_311_n N_A_157_349#_c_469_n 0.00318866f $X=2.25 $Y=2.45 $X2=2.735
+ $Y2=2.62
cc_294 N_CK_M1008_g N_A_157_349#_c_469_n 0.00395773f $X=2.25 $Y=3.235 $X2=2.735
+ $Y2=2.62
cc_295 N_CK_c_312_n N_A_157_349#_c_469_n 0.00643904f $X=2.305 $Y=2.12 $X2=2.735
+ $Y2=2.62
cc_296 N_CK_c_327_n N_A_157_349#_c_469_n 0.0277441f $X=2.395 $Y=2.11 $X2=2.735
+ $Y2=2.62
cc_297 CK N_A_157_349#_c_469_n 0.00256489f $X=2.395 $Y=2.11 $X2=2.735 $Y2=2.62
cc_298 N_CK_c_311_n N_A_157_349#_c_470_n 0.0016621f $X=2.25 $Y=2.45 $X2=2.735
+ $Y2=1.725
cc_299 N_CK_c_312_n N_A_157_349#_c_470_n 0.00536103f $X=2.305 $Y=2.12 $X2=2.735
+ $Y2=1.725
cc_300 N_CK_c_327_n N_A_157_349#_c_470_n 0.00607622f $X=2.395 $Y=2.11 $X2=2.735
+ $Y2=1.725
cc_301 CK N_A_157_349#_c_470_n 7.74944e-19 $X=2.395 $Y=2.11 $X2=2.735 $Y2=1.725
cc_302 N_CK_c_311_n N_A_157_349#_c_482_n 0.00233394f $X=2.25 $Y=2.45 $X2=2.735
+ $Y2=2.705
cc_303 N_CK_c_327_n N_A_157_349#_c_482_n 0.00601935f $X=2.395 $Y=2.11 $X2=2.735
+ $Y2=2.705
cc_304 N_CK_c_324_n N_A_157_349#_c_471_n 0.00321055f $X=0.92 $Y=1.37 $X2=1.545
+ $Y2=1.725
cc_305 N_CK_c_325_n N_A_157_349#_c_471_n 6.0961e-19 $X=1.315 $Y=2.11 $X2=1.545
+ $Y2=1.725
cc_306 N_CK_c_328_n N_A_157_349#_c_471_n 4.76324e-19 $X=1.4 $Y=2.11 $X2=1.545
+ $Y2=1.725
cc_307 N_CK_c_330_n N_A_157_349#_c_471_n 0.0296305f $X=1.545 $Y=2.11 $X2=1.545
+ $Y2=1.725
cc_308 N_CK_c_311_n N_A_157_349#_c_472_n 2.36275e-19 $X=2.25 $Y=2.45 $X2=2.465
+ $Y2=1.74
cc_309 N_CK_c_312_n N_A_157_349#_c_472_n 0.00216028f $X=2.305 $Y=2.12 $X2=2.465
+ $Y2=1.74
cc_310 N_CK_c_327_n N_A_157_349#_c_472_n 0.00129914f $X=2.395 $Y=2.11 $X2=2.465
+ $Y2=1.74
cc_311 CK N_A_157_349#_c_472_n 0.0226506f $X=2.395 $Y=2.11 $X2=2.465 $Y2=1.74
cc_312 N_CK_c_312_n N_A_157_349#_c_473_n 0.00278025f $X=2.305 $Y=2.12 $X2=2.32
+ $Y2=1.74
cc_313 N_CK_c_323_n N_A_157_349#_c_473_n 2.64649e-19 $X=2.277 $Y=1.355 $X2=2.32
+ $Y2=1.74
cc_314 N_CK_c_329_n N_A_157_349#_c_473_n 0.0538111f $X=2.25 $Y=2.11 $X2=2.32
+ $Y2=1.74
cc_315 CK N_A_157_349#_c_473_n 0.00582134f $X=2.395 $Y=2.11 $X2=2.32 $Y2=1.74
cc_316 N_CK_c_312_n N_A_349_89#_M1003_g 0.00866378f $X=2.305 $Y=2.12 $X2=1.82
+ $Y2=0.835
cc_317 N_CK_c_318_n N_A_349_89#_M1003_g 0.0243817f $X=2.277 $Y=1.205 $X2=1.82
+ $Y2=0.835
cc_318 N_CK_c_311_n N_A_349_89#_M1015_g 0.0421262f $X=2.25 $Y=2.45 $X2=1.82
+ $Y2=3.235
cc_319 N_CK_c_312_n N_A_349_89#_M1015_g 0.0139901f $X=2.305 $Y=2.12 $X2=1.82
+ $Y2=3.235
cc_320 N_CK_c_317_n N_A_349_89#_M1015_g 0.113563f $X=1.4 $Y=2.285 $X2=1.82
+ $Y2=3.235
cc_321 N_CK_c_327_n N_A_349_89#_M1015_g 5.87562e-19 $X=2.395 $Y=2.11 $X2=1.82
+ $Y2=3.235
cc_322 N_CK_c_328_n N_A_349_89#_M1015_g 0.0022769f $X=1.4 $Y=2.11 $X2=1.82
+ $Y2=3.235
cc_323 N_CK_c_329_n N_A_349_89#_M1015_g 0.00269314f $X=2.25 $Y=2.11 $X2=1.82
+ $Y2=3.235
cc_324 N_CK_c_330_n N_A_349_89#_M1015_g 0.00113587f $X=1.545 $Y=2.11 $X2=1.82
+ $Y2=3.235
cc_325 N_CK_c_312_n N_A_349_89#_c_603_n 0.0205813f $X=2.305 $Y=2.12 $X2=1.88
+ $Y2=1.74
cc_326 N_CK_c_329_n N_A_349_89#_c_603_n 7.38456e-19 $X=2.25 $Y=2.11 $X2=1.88
+ $Y2=1.74
cc_327 N_CK_c_312_n N_A_349_89#_c_607_n 8.19109e-19 $X=2.305 $Y=2.12 $X2=1.882
+ $Y2=1.812
cc_328 N_CK_c_311_n N_A_349_89#_c_608_n 0.00276728f $X=2.25 $Y=2.45 $X2=1.88
+ $Y2=2.48
cc_329 N_CK_c_312_n N_A_349_89#_c_608_n 0.00446139f $X=2.305 $Y=2.12 $X2=1.88
+ $Y2=2.48
cc_330 N_CK_c_317_n N_A_349_89#_c_608_n 0.00225599f $X=1.4 $Y=2.285 $X2=1.88
+ $Y2=2.48
cc_331 N_CK_c_327_n N_A_349_89#_c_608_n 0.0149594f $X=2.395 $Y=2.11 $X2=1.88
+ $Y2=2.48
cc_332 N_CK_c_328_n N_A_349_89#_c_608_n 0.0150983f $X=1.4 $Y=2.11 $X2=1.88
+ $Y2=2.48
cc_333 N_CK_c_329_n N_A_349_89#_c_608_n 0.014171f $X=2.25 $Y=2.11 $X2=1.88
+ $Y2=2.48
cc_334 N_CK_c_330_n N_A_349_89#_c_608_n 0.00206546f $X=1.545 $Y=2.11 $X2=1.88
+ $Y2=2.48
cc_335 CK N_A_349_89#_c_608_n 0.00191287f $X=2.395 $Y=2.11 $X2=1.88 $Y2=2.48
cc_336 N_CK_c_311_n N_A_349_89#_c_615_n 0.00433056f $X=2.25 $Y=2.45 $X2=2.755
+ $Y2=2.48
cc_337 N_CK_M1008_g N_A_349_89#_c_615_n 0.00888384f $X=2.25 $Y=3.235 $X2=2.755
+ $Y2=2.48
cc_338 N_CK_c_327_n N_A_349_89#_c_615_n 0.00642492f $X=2.395 $Y=2.11 $X2=2.755
+ $Y2=2.48
cc_339 N_CK_c_329_n N_A_349_89#_c_615_n 0.0190773f $X=2.25 $Y=2.11 $X2=2.755
+ $Y2=2.48
cc_340 CK N_A_349_89#_c_615_n 0.025144f $X=2.395 $Y=2.11 $X2=2.755 $Y2=2.48
cc_341 N_CK_c_311_n N_A_349_89#_c_616_n 4.83733e-19 $X=2.25 $Y=2.45 $X2=2.025
+ $Y2=2.48
cc_342 N_CK_M1008_g N_A_349_89#_c_616_n 4.63789e-19 $X=2.25 $Y=3.235 $X2=2.025
+ $Y2=2.48
cc_343 N_CK_c_317_n N_A_349_89#_c_616_n 0.00405956f $X=1.4 $Y=2.285 $X2=2.025
+ $Y2=2.48
cc_344 N_CK_c_327_n N_A_349_89#_c_616_n 7.97287e-19 $X=2.395 $Y=2.11 $X2=2.025
+ $Y2=2.48
cc_345 N_CK_c_328_n N_A_349_89#_c_616_n 0.0025579f $X=1.4 $Y=2.11 $X2=2.025
+ $Y2=2.48
cc_346 N_CK_c_329_n N_A_349_89#_c_616_n 0.0252583f $X=2.25 $Y=2.11 $X2=2.025
+ $Y2=2.48
cc_347 N_CK_c_327_n N_A_349_89#_c_617_n 0.00120049f $X=2.395 $Y=2.11 $X2=2.827
+ $Y2=2.395
cc_348 CK N_A_349_89#_c_617_n 0.0189169f $X=2.395 $Y=2.11 $X2=2.827 $Y2=2.395
cc_349 N_A_157_349#_M1010_g N_A_349_89#_M1003_g 0.0464104f $X=1.46 $Y=0.835
+ $X2=1.82 $Y2=0.835
cc_350 N_A_157_349#_c_463_n N_A_349_89#_c_603_n 0.0464104f $X=1.4 $Y=1.74
+ $X2=1.88 $Y2=1.74
cc_351 N_A_157_349#_c_464_n N_A_349_89#_c_603_n 8.11121e-19 $X=1.4 $Y=1.74
+ $X2=1.88 $Y2=1.74
cc_352 N_A_157_349#_c_470_n N_A_349_89#_c_603_n 6.38549e-19 $X=2.735 $Y=1.725
+ $X2=1.88 $Y2=1.74
cc_353 N_A_157_349#_c_471_n N_A_349_89#_c_603_n 9.00828e-19 $X=1.545 $Y=1.725
+ $X2=1.88 $Y2=1.74
cc_354 N_A_157_349#_c_472_n N_A_349_89#_c_603_n 4.49351e-19 $X=2.465 $Y=1.74
+ $X2=1.88 $Y2=1.74
cc_355 N_A_157_349#_c_473_n N_A_349_89#_c_603_n 0.00295157f $X=2.32 $Y=1.74
+ $X2=1.88 $Y2=1.74
cc_356 N_A_157_349#_c_463_n N_A_349_89#_c_607_n 7.47762e-19 $X=1.4 $Y=1.74
+ $X2=1.882 $Y2=1.812
cc_357 N_A_157_349#_c_464_n N_A_349_89#_c_607_n 0.0079274f $X=1.4 $Y=1.74
+ $X2=1.882 $Y2=1.812
cc_358 N_A_157_349#_c_465_n N_A_349_89#_c_607_n 0.00183874f $X=2.465 $Y=0.74
+ $X2=1.882 $Y2=1.812
cc_359 N_A_157_349#_c_470_n N_A_349_89#_c_607_n 0.00400058f $X=2.735 $Y=1.725
+ $X2=1.882 $Y2=1.812
cc_360 N_A_157_349#_c_471_n N_A_349_89#_c_607_n 0.00135239f $X=1.545 $Y=1.725
+ $X2=1.882 $Y2=1.812
cc_361 N_A_157_349#_c_472_n N_A_349_89#_c_607_n 0.00102352f $X=2.465 $Y=1.74
+ $X2=1.882 $Y2=1.812
cc_362 N_A_157_349#_c_473_n N_A_349_89#_c_607_n 0.0115044f $X=2.32 $Y=1.74
+ $X2=1.882 $Y2=1.812
cc_363 N_A_157_349#_c_463_n N_A_349_89#_c_608_n 5.35826e-19 $X=1.4 $Y=1.74
+ $X2=1.88 $Y2=2.48
cc_364 N_A_157_349#_c_464_n N_A_349_89#_c_608_n 6.26362e-19 $X=1.4 $Y=1.74
+ $X2=1.88 $Y2=2.48
cc_365 N_A_157_349#_c_470_n N_A_349_89#_c_608_n 2.40837e-19 $X=2.735 $Y=1.725
+ $X2=1.88 $Y2=2.48
cc_366 N_A_157_349#_c_471_n N_A_349_89#_c_608_n 0.00136024f $X=1.545 $Y=1.725
+ $X2=1.88 $Y2=2.48
cc_367 N_A_157_349#_c_472_n N_A_349_89#_c_608_n 0.0012974f $X=2.465 $Y=1.74
+ $X2=1.88 $Y2=2.48
cc_368 N_A_157_349#_c_470_n N_A_349_89#_c_609_n 0.00107657f $X=2.735 $Y=1.725
+ $X2=3.415 $Y2=0.74
cc_369 N_A_157_349#_c_469_n N_A_349_89#_c_612_n 0.0168304f $X=2.735 $Y=2.62
+ $X2=3.415 $Y2=2.935
cc_370 N_A_157_349#_c_470_n N_A_349_89#_c_614_n 0.0038359f $X=2.735 $Y=1.725
+ $X2=3.415 $Y2=1.74
cc_371 N_A_157_349#_c_469_n N_A_349_89#_c_615_n 0.0136501f $X=2.735 $Y=2.62
+ $X2=2.755 $Y2=2.48
cc_372 N_A_157_349#_c_470_n N_A_349_89#_c_615_n 0.0020334f $X=2.735 $Y=1.725
+ $X2=2.755 $Y2=2.48
cc_373 N_A_157_349#_c_482_n N_A_349_89#_c_615_n 0.0134665f $X=2.735 $Y=2.705
+ $X2=2.755 $Y2=2.48
cc_374 N_A_157_349#_c_472_n N_A_349_89#_c_615_n 0.00360662f $X=2.465 $Y=1.74
+ $X2=2.755 $Y2=2.48
cc_375 N_A_157_349#_c_469_n N_A_349_89#_c_617_n 0.0185071f $X=2.735 $Y=2.62
+ $X2=2.827 $Y2=2.395
cc_376 N_A_157_349#_c_470_n N_A_349_89#_c_619_n 0.00779877f $X=2.735 $Y=1.725
+ $X2=2.9 $Y2=1.74
cc_377 N_A_157_349#_c_472_n N_A_349_89#_c_619_n 0.0198607f $X=2.465 $Y=1.74
+ $X2=2.9 $Y2=1.74
cc_378 N_A_349_89#_c_598_n N_ON_M1009_g 0.0154242f $X=4.1 $Y=1.905 $X2=4.58
+ $Y2=0.835
cc_379 N_A_349_89#_M1007_g N_ON_M1009_g 0.0253161f $X=4.15 $Y=0.835 $X2=4.58
+ $Y2=0.835
cc_380 N_A_349_89#_c_613_n N_ON_M1009_g 6.49773e-19 $X=4.035 $Y=1.74 $X2=4.58
+ $Y2=0.835
cc_381 N_A_349_89#_c_605_n N_ON_M1001_g 0.00624123f $X=4.125 $Y=2.36 $X2=4.58
+ $Y2=3.235
cc_382 N_A_349_89#_c_606_n N_ON_M1001_g 0.0506335f $X=4.125 $Y=2.49 $X2=4.58
+ $Y2=3.235
cc_383 N_A_349_89#_c_598_n N_ON_c_763_n 0.0212294f $X=4.1 $Y=1.905 $X2=4.52
+ $Y2=2.015
cc_384 N_A_349_89#_c_598_n N_ON_c_764_n 0.00188672f $X=4.1 $Y=1.905 $X2=3.935
+ $Y2=0.74
cc_385 N_A_349_89#_M1007_g N_ON_c_764_n 0.00981805f $X=4.15 $Y=0.835 $X2=3.935
+ $Y2=0.74
cc_386 N_A_349_89#_c_609_n N_ON_c_764_n 0.0322441f $X=3.415 $Y=0.74 $X2=3.935
+ $Y2=0.74
cc_387 N_A_349_89#_c_598_n N_ON_c_767_n 0.00289364f $X=4.1 $Y=1.905 $X2=3.935
+ $Y2=2.195
cc_388 N_A_349_89#_c_612_n N_ON_c_767_n 0.00525727f $X=3.415 $Y=2.935 $X2=3.935
+ $Y2=2.195
cc_389 N_A_349_89#_c_613_n N_ON_c_767_n 0.0101349f $X=4.035 $Y=1.74 $X2=3.935
+ $Y2=2.195
cc_390 N_A_349_89#_c_620_n N_ON_c_767_n 3.37612e-19 $X=4.035 $Y=1.74 $X2=3.935
+ $Y2=2.195
cc_391 N_A_349_89#_c_605_n N_ON_c_768_n 0.0120965f $X=4.125 $Y=2.36 $X2=3.935
+ $Y2=3.615
cc_392 N_A_349_89#_c_606_n N_ON_c_768_n 0.0210894f $X=4.125 $Y=2.49 $X2=3.935
+ $Y2=3.615
cc_393 N_A_349_89#_c_612_n N_ON_c_768_n 0.0721092f $X=3.415 $Y=2.935 $X2=3.935
+ $Y2=3.615
cc_394 N_A_349_89#_c_598_n N_ON_c_769_n 0.0192889f $X=4.1 $Y=1.905 $X2=4.43
+ $Y2=1.4
cc_395 N_A_349_89#_c_613_n N_ON_c_769_n 0.0110497f $X=4.035 $Y=1.74 $X2=4.43
+ $Y2=1.4
cc_396 N_A_349_89#_c_620_n N_ON_c_769_n 0.00387586f $X=4.035 $Y=1.74 $X2=4.43
+ $Y2=1.4
cc_397 N_A_349_89#_c_598_n N_ON_c_771_n 0.00308111f $X=4.1 $Y=1.905 $X2=4.02
+ $Y2=1.4
cc_398 N_A_349_89#_c_609_n N_ON_c_771_n 0.00869401f $X=3.415 $Y=0.74 $X2=4.02
+ $Y2=1.4
cc_399 N_A_349_89#_c_613_n N_ON_c_771_n 0.0120752f $X=4.035 $Y=1.74 $X2=4.02
+ $Y2=1.4
cc_400 N_A_349_89#_c_618_n N_ON_c_771_n 0.00132729f $X=3.9 $Y=1.74 $X2=4.02
+ $Y2=1.4
cc_401 N_A_349_89#_c_620_n N_ON_c_771_n 0.00306734f $X=4.035 $Y=1.74 $X2=4.02
+ $Y2=1.4
cc_402 N_A_349_89#_c_598_n N_ON_c_772_n 2.65797e-19 $X=4.1 $Y=1.905 $X2=4.435
+ $Y2=2.11
cc_403 N_A_349_89#_c_605_n N_ON_c_772_n 0.0141863f $X=4.125 $Y=2.36 $X2=4.435
+ $Y2=2.11
cc_404 N_A_349_89#_c_606_n N_ON_c_772_n 0.00208656f $X=4.125 $Y=2.49 $X2=4.435
+ $Y2=2.11
cc_405 N_A_349_89#_c_613_n N_ON_c_772_n 0.00957264f $X=4.035 $Y=1.74 $X2=4.435
+ $Y2=2.11
cc_406 N_A_349_89#_c_620_n N_ON_c_772_n 0.00261089f $X=4.035 $Y=1.74 $X2=4.435
+ $Y2=2.11
cc_407 N_A_349_89#_c_598_n N_ON_c_773_n 0.00356545f $X=4.1 $Y=1.905 $X2=4.517
+ $Y2=1.658
cc_408 N_A_349_89#_c_613_n N_ON_c_773_n 0.00537589f $X=4.035 $Y=1.74 $X2=4.517
+ $Y2=1.658
cc_409 N_A_349_89#_c_620_n N_ON_c_773_n 0.00199559f $X=4.035 $Y=1.74 $X2=4.517
+ $Y2=1.658
cc_410 N_A_349_89#_c_598_n N_ON_c_774_n 0.001785f $X=4.1 $Y=1.905 $X2=4.52
+ $Y2=2.015
cc_411 N_A_349_89#_c_613_n N_ON_c_774_n 0.004679f $X=4.035 $Y=1.74 $X2=4.52
+ $Y2=2.015
cc_412 N_A_349_89#_c_620_n N_ON_c_774_n 0.00189693f $X=4.035 $Y=1.74 $X2=4.52
+ $Y2=2.015
cc_413 N_A_349_89#_c_598_n ON 0.00197254f $X=4.1 $Y=1.905 $X2=3.935 $Y2=2.11
cc_414 N_A_349_89#_c_605_n ON 0.0039793f $X=4.125 $Y=2.36 $X2=3.935 $Y2=2.11
cc_415 N_A_349_89#_c_612_n ON 0.00761812f $X=3.415 $Y=2.935 $X2=3.935 $Y2=2.11
cc_416 N_A_349_89#_c_613_n ON 0.00222181f $X=4.035 $Y=1.74 $X2=3.935 $Y2=2.11
cc_417 N_A_349_89#_c_618_n ON 0.0192933f $X=3.9 $Y=1.74 $X2=3.935 $Y2=2.11
cc_418 N_A_349_89#_c_620_n ON 0.0183431f $X=4.035 $Y=1.74 $X2=3.935 $Y2=2.11
cc_419 N_A_349_89#_c_606_n Q 0.00101257f $X=4.125 $Y=2.49 $X2=4.795 $Y2=2.48
cc_420 N_ON_M1009_g N_Q_c_839_n 0.0054637f $X=4.58 $Y=0.835 $X2=4.827 $Y2=1.155
cc_421 N_ON_M1001_g N_Q_c_840_n 0.0237707f $X=4.58 $Y=3.235 $X2=4.795 $Y2=2.48
cc_422 N_ON_M1009_g N_Q_c_841_n 0.0314212f $X=4.58 $Y=0.835 $X2=4.827 $Y2=2.395
cc_423 N_ON_c_769_n N_Q_c_841_n 0.0135849f $X=4.43 $Y=1.4 $X2=4.827 $Y2=2.395
cc_424 N_ON_c_772_n N_Q_c_841_n 0.0135427f $X=4.435 $Y=2.11 $X2=4.827 $Y2=2.395
cc_425 N_ON_c_773_n N_Q_c_841_n 0.0380597f $X=4.517 $Y=1.658 $X2=4.827 $Y2=2.395
cc_426 N_ON_M1001_g Q 0.0138443f $X=4.58 $Y=3.235 $X2=4.795 $Y2=2.48
cc_427 N_ON_c_768_n Q 0.00547636f $X=3.935 $Y=3.615 $X2=4.795 $Y2=2.48
cc_428 N_ON_c_772_n Q 0.00264943f $X=4.435 $Y=2.11 $X2=4.795 $Y2=2.48
