* File: sky130_osu_sc_18T_ls__ndlat_l.pex.spice
* Created: Thu Mar 10 13:45:31 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%GND 1 2 3 49 51 58 60 70 72 82 95 97 99
+ 101 103 107
r105 105 107 0.00465721 $w=3.05e-07 $l=1e-08 $layer=MET1_cond $X=4.42 $Y=0.152
+ $X2=4.43 $Y2=0.152
r106 103 105 0.323676 $w=3.05e-07 $l=6.95e-07 $layer=MET1_cond $X=3.725 $Y=0.152
+ $X2=4.42 $Y2=0.152
r107 101 103 0.312033 $w=3.05e-07 $l=6.7e-07 $layer=MET1_cond $X=3.055 $Y=0.152
+ $X2=3.725 $Y2=0.152
r108 99 101 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=2.375 $Y=0.152
+ $X2=3.055 $Y2=0.152
r109 97 99 0.321348 $w=3.05e-07 $l=6.9e-07 $layer=MET1_cond $X=1.685 $Y=0.152
+ $X2=2.375 $Y2=0.152
r110 95 97 0.309705 $w=3.05e-07 $l=6.65e-07 $layer=MET1_cond $X=1.02 $Y=0.152
+ $X2=1.685 $Y2=0.152
r111 80 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.365 $Y=0.305
+ $X2=4.365 $Y2=0.865
r112 73 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.152
+ $X2=2.895 $Y2=0.152
r113 68 87 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.895 $Y=0.305
+ $X2=2.895 $Y2=0.152
r114 68 70 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.895 $Y=0.305
+ $X2=2.895 $Y2=0.825
r115 61 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.152
+ $X2=1.145 $Y2=0.152
r116 60 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.152
+ $X2=2.895 $Y2=0.152
r117 56 86 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.145 $Y=0.305
+ $X2=1.145 $Y2=0.152
r118 56 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.145 $Y=0.305
+ $X2=1.145 $Y2=0.825
r119 51 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.152
+ $X2=1.145 $Y2=0.152
r120 49 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r121 49 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r122 49 80 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.365 $Y2=0.305
r123 49 72 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.28 $Y2=0.152
r124 49 72 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.28 $Y2=0.152
r125 49 73 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=3.06 $Y=0.152 $X2=2.98
+ $Y2=0.152
r126 49 60 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.81 $Y2=0.152
r127 49 61 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.23 $Y2=0.152
r128 49 51 1.6 $w=3.05e-07 $l=4e-08 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=1.06
+ $Y2=0.152
r129 3 82 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.575 $X2=4.365 $Y2=0.865
r130 2 70 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.575 $X2=2.895 $Y2=0.825
r131 1 58 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.575 $X2=1.145 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%VDD 1 2 3 37 41 47 51 59 63 71 80 86 88
+ 90 94
r65 92 94 0.00232861 $w=3.05e-07 $l=5e-09 $layer=MET1_cond $X=4.42 $Y=6.507
+ $X2=4.425 $Y2=6.507
r66 90 92 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=3.735 $Y=6.507
+ $X2=4.42 $Y2=6.507
r67 88 90 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=3.055 $Y=6.507
+ $X2=3.735 $Y2=6.507
r68 86 88 0.314362 $w=3.05e-07 $l=6.75e-07 $layer=MET1_cond $X=2.38 $Y=6.507
+ $X2=3.055 $Y2=6.507
r69 83 86 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=1.02 $Y=6.507
+ $X2=2.38 $Y2=6.507
r70 80 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.42 $Y=6.47
+ $X2=4.42 $Y2=6.47
r71 71 74 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.365 $Y=4.465
+ $X2=4.365 $Y2=5.825
r72 69 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.365 $Y=6.355
+ $X2=4.365 $Y2=6.507
r73 69 74 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.365 $Y=6.355
+ $X2=4.365 $Y2=5.825
r74 66 68 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=6.507
+ $X2=3.74 $Y2=6.507
r75 64 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=6.507
+ $X2=2.895 $Y2=6.507
r76 64 66 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=2.98 $Y=6.507 $X2=3.06
+ $Y2=6.507
r77 63 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=6.507
+ $X2=4.365 $Y2=6.507
r78 63 68 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=4.28 $Y=6.507
+ $X2=3.74 $Y2=6.507
r79 59 62 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.895 $Y=3.455
+ $X2=2.895 $Y2=5.835
r80 57 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.895 $Y=6.355
+ $X2=2.895 $Y2=6.507
r81 57 62 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.895 $Y=6.355
+ $X2=2.895 $Y2=5.835
r82 54 56 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=6.507
+ $X2=2.38 $Y2=6.507
r83 52 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=6.507
+ $X2=1.145 $Y2=6.507
r84 52 54 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.23 $Y=6.507 $X2=1.7
+ $Y2=6.507
r85 51 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=6.507
+ $X2=2.895 $Y2=6.507
r86 51 56 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.81 $Y=6.507
+ $X2=2.38 $Y2=6.507
r87 47 50 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.145 $Y=3.795
+ $X2=1.145 $Y2=5.835
r88 45 77 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.145 $Y=6.355
+ $X2=1.145 $Y2=6.507
r89 45 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.145 $Y=6.355
+ $X2=1.145 $Y2=5.835
r90 43 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r91 41 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=6.507
+ $X2=1.145 $Y2=6.507
r92 41 43 1.6 $w=3.05e-07 $l=4e-08 $layer=LI1_cond $X=1.06 $Y=6.507 $X2=1.02
+ $Y2=6.507
r93 37 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r94 37 68 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r95 37 66 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r96 37 56 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r97 37 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r98 37 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r99 3 74 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=4.085 $X2=4.365 $Y2=5.825
r100 3 71 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=4.085 $X2=4.365 $Y2=4.465
r101 2 62 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.755
+ $Y=3.085 $X2=2.895 $Y2=5.835
r102 2 59 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.755
+ $Y=3.085 $X2=2.895 $Y2=3.455
r103 1 50 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=1.005 $Y=3.085 $X2=1.145 $Y2=5.835
r104 1 47 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=1.005 $Y=3.085 $X2=1.145 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_161_337# 1 3 13 16 18 19 21 22 23 24
+ 25 27 28 30 31 32 35 39
r82 39 41 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=2.02 $Y=3.455
+ $X2=2.02 $Y2=5.835
r83 37 39 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=2.02 $Y=3.27
+ $X2=2.02 $Y2=3.455
r84 33 35 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=2.02 $Y=1.345
+ $X2=2.02 $Y2=0.825
r85 31 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.85 $Y=1.43
+ $X2=2.02 $Y2=1.345
r86 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.85 $Y=1.43
+ $X2=1.57 $Y2=1.43
r87 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=1.515
+ $X2=1.57 $Y2=1.43
r88 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.485 $Y=1.515
+ $X2=1.485 $Y2=1.765
r89 27 37 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.85 $Y=3.185
+ $X2=2.02 $Y2=3.27
r90 27 28 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.85 $Y=3.185
+ $X2=1.025 $Y2=3.185
r91 26 44 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.025 $Y=1.85
+ $X2=0.94 $Y2=1.81
r92 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.4 $Y=1.85
+ $X2=1.485 $Y2=1.765
r93 25 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.4 $Y=1.85
+ $X2=1.025 $Y2=1.85
r94 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.94 $Y=3.1
+ $X2=1.025 $Y2=3.185
r95 23 44 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=1.935
+ $X2=0.94 $Y2=1.81
r96 23 24 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=0.94 $Y=1.935
+ $X2=0.94 $Y2=3.1
r97 21 22 56.3681 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=0.905 $Y=2.805
+ $X2=0.905 $Y2=2.975
r98 20 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.88 $Y=2.015
+ $X2=0.88 $Y2=2.805
r99 18 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.85 $X2=0.94 $Y2=1.85
r100 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.85
+ $X2=0.94 $Y2=2.015
r101 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.85
+ $X2=0.94 $Y2=1.685
r102 16 22 517.347 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=0.93 $Y=4.585
+ $X2=0.93 $Y2=2.975
r103 13 19 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.93 $Y=1.075
+ $X2=0.93 $Y2=1.685
r104 3 41 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.795
+ $Y=3.085 $X2=2.02 $Y2=5.835
r105 3 39 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.795
+ $Y=3.085 $X2=2.02 $Y2=3.455
r106 1 35 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.795
+ $Y=0.575 $X2=2.02 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%D 3 7 10 14 20
c51 7 0 1.64001e-19 $X=1.36 $Y=4.585
c52 3 0 1.3839e-19 $X=1.36 $Y=1.075
r53 20 23 0.00169837 $w=3.68e-07 $l=5e-09 $layer=MET1_cond $X=1.352 $Y=2.59
+ $X2=1.352 $Y2=2.595
r54 17 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.3 $Y=2.595 $X2=1.3
+ $Y2=2.595
r55 14 17 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.3 $Y=2.425 $X2=1.3
+ $Y2=2.595
r56 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.3
+ $Y=2.425 $X2=1.3 $Y2=2.425
r57 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=2.425
+ $X2=1.3 $Y2=2.59
r58 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=2.425
+ $X2=1.3 $Y2=2.26
r59 7 12 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=1.36 $Y=4.585
+ $X2=1.36 $Y2=2.59
r60 3 11 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.36 $Y=1.075
+ $X2=1.36 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%CK 3 7 8 10 13 15 18 22 23 25 26 30 31
+ 33 37 44 46 47 49
c123 44 0 9.95038e-20 $X=1.86 $Y=2.765
c124 31 0 1.3839e-19 $X=1.945 $Y=1.85
c125 30 0 1.64001e-19 $X=1.86 $Y=2.68
c126 25 0 1.9983e-19 $X=3.137 $Y=2.78
c127 18 0 1.47633e-20 $X=1.78 $Y=2.765
r128 47 49 0.0928211 $w=2.16e-07 $l=1.50997e-07 $layer=MET1_cond $X=2.41 $Y=1.85
+ $X2=2.26 $Y2=1.852
r129 46 53 0.101772 $w=2.27e-07 $l=1.71493e-07 $layer=MET1_cond $X=3.075 $Y=1.85
+ $X2=3.245 $Y2=1.847
r130 46 47 0.640317 $w=1.7e-07 $l=6.65e-07 $layer=MET1_cond $X=3.075 $Y=1.85
+ $X2=2.41 $Y2=1.85
r131 42 44 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.78 $Y=2.765
+ $X2=1.86 $Y2=2.765
r132 37 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.245 $Y=1.85
+ $X2=3.245 $Y2=1.85
r133 33 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.26 $Y=1.85
+ $X2=2.26 $Y2=1.85
r134 31 33 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.945 $Y=1.85
+ $X2=2.26 $Y2=1.85
r135 30 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=2.68
+ $X2=1.86 $Y2=2.765
r136 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.86 $Y=1.935
+ $X2=1.945 $Y2=1.85
r137 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.86 $Y=1.935
+ $X2=1.86 $Y2=2.68
r138 28 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.85 $X2=3.245 $Y2=1.85
r139 25 26 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=3.137 $Y=2.78
+ $X2=3.137 $Y2=2.93
r140 22 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.85 $X2=2.26 $Y2=1.85
r141 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.85
+ $X2=2.26 $Y2=1.685
r142 18 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=2.765 $X2=1.78 $Y2=2.765
r143 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=2.765
+ $X2=1.78 $Y2=2.93
r144 15 28 38.6212 $w=3.33e-07 $l=1.89222e-07 $layer=POLY_cond $X=3.165 $Y=2.015
+ $X2=3.217 $Y2=1.85
r145 15 25 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=3.165 $Y=2.015
+ $X2=3.165 $Y2=2.78
r146 13 26 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.11 $Y=4.585
+ $X2=3.11 $Y2=2.93
r147 8 28 41.516 $w=3.33e-07 $l=2.32422e-07 $layer=POLY_cond $X=3.11 $Y=1.665
+ $X2=3.217 $Y2=1.85
r148 8 10 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=1.075
r149 7 23 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.32 $Y=1.075
+ $X2=2.32 $Y2=1.685
r150 3 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.72 $Y=4.585
+ $X2=1.72 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_329_89# 1 3 11 13 14 19 22 23 26 33
+ 37 44 47 51 53 54 59
c124 54 0 1.47633e-20 $X=2.405 $Y=2.59
c125 22 0 1.2087e-19 $X=2.26 $Y=2.765
c126 13 0 9.95038e-20 $X=2.125 $Y=2.3
r127 54 56 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.405 $Y=2.59
+ $X2=2.26 $Y2=2.59
r128 53 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.18 $Y=2.59
+ $X2=3.325 $Y2=2.59
r129 53 54 0.746234 $w=1.7e-07 $l=7.75e-07 $layer=MET1_cond $X=3.18 $Y=2.59
+ $X2=2.405 $Y2=2.59
r130 49 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.325 $Y=2.27
+ $X2=3.595 $Y2=2.27
r131 45 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.325 $Y=1.42
+ $X2=3.595 $Y2=1.42
r132 44 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=2.185
+ $X2=3.595 $Y2=2.27
r133 43 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=1.505
+ $X2=3.595 $Y2=1.42
r134 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.595 $Y=1.505
+ $X2=3.595 $Y2=2.185
r135 39 41 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.325 $Y=3.455
+ $X2=3.325 $Y2=5.835
r136 37 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.325 $Y=2.59
+ $X2=3.325 $Y2=2.59
r137 37 39 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.325 $Y=2.59
+ $X2=3.325 $Y2=3.455
r138 35 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.355
+ $X2=3.325 $Y2=2.27
r139 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.325 $Y=2.355
+ $X2=3.325 $Y2=2.59
r140 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.335
+ $X2=3.325 $Y2=1.42
r141 31 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.325 $Y=1.335
+ $X2=3.325 $Y2=0.825
r142 26 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.26 $Y=2.59
+ $X2=2.26 $Y2=2.59
r143 26 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.26 $Y=2.59
+ $X2=2.26 $Y2=2.765
r144 22 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=2.765 $X2=2.26 $Y2=2.765
r145 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=2.765
+ $X2=2.26 $Y2=2.93
r146 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=2.765
+ $X2=2.26 $Y2=2.6
r147 19 24 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.32 $Y=4.585
+ $X2=2.32 $Y2=2.93
r148 15 23 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.2 $Y=2.375
+ $X2=2.2 $Y2=2.6
r149 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=2.3
+ $X2=2.2 $Y2=2.375
r150 13 14 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.125 $Y=2.3
+ $X2=1.795 $Y2=2.3
r151 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.72 $Y=2.225
+ $X2=1.795 $Y2=2.3
r152 9 11 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=1.72 $Y=2.225
+ $X2=1.72 $Y2=1.075
r153 3 41 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.185
+ $Y=3.085 $X2=3.325 $Y2=5.835
r154 3 39 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.185
+ $Y=3.085 $X2=3.325 $Y2=3.455
r155 1 33 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.185
+ $Y=0.575 $X2=3.325 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%A_118_115# 1 3 11 15 23 27 29 33 34 37
+ 38 39 43 46 50 55 60 66 69 74 75 79 82 84
c154 82 0 1.2087e-19 $X=2.595 $Y=2.22
c155 60 0 1.9983e-19 $X=4.035 $Y=2.22
c156 38 0 8.77106e-20 $X=4.125 $Y=3.855
c157 33 0 1.18035e-19 $X=4.035 $Y=2.22
r158 81 82 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.74 $Y=2.22
+ $X2=2.595 $Y2=2.22
r159 79 82 2.2896 $w=1.4e-07 $l=1.85e-06 $layer=MET1_cond $X=0.745 $Y=2.2
+ $X2=2.595 $Y2=2.2
r160 77 79 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.6 $Y=2.22
+ $X2=0.745 $Y2=2.22
r161 75 81 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=2.89 $Y=2.22
+ $X2=2.74 $Y2=2.22
r162 74 84 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.89 $Y=2.22
+ $X2=4.035 $Y2=2.22
r163 74 75 1.23762 $w=1.4e-07 $l=1e-06 $layer=MET1_cond $X=3.89 $Y=2.22 $X2=2.89
+ $Y2=2.22
r164 69 71 8.33135 $w=2.83e-07 $l=1.6e-07 $layer=LI1_cond $X=0.657 $Y=3.795
+ $X2=0.657 $Y2=3.955
r165 69 70 12.1728 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.657 $Y=3.795
+ $X2=0.657 $Y2=3.54
r166 64 66 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.6 $Y=1.395
+ $X2=0.715 $Y2=1.395
r167 60 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.035 $Y=2.22
+ $X2=4.035 $Y2=2.22
r168 55 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.74 $Y=2.22
+ $X2=2.74 $Y2=2.22
r169 50 52 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=5.835
r170 50 71 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=3.955
r171 44 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=1.31
+ $X2=0.715 $Y2=1.395
r172 44 46 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.715 $Y=1.31
+ $X2=0.715 $Y2=0.825
r173 43 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.6 $Y=2.22 $X2=0.6
+ $Y2=2.22
r174 43 70 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.6 $Y=2.22
+ $X2=0.6 $Y2=3.54
r175 40 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=1.48 $X2=0.6
+ $Y2=1.395
r176 40 43 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.6 $Y=1.48 $X2=0.6
+ $Y2=2.22
r177 38 39 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=3.855
+ $X2=4.125 $Y2=4.005
r178 36 37 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=1.65
+ $X2=4.125 $Y2=1.8
r179 35 38 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=4.1 $Y=2.385
+ $X2=4.1 $Y2=3.855
r180 34 37 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.1 $Y=2.055
+ $X2=4.1 $Y2=1.8
r181 33 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=2.22 $X2=4.035 $Y2=2.22
r182 33 35 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.037 $Y=2.22
+ $X2=4.037 $Y2=2.385
r183 33 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.037 $Y=2.22
+ $X2=4.037 $Y2=2.055
r184 29 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=2.22 $X2=2.74 $Y2=2.22
r185 29 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=2.22
+ $X2=2.74 $Y2=2.385
r186 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=2.22
+ $X2=2.74 $Y2=2.055
r187 27 39 347.04 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=4.15 $Y=5.085
+ $X2=4.15 $Y2=4.005
r188 23 36 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=4.15 $Y=0.945
+ $X2=4.15 $Y2=1.65
r189 15 31 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=2.68 $Y=4.585
+ $X2=2.68 $Y2=2.385
r190 11 30 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.68 $Y=1.075
+ $X2=2.68 $Y2=2.055
r191 3 52 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.59
+ $Y=3.085 $X2=0.715 $Y2=5.835
r192 3 50 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.59
+ $Y=3.085 $X2=0.715 $Y2=4.135
r193 3 69 600 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=3.085 $X2=0.715 $Y2=3.795
r194 1 46 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.575 $X2=0.715 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c67 44 0 8.77106e-20 $X=3.94 $Y=3.96
c68 33 0 1.18035e-19 $X=4.435 $Y=1.85
r69 42 44 0.00296209 $w=2.11e-07 $l=5e-09 $layer=MET1_cond $X=3.935 $Y=3.96
+ $X2=3.94 $Y2=3.96
r70 38 40 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=4.52 $Y=3.68
+ $X2=4.52 $Y2=2.22
r71 37 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.52 $Y=1.935
+ $X2=4.52 $Y2=2.22
r72 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=3.765
+ $X2=4.52 $Y2=3.68
r73 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=3.765
+ $X2=4.02 $Y2=3.765
r74 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=1.85
+ $X2=4.52 $Y2=1.935
r75 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=1.85
+ $X2=4.02 $Y2=1.85
r76 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.935 $Y=4.465
+ $X2=3.935 $Y2=5.825
r77 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=3.96
+ $X2=3.935 $Y2=3.96
r78 27 29 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.935 $Y=3.96
+ $X2=3.935 $Y2=4.465
r79 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=3.85
+ $X2=4.02 $Y2=3.765
r80 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.935 $Y=3.85
+ $X2=3.935 $Y2=3.96
r81 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=1.765
+ $X2=4.02 $Y2=1.85
r82 21 23 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=3.935 $Y=1.765
+ $X2=3.935 $Y2=0.865
r83 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=2.22 $X2=4.52 $Y2=2.22
r84 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.22
+ $X2=4.52 $Y2=2.385
r85 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.22
+ $X2=4.52 $Y2=2.055
r86 15 20 1384.47 $w=1.5e-07 $l=2.7e-06 $layer=POLY_cond $X=4.58 $Y=5.085
+ $X2=4.58 $Y2=2.385
r87 11 19 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=4.58 $Y=0.945
+ $X2=4.58 $Y2=2.055
r88 3 31 240 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=3.81
+ $Y=4.085 $X2=3.935 $Y2=5.825
r89 3 29 240 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=3.81
+ $Y=4.085 $X2=3.935 $Y2=4.465
r90 1 23 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=3.81
+ $Y=0.575 $X2=3.935 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__NDLAT_L%Q 1 3 11 15 17 24 25 28
r19 24 25 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=4.86 $Y=1.335
+ $X2=4.86 $Y2=4.16
r20 23 24 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.827 $Y=1.165
+ $X2=4.827 $Y2=1.335
r21 17 19 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.795 $Y=4.465
+ $X2=4.795 $Y2=5.825
r22 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.795 $Y=4.33
+ $X2=4.795 $Y2=4.33
r23 15 25 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.827 $Y=4.33
+ $X2=4.827 $Y2=4.16
r24 15 17 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.795 $Y=4.33
+ $X2=4.795 $Y2=4.465
r25 11 23 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.795 $Y=0.865
+ $X2=4.795 $Y2=1.165
r26 3 19 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=4.655
+ $Y=4.085 $X2=4.795 $Y2=5.825
r27 3 17 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=4.655
+ $Y=4.085 $X2=4.795 $Y2=4.465
r28 1 11 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.575 $X2=4.795 $Y2=0.865
.ends

