* File: sky130_osu_sc_15T_ms__or2_l.pex.spice
* Created: Fri Nov 12 14:46:25 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__OR2_L%GND 1 2 21 25 27 35 42 44 47
r35 44 47 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r36 33 42 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r37 33 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.74
r38 27 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r39 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r40 21 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r41 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r42 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r43 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r44 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r45 2 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.74
r46 1 25 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_L%VDD 1 13 15 24 28 30 33
r25 30 33 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r26 22 28 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r27 22 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r28 20 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r29 17 20 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r30 15 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r31 15 20 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r32 13 20 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r33 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r34 1 24 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=3.565 $X2=1.12 $Y2=4.565
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_L%B 3 7 12 15 21
c29 15 0 1.87787e-19 $X=0.27 $Y=2.415
r30 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.7 $X2=0.27
+ $Y2=2.7
r31 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.415
+ $X2=0.27 $Y2=2.7
r32 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.415 $X2=0.27 $Y2=2.415
r33 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.415
+ $X2=0.475 $Y2=2.415
r34 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.58
+ $X2=0.475 $Y2=2.415
r35 5 7 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=0.475 $Y=2.58
+ $X2=0.475 $Y2=4.195
r36 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.25
+ $X2=0.475 $Y2=2.415
r37 1 3 725.564 $w=1.5e-07 $l=1.415e-06 $layer=POLY_cond $X=0.475 $Y=2.25
+ $X2=0.475 $Y2=0.835
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_L%A 3 7 10 14 20
r42 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=3.07
+ $X2=0.95 $Y2=3.07
r43 14 17 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=2.125
+ $X2=0.95 $Y2=3.07
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.125 $X2=0.95 $Y2=2.125
r45 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.125
+ $X2=0.95 $Y2=2.29
r46 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.125
+ $X2=0.95 $Y2=1.96
r47 7 12 976.819 $w=1.5e-07 $l=1.905e-06 $layer=POLY_cond $X=0.905 $Y=4.195
+ $X2=0.905 $Y2=2.29
r48 3 11 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=0.905 $Y=0.835
+ $X2=0.905 $Y2=1.96
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_L%A_27_713# 1 3 11 15 17 19 20 25 27 28 30
+ 33 37 39
c71 27 0 1.87787e-19 $X=0.525 $Y=3.37
r72 35 39 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.675
+ $X2=0.65 $Y2=1.675
r73 35 37 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.675
+ $X2=1.43 $Y2=1.675
r74 31 39 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.65 $Y2=1.675
r75 31 33 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.69 $Y2=0.74
r76 29 39 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.65 $Y2=1.675
r77 29 30 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=3.285
r78 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.37
+ $X2=0.61 $Y2=3.285
r79 27 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.37
+ $X2=0.345 $Y2=3.37
r80 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.345 $Y2=3.37
r81 23 25 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=4.565
r82 22 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.675 $X2=1.43 $Y2=1.675
r83 19 20 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.55
+ $X2=1.352 $Y2=2.7
r84 17 22 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.412 $Y2=1.675
r85 17 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=2.55
r86 15 20 766.585 $w=1.5e-07 $l=1.495e-06 $layer=POLY_cond $X=1.335 $Y=4.195
+ $X2=1.335 $Y2=2.7
r87 9 22 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.412 $Y2=1.675
r88 9 11 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.835
r89 3 25 600 $w=1.7e-07 $l=1.06066e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=3.565 $X2=0.26 $Y2=4.565
r90 1 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_L%Y 1 3 10 16 24 27 30
r34 22 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r35 22 24 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r36 21 27 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r37 21 24 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r38 16 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r39 16 19 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=4.565
r40 13 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r41 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.22
r42 3 19 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=3.565 $X2=1.55 $Y2=4.565
r43 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

