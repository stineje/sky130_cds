* File: sky130_osu_sc_12T_ms__or2_4.pxi.spice
* Created: Fri Nov 12 15:26:19 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__OR2_4%GND N_GND_M1003_s N_GND_M1000_d N_GND_M1009_s
+ N_GND_M1011_s N_GND_M1003_b N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p
+ N_GND_c_24_p N_GND_c_32_p N_GND_c_38_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_MS__OR2_4%GND
x_PM_SKY130_OSU_SC_12T_MS__OR2_4%VDD N_VDD_M1007_d N_VDD_M1005_d N_VDD_M1008_d
+ N_VDD_M1002_b N_VDD_c_78_p N_VDD_c_84_p N_VDD_c_91_p N_VDD_c_97_p
+ N_VDD_c_103_p N_VDD_c_108_p VDD N_VDD_c_79_p
+ PM_SKY130_OSU_SC_12T_MS__OR2_4%VDD
x_PM_SKY130_OSU_SC_12T_MS__OR2_4%B N_B_M1003_g N_B_M1002_g N_B_c_129_n
+ N_B_c_130_n B PM_SKY130_OSU_SC_12T_MS__OR2_4%B
x_PM_SKY130_OSU_SC_12T_MS__OR2_4%A N_A_M1000_g N_A_M1007_g N_A_c_157_n
+ N_A_c_158_n A PM_SKY130_OSU_SC_12T_MS__OR2_4%A
x_PM_SKY130_OSU_SC_12T_MS__OR2_4%A_27_521# N_A_27_521#_M1003_d
+ N_A_27_521#_M1002_s N_A_27_521#_M1001_g N_A_27_521#_c_231_n
+ N_A_27_521#_M1004_g N_A_27_521#_c_200_n N_A_27_521#_c_201_n
+ N_A_27_521#_M1009_g N_A_27_521#_c_236_n N_A_27_521#_M1005_g
+ N_A_27_521#_c_206_n N_A_27_521#_c_208_n N_A_27_521#_c_209_n
+ N_A_27_521#_M1010_g N_A_27_521#_c_243_n N_A_27_521#_M1006_g
+ N_A_27_521#_c_214_n N_A_27_521#_c_215_n N_A_27_521#_M1011_g
+ N_A_27_521#_c_248_n N_A_27_521#_M1008_g N_A_27_521#_c_220_n
+ N_A_27_521#_c_221_n N_A_27_521#_c_222_n N_A_27_521#_c_223_n
+ N_A_27_521#_c_255_n N_A_27_521#_c_259_n N_A_27_521#_c_261_n
+ N_A_27_521#_c_224_n N_A_27_521#_c_225_n N_A_27_521#_c_228_n
+ N_A_27_521#_c_230_n PM_SKY130_OSU_SC_12T_MS__OR2_4%A_27_521#
x_PM_SKY130_OSU_SC_12T_MS__OR2_4%Y N_Y_M1001_d N_Y_M1010_d N_Y_M1004_s
+ N_Y_M1006_s N_Y_c_334_n N_Y_c_338_n N_Y_c_339_n N_Y_c_343_n N_Y_c_344_n
+ N_Y_c_348_n Y N_Y_c_350_n N_Y_c_354_n N_Y_c_355_n N_Y_c_359_n
+ PM_SKY130_OSU_SC_12T_MS__OR2_4%Y
cc_1 N_GND_M1003_b N_B_M1003_g 0.083817f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_B_M1003_g 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_B_M1003_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.835
cc_4 N_GND_c_4_p N_B_M1003_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=0.835
cc_5 N_GND_M1003_b N_B_M1002_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_6 N_GND_M1003_b N_B_c_129_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.195
cc_7 N_GND_M1003_b N_B_c_130_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.195
cc_8 N_GND_M1003_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.48
cc_9 N_GND_M1003_b N_A_M1000_g 0.0440597f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.835
cc_10 N_GND_c_3_p N_A_M1000_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.835
cc_11 N_GND_c_11_p N_A_M1000_g 0.00308284f $X=1.12 $Y=0.755 $X2=0.905 $Y2=0.835
cc_12 N_GND_c_4_p N_A_M1000_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.905 $Y2=0.835
cc_13 N_GND_M1003_b N_A_M1007_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_14 N_GND_M1003_b N_A_c_157_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.905
cc_15 N_GND_M1003_b N_A_c_158_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.905
cc_16 N_GND_M1003_b N_A_27_521#_M1001_g 0.0207501f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.835
cc_17 N_GND_c_11_p N_A_27_521#_M1001_g 0.00308284f $X=1.12 $Y=0.755 $X2=1.335
+ $Y2=0.835
cc_18 N_GND_c_18_p N_A_27_521#_M1001_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.835
cc_19 N_GND_c_4_p N_A_27_521#_M1001_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.335
+ $Y2=0.835
cc_20 N_GND_M1003_b N_A_27_521#_c_200_n 0.0466273f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.33
cc_21 N_GND_M1003_b N_A_27_521#_c_201_n 0.00954592f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.405
cc_22 N_GND_M1003_b N_A_27_521#_M1009_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.835
cc_23 N_GND_c_18_p N_A_27_521#_M1009_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.835
cc_24 N_GND_c_24_p N_A_27_521#_M1009_g 0.00311745f $X=1.98 $Y=0.755 $X2=1.765
+ $Y2=0.835
cc_25 N_GND_c_4_p N_A_27_521#_M1009_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.765
+ $Y2=0.835
cc_26 N_GND_M1003_b N_A_27_521#_c_206_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.365
cc_27 N_GND_c_24_p N_A_27_521#_c_206_n 0.00256938f $X=1.98 $Y=0.755 $X2=2.12
+ $Y2=1.365
cc_28 N_GND_M1003_b N_A_27_521#_c_208_n 0.0439685f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.365
cc_29 N_GND_M1003_b N_A_27_521#_c_209_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.405
cc_30 N_GND_M1003_b N_A_27_521#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.835
cc_31 N_GND_c_24_p N_A_27_521#_M1010_g 0.00311745f $X=1.98 $Y=0.755 $X2=2.195
+ $Y2=0.835
cc_32 N_GND_c_32_p N_A_27_521#_M1010_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.835
cc_33 N_GND_c_4_p N_A_27_521#_M1010_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.195
+ $Y2=0.835
cc_34 N_GND_M1003_b N_A_27_521#_c_214_n 0.0369419f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.365
cc_35 N_GND_M1003_b N_A_27_521#_c_215_n 0.0268552f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.405
cc_36 N_GND_M1003_b N_A_27_521#_M1011_g 0.0264941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.835
cc_37 N_GND_c_32_p N_A_27_521#_M1011_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.835
cc_38 N_GND_c_38_p N_A_27_521#_M1011_g 0.00502587f $X=2.84 $Y=0.755 $X2=2.625
+ $Y2=0.835
cc_39 N_GND_c_4_p N_A_27_521#_M1011_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.625
+ $Y2=0.835
cc_40 N_GND_M1003_b N_A_27_521#_c_220_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.405
cc_41 N_GND_M1003_b N_A_27_521#_c_221_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.405
cc_42 N_GND_M1003_b N_A_27_521#_c_222_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.365
cc_43 N_GND_M1003_b N_A_27_521#_c_223_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.405
cc_44 N_GND_M1003_b N_A_27_521#_c_224_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.065
cc_45 N_GND_M1003_b N_A_27_521#_c_225_n 0.00710171f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.755
cc_46 N_GND_c_3_p N_A_27_521#_c_225_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.755
cc_47 N_GND_c_4_p N_A_27_521#_c_225_n 0.00475776f $X=2.38 $Y=0.19 $X2=0.69
+ $Y2=0.755
cc_48 N_GND_M1003_b N_A_27_521#_c_228_n 0.0190355f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_49 N_GND_c_11_p N_A_27_521#_c_228_n 0.00702738f $X=1.12 $Y=0.755 $X2=1.43
+ $Y2=1.455
cc_50 N_GND_M1003_b N_A_27_521#_c_230_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.455
cc_51 N_GND_M1003_b N_Y_c_334_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_52 N_GND_c_18_p N_Y_c_334_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_53 N_GND_c_24_p N_Y_c_334_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=0.755
cc_54 N_GND_c_4_p N_Y_c_334_n 0.0047139f $X=2.38 $Y=0.19 $X2=1.55 $Y2=0.755
cc_55 N_GND_M1003_b N_Y_c_338_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_56 N_GND_M1003_b N_Y_c_339_n 0.00154299f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.755
cc_57 N_GND_c_24_p N_Y_c_339_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=2.41 $Y2=0.755
cc_58 N_GND_c_32_p N_Y_c_339_n 0.00718527f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.755
cc_59 N_GND_c_4_p N_Y_c_339_n 0.0047139f $X=2.38 $Y=0.19 $X2=2.41 $Y2=0.755
cc_60 N_GND_M1003_b N_Y_c_343_n 0.0152877f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.11
cc_61 N_GND_M1003_b N_Y_c_344_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.115
cc_62 N_GND_c_11_p N_Y_c_344_n 0.00134236f $X=1.12 $Y=0.755 $X2=1.55 $Y2=1.115
cc_63 N_GND_c_18_p N_Y_c_344_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.55 $Y2=1.115
cc_64 N_GND_c_24_p N_Y_c_344_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=1.115
cc_65 N_GND_M1003_b N_Y_c_348_n 0.00463624f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.995
cc_66 N_GND_M1003_b Y 0.0305055f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.74
cc_67 N_GND_M1009_s N_Y_c_350_n 0.0100329f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1
cc_68 N_GND_c_18_p N_Y_c_350_n 0.0028844f $X=1.895 $Y=0.152 $X2=2.265 $Y2=1
cc_69 N_GND_c_24_p N_Y_c_350_n 0.0142303f $X=1.98 $Y=0.755 $X2=2.265 $Y2=1
cc_70 N_GND_c_32_p N_Y_c_350_n 0.0028844f $X=2.755 $Y=0.152 $X2=2.265 $Y2=1
cc_71 N_GND_M1003_b N_Y_c_354_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.11
cc_72 N_GND_M1003_b N_Y_c_355_n 0.00409378f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.115
cc_73 N_GND_c_24_p N_Y_c_355_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=2.41 $Y2=1.115
cc_74 N_GND_c_32_p N_Y_c_355_n 0.00245319f $X=2.755 $Y=0.152 $X2=2.41 $Y2=1.115
cc_75 N_GND_c_38_p N_Y_c_355_n 0.00134236f $X=2.84 $Y=0.755 $X2=2.41 $Y2=1.115
cc_76 N_GND_M1003_b N_Y_c_359_n 0.06145f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.995
cc_77 N_VDD_M1002_b N_B_M1002_g 0.0260091f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_78 N_VDD_c_78_p N_B_M1002_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.235
cc_79 N_VDD_c_79_p N_B_M1002_g 0.00468827f $X=2.38 $Y=4.25 $X2=0.475 $Y2=3.235
cc_80 N_VDD_M1002_b N_B_c_130_n 0.00375034f $X=-0.045 $Y=2.425 $X2=0.27
+ $Y2=2.195
cc_81 N_VDD_M1002_b B 0.0108395f $X=-0.045 $Y=2.425 $X2=0.27 $Y2=2.48
cc_82 N_VDD_M1002_b N_A_M1007_g 0.0195137f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_83 N_VDD_c_78_p N_A_M1007_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.235
cc_84 N_VDD_c_84_p N_A_M1007_g 0.00337744f $X=1.12 $Y=3.635 $X2=0.905 $Y2=3.235
cc_85 N_VDD_c_79_p N_A_M1007_g 0.00468827f $X=2.38 $Y=4.25 $X2=0.905 $Y2=3.235
cc_86 N_VDD_M1002_b N_A_c_158_n 0.00153494f $X=-0.045 $Y=2.425 $X2=0.95
+ $Y2=1.905
cc_87 N_VDD_M1007_d A 0.0077995f $X=0.98 $Y=2.605 $X2=0.95 $Y2=2.85
cc_88 N_VDD_c_84_p A 0.00247404f $X=1.12 $Y=3.635 $X2=0.95 $Y2=2.85
cc_89 N_VDD_M1002_b N_A_27_521#_c_231_n 0.0170965f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.48
cc_90 N_VDD_c_84_p N_A_27_521#_c_231_n 0.00337744f $X=1.12 $Y=3.635 $X2=1.335
+ $Y2=2.48
cc_91 N_VDD_c_91_p N_A_27_521#_c_231_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335
+ $Y2=2.48
cc_92 N_VDD_c_79_p N_A_27_521#_c_231_n 0.00468827f $X=2.38 $Y=4.25 $X2=1.335
+ $Y2=2.48
cc_93 N_VDD_M1002_b N_A_27_521#_c_201_n 0.00428234f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_94 N_VDD_M1002_b N_A_27_521#_c_236_n 0.017006f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.48
cc_95 N_VDD_c_84_p N_A_27_521#_c_236_n 3.67508e-19 $X=1.12 $Y=3.635 $X2=1.765
+ $Y2=2.48
cc_96 N_VDD_c_91_p N_A_27_521#_c_236_n 0.00610567f $X=1.895 $Y=4.287 $X2=1.765
+ $Y2=2.48
cc_97 N_VDD_c_97_p N_A_27_521#_c_236_n 0.0035715f $X=1.98 $Y=2.955 $X2=1.765
+ $Y2=2.48
cc_98 N_VDD_c_79_p N_A_27_521#_c_236_n 0.00470215f $X=2.38 $Y=4.25 $X2=1.765
+ $Y2=2.48
cc_99 N_VDD_M1002_b N_A_27_521#_c_209_n 0.00396043f $X=-0.045 $Y=2.425 $X2=2.12
+ $Y2=2.405
cc_100 N_VDD_c_97_p N_A_27_521#_c_209_n 0.00379272f $X=1.98 $Y=2.955 $X2=2.12
+ $Y2=2.405
cc_101 N_VDD_M1002_b N_A_27_521#_c_243_n 0.0166898f $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.48
cc_102 N_VDD_c_97_p N_A_27_521#_c_243_n 0.00337744f $X=1.98 $Y=2.955 $X2=2.195
+ $Y2=2.48
cc_103 N_VDD_c_103_p N_A_27_521#_c_243_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.195
+ $Y2=2.48
cc_104 N_VDD_c_79_p N_A_27_521#_c_243_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.195
+ $Y2=2.48
cc_105 N_VDD_M1002_b N_A_27_521#_c_215_n 0.00840215f $X=-0.045 $Y=2.425 $X2=2.55
+ $Y2=2.405
cc_106 N_VDD_M1002_b N_A_27_521#_c_248_n 0.0209036f $X=-0.045 $Y=2.425 $X2=2.625
+ $Y2=2.48
cc_107 N_VDD_c_103_p N_A_27_521#_c_248_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.625
+ $Y2=2.48
cc_108 N_VDD_c_108_p N_A_27_521#_c_248_n 0.00636672f $X=2.84 $Y=2.955 $X2=2.625
+ $Y2=2.48
cc_109 N_VDD_c_79_p N_A_27_521#_c_248_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.625
+ $Y2=2.48
cc_110 N_VDD_M1002_b N_A_27_521#_c_220_n 0.0021704f $X=-0.045 $Y=2.425 $X2=1.352
+ $Y2=2.405
cc_111 N_VDD_M1002_b N_A_27_521#_c_221_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=1.765 $Y2=2.405
cc_112 N_VDD_M1002_b N_A_27_521#_c_223_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=2.195 $Y2=2.405
cc_113 N_VDD_M1002_b N_A_27_521#_c_255_n 0.00156053f $X=-0.045 $Y=2.425 $X2=0.26
+ $Y2=3.295
cc_114 N_VDD_c_78_p N_A_27_521#_c_255_n 0.00736239f $X=1.035 $Y=4.287 $X2=0.26
+ $Y2=3.295
cc_115 N_VDD_c_79_p N_A_27_521#_c_255_n 0.00476261f $X=2.38 $Y=4.25 $X2=0.26
+ $Y2=3.295
cc_116 N_VDD_M1002_b N_A_27_521#_c_224_n 0.00106577f $X=-0.045 $Y=2.425 $X2=0.61
+ $Y2=3.065
cc_117 N_VDD_M1002_b N_Y_c_338_n 0.00367096f $X=-0.045 $Y=2.425 $X2=1.55
+ $Y2=2.11
cc_118 N_VDD_c_91_p N_Y_c_338_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.11
cc_119 N_VDD_c_79_p N_Y_c_338_n 0.00475776f $X=2.38 $Y=4.25 $X2=1.55 $Y2=2.11
cc_120 N_VDD_M1002_b N_Y_c_343_n 0.00380347f $X=-0.045 $Y=2.425 $X2=2.41
+ $Y2=2.11
cc_121 N_VDD_c_103_p N_Y_c_343_n 0.00734006f $X=2.755 $Y=4.287 $X2=2.41 $Y2=2.11
cc_122 N_VDD_c_79_p N_Y_c_343_n 0.00475776f $X=2.38 $Y=4.25 $X2=2.41 $Y2=2.11
cc_123 N_VDD_c_97_p N_Y_c_354_n 0.00634153f $X=1.98 $Y=2.955 $X2=2.265 $Y2=2.11
cc_124 N_B_M1003_g N_A_M1000_g 0.0358421f $X=0.475 $Y=0.835 $X2=0.905 $Y2=0.835
cc_125 N_B_c_129_n N_A_M1007_g 0.0819064f $X=0.475 $Y=2.195 $X2=0.905 $Y2=3.235
cc_126 N_B_M1003_g N_A_c_157_n 0.0148656f $X=0.475 $Y=0.835 $X2=0.95 $Y2=1.905
cc_127 N_B_M1003_g N_A_c_158_n 0.00121111f $X=0.475 $Y=0.835 $X2=0.95 $Y2=1.905
cc_128 N_B_M1002_g N_A_27_521#_c_259_n 0.0136492f $X=0.475 $Y=3.235 $X2=0.525
+ $Y2=3.15
cc_129 B N_A_27_521#_c_259_n 0.00520961f $X=0.27 $Y=2.48 $X2=0.525 $Y2=3.15
cc_130 N_B_c_130_n N_A_27_521#_c_261_n 0.00369517f $X=0.27 $Y=2.195 $X2=0.345
+ $Y2=3.15
cc_131 B N_A_27_521#_c_261_n 0.00431991f $X=0.27 $Y=2.48 $X2=0.345 $Y2=3.15
cc_132 N_B_M1003_g N_A_27_521#_c_224_n 0.0231435f $X=0.475 $Y=0.835 $X2=0.61
+ $Y2=3.065
cc_133 N_B_M1002_g N_A_27_521#_c_224_n 0.026563f $X=0.475 $Y=3.235 $X2=0.61
+ $Y2=3.065
cc_134 N_B_c_129_n N_A_27_521#_c_224_n 0.00764878f $X=0.475 $Y=2.195 $X2=0.61
+ $Y2=3.065
cc_135 N_B_c_130_n N_A_27_521#_c_224_n 0.0350086f $X=0.27 $Y=2.195 $X2=0.61
+ $Y2=3.065
cc_136 B N_A_27_521#_c_224_n 0.00758489f $X=0.27 $Y=2.48 $X2=0.61 $Y2=3.065
cc_137 N_B_M1003_g N_A_27_521#_c_225_n 0.00713391f $X=0.475 $Y=0.835 $X2=0.69
+ $Y2=0.755
cc_138 N_B_M1003_g N_A_27_521#_c_230_n 0.0113001f $X=0.475 $Y=0.835 $X2=0.65
+ $Y2=1.455
cc_139 N_A_M1000_g N_A_27_521#_M1001_g 0.0265272f $X=0.905 $Y=0.835 $X2=1.335
+ $Y2=0.835
cc_140 A N_A_27_521#_c_231_n 0.00374181f $X=0.95 $Y=2.85 $X2=1.335 $Y2=2.48
cc_141 N_A_M1007_g N_A_27_521#_c_200_n 0.00914307f $X=0.905 $Y=3.235 $X2=1.37
+ $Y2=2.33
cc_142 N_A_c_157_n N_A_27_521#_c_200_n 0.0204279f $X=0.95 $Y=1.905 $X2=1.37
+ $Y2=2.33
cc_143 N_A_c_158_n N_A_27_521#_c_200_n 0.00375034f $X=0.95 $Y=1.905 $X2=1.37
+ $Y2=2.33
cc_144 N_A_M1000_g N_A_27_521#_c_208_n 0.0119161f $X=0.905 $Y=0.835 $X2=1.84
+ $Y2=1.365
cc_145 N_A_M1007_g N_A_27_521#_c_220_n 0.0533175f $X=0.905 $Y=3.235 $X2=1.352
+ $Y2=2.405
cc_146 N_A_c_158_n N_A_27_521#_c_220_n 0.00358357f $X=0.95 $Y=1.905 $X2=1.352
+ $Y2=2.405
cc_147 N_A_M1007_g N_A_27_521#_c_259_n 0.00457566f $X=0.905 $Y=3.235 $X2=0.525
+ $Y2=3.15
cc_148 N_A_M1000_g N_A_27_521#_c_224_n 0.00429604f $X=0.905 $Y=0.835 $X2=0.61
+ $Y2=3.065
cc_149 N_A_M1007_g N_A_27_521#_c_224_n 0.00776428f $X=0.905 $Y=3.235 $X2=0.61
+ $Y2=3.065
cc_150 N_A_c_157_n N_A_27_521#_c_224_n 0.0021255f $X=0.95 $Y=1.905 $X2=0.61
+ $Y2=3.065
cc_151 N_A_c_158_n N_A_27_521#_c_224_n 0.0822139f $X=0.95 $Y=1.905 $X2=0.61
+ $Y2=3.065
cc_152 A N_A_27_521#_c_224_n 0.00866797f $X=0.95 $Y=2.85 $X2=0.61 $Y2=3.065
cc_153 N_A_M1000_g N_A_27_521#_c_225_n 0.00713391f $X=0.905 $Y=0.835 $X2=0.69
+ $Y2=0.755
cc_154 N_A_M1000_g N_A_27_521#_c_228_n 0.0163305f $X=0.905 $Y=0.835 $X2=1.43
+ $Y2=1.455
cc_155 N_A_c_157_n N_A_27_521#_c_228_n 0.00276813f $X=0.95 $Y=1.905 $X2=1.43
+ $Y2=1.455
cc_156 N_A_c_158_n N_A_27_521#_c_228_n 0.0114342f $X=0.95 $Y=1.905 $X2=1.43
+ $Y2=1.455
cc_157 A A_110_521# 0.0123256f $X=0.95 $Y=2.85 $X2=0.55 $Y2=2.605
cc_158 N_A_c_158_n N_Y_c_338_n 0.0206732f $X=0.95 $Y=1.905 $X2=1.55 $Y2=2.11
cc_159 A N_Y_c_338_n 0.00659455f $X=0.95 $Y=2.85 $X2=1.55 $Y2=2.11
cc_160 N_A_M1000_g N_Y_c_344_n 8.01483e-19 $X=0.905 $Y=0.835 $X2=1.55 $Y2=1.115
cc_161 N_A_c_157_n N_Y_c_348_n 3.73261e-19 $X=0.95 $Y=1.905 $X2=1.55 $Y2=1.995
cc_162 N_A_c_158_n N_Y_c_348_n 0.0059581f $X=0.95 $Y=1.905 $X2=1.55 $Y2=1.995
cc_163 N_A_M1000_g Y 6.73508e-19 $X=0.905 $Y=0.835 $X2=1.555 $Y2=1.74
cc_164 N_A_c_158_n Y 0.00825539f $X=0.95 $Y=1.905 $X2=1.555 $Y2=1.74
cc_165 N_A_27_521#_c_259_n A_110_521# 0.00613297f $X=0.525 $Y=3.15 $X2=0.55
+ $Y2=2.605
cc_166 N_A_27_521#_c_224_n A_110_521# 0.00377193f $X=0.61 $Y=3.065 $X2=0.55
+ $Y2=2.605
cc_167 N_A_27_521#_M1001_g N_Y_c_334_n 0.00182852f $X=1.335 $Y=0.835 $X2=1.55
+ $Y2=0.755
cc_168 N_A_27_521#_M1009_g N_Y_c_334_n 0.00182852f $X=1.765 $Y=0.835 $X2=1.55
+ $Y2=0.755
cc_169 N_A_27_521#_c_208_n N_Y_c_334_n 0.0016986f $X=1.84 $Y=1.365 $X2=1.55
+ $Y2=0.755
cc_170 N_A_27_521#_c_228_n N_Y_c_334_n 0.00498892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_171 N_A_27_521#_c_231_n N_Y_c_338_n 0.0020967f $X=1.335 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_172 N_A_27_521#_c_200_n N_Y_c_338_n 0.00744772f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_173 N_A_27_521#_c_201_n N_Y_c_338_n 0.0168228f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_174 N_A_27_521#_c_236_n N_Y_c_338_n 0.00375894f $X=1.765 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_175 N_A_27_521#_c_208_n N_Y_c_338_n 0.0013767f $X=1.84 $Y=1.365 $X2=1.55
+ $Y2=2.11
cc_176 N_A_27_521#_c_228_n N_Y_c_338_n 0.00273485f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_177 N_A_27_521#_M1010_g N_Y_c_339_n 0.00182852f $X=2.195 $Y=0.835 $X2=2.41
+ $Y2=0.755
cc_178 N_A_27_521#_c_214_n N_Y_c_339_n 0.00274041f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=0.755
cc_179 N_A_27_521#_M1011_g N_Y_c_339_n 0.00182852f $X=2.625 $Y=0.835 $X2=2.41
+ $Y2=0.755
cc_180 N_A_27_521#_c_243_n N_Y_c_343_n 0.00375894f $X=2.195 $Y=2.48 $X2=2.41
+ $Y2=2.11
cc_181 N_A_27_521#_c_214_n N_Y_c_343_n 0.00250559f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=2.11
cc_182 N_A_27_521#_c_215_n N_Y_c_343_n 0.0206674f $X=2.55 $Y=2.405 $X2=2.41
+ $Y2=2.11
cc_183 N_A_27_521#_c_248_n N_Y_c_343_n 0.00375894f $X=2.625 $Y=2.48 $X2=2.41
+ $Y2=2.11
cc_184 N_A_27_521#_M1001_g N_Y_c_344_n 0.00481614f $X=1.335 $Y=0.835 $X2=1.55
+ $Y2=1.115
cc_185 N_A_27_521#_M1009_g N_Y_c_344_n 0.00198614f $X=1.765 $Y=0.835 $X2=1.55
+ $Y2=1.115
cc_186 N_A_27_521#_c_228_n N_Y_c_344_n 0.00238892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1.115
cc_187 N_A_27_521#_c_200_n N_Y_c_348_n 0.00821104f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=1.995
cc_188 N_A_27_521#_c_201_n N_Y_c_348_n 0.00229755f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=1.995
cc_189 N_A_27_521#_c_208_n N_Y_c_348_n 0.00174847f $X=1.84 $Y=1.365 $X2=1.55
+ $Y2=1.995
cc_190 N_A_27_521#_c_228_n N_Y_c_348_n 0.00181779f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1.995
cc_191 N_A_27_521#_M1001_g Y 0.00251111f $X=1.335 $Y=0.835 $X2=1.555 $Y2=1.74
cc_192 N_A_27_521#_c_200_n Y 0.00892438f $X=1.37 $Y=2.33 $X2=1.555 $Y2=1.74
cc_193 N_A_27_521#_M1009_g Y 0.00251111f $X=1.765 $Y=0.835 $X2=1.555 $Y2=1.74
cc_194 N_A_27_521#_c_208_n Y 0.012793f $X=1.84 $Y=1.365 $X2=1.555 $Y2=1.74
cc_195 N_A_27_521#_c_228_n Y 0.0147088f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_196 N_A_27_521#_M1009_g N_Y_c_350_n 0.00873177f $X=1.765 $Y=0.835 $X2=2.265
+ $Y2=1
cc_197 N_A_27_521#_c_206_n N_Y_c_350_n 0.00213861f $X=2.12 $Y=1.365 $X2=2.265
+ $Y2=1
cc_198 N_A_27_521#_M1010_g N_Y_c_350_n 0.00873177f $X=2.195 $Y=0.835 $X2=2.265
+ $Y2=1
cc_199 N_A_27_521#_c_208_n N_Y_c_354_n 0.0121767f $X=1.84 $Y=1.365 $X2=2.265
+ $Y2=2.11
cc_200 N_A_27_521#_c_221_n N_Y_c_354_n 0.0158479f $X=1.765 $Y=2.405 $X2=2.265
+ $Y2=2.11
cc_201 N_A_27_521#_M1010_g N_Y_c_355_n 0.00198614f $X=2.195 $Y=0.835 $X2=2.41
+ $Y2=1.115
cc_202 N_A_27_521#_M1011_g N_Y_c_355_n 0.00878256f $X=2.625 $Y=0.835 $X2=2.41
+ $Y2=1.115
cc_203 N_A_27_521#_M1010_g N_Y_c_359_n 0.00251111f $X=2.195 $Y=0.835 $X2=2.41
+ $Y2=1.995
cc_204 N_A_27_521#_c_214_n N_Y_c_359_n 0.0184054f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=1.995
cc_205 N_A_27_521#_M1011_g N_Y_c_359_n 0.00251111f $X=2.625 $Y=0.835 $X2=2.41
+ $Y2=1.995
cc_206 N_A_27_521#_c_222_n N_Y_c_359_n 0.00140336f $X=2.195 $Y=1.365 $X2=2.41
+ $Y2=1.995
cc_207 N_A_27_521#_c_223_n N_Y_c_359_n 0.00372651f $X=2.195 $Y=2.405 $X2=2.41
+ $Y2=1.995
