magic
tech sky130A
magscale 1 2
timestamp 1612371069
<< nwell >>
rect -9 529 1435 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 252 115 282 243
rect 338 115 368 243
rect 410 115 440 243
rect 496 115 526 243
rect 582 115 612 243
rect 668 115 698 243
rect 754 115 784 243
rect 840 115 870 243
rect 922 115 952 243
rect 1004 115 1034 243
rect 1102 115 1132 225
rect 1292 115 1322 225
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
rect 338 565 368 965
rect 410 565 440 965
rect 496 565 526 965
rect 582 565 612 965
rect 668 565 698 965
rect 754 565 784 965
rect 840 565 870 965
rect 922 565 952 965
rect 1004 565 1034 965
rect 1102 713 1132 965
rect 1292 713 1322 965
<< ndiff >>
rect 27 228 80 243
rect 27 131 35 228
rect 69 131 80 228
rect 27 115 80 131
rect 110 165 166 243
rect 110 131 121 165
rect 155 131 166 165
rect 110 115 166 131
rect 196 228 252 243
rect 196 131 207 228
rect 241 131 252 228
rect 196 115 252 131
rect 282 228 338 243
rect 282 131 293 228
rect 327 131 338 228
rect 282 115 338 131
rect 368 115 410 243
rect 440 228 496 243
rect 440 131 451 228
rect 485 131 496 228
rect 440 115 496 131
rect 526 228 582 243
rect 526 131 537 228
rect 571 131 582 228
rect 526 115 582 131
rect 612 165 668 243
rect 612 131 623 165
rect 657 131 668 165
rect 612 115 668 131
rect 698 228 754 243
rect 698 131 709 228
rect 743 131 754 228
rect 698 115 754 131
rect 784 165 840 243
rect 784 131 795 165
rect 829 131 840 165
rect 784 115 840 131
rect 870 115 922 243
rect 952 115 1004 243
rect 1034 228 1087 243
rect 1034 131 1045 228
rect 1079 225 1087 228
rect 1079 131 1102 225
rect 1034 115 1102 131
rect 1132 165 1185 225
rect 1132 131 1143 165
rect 1177 131 1185 165
rect 1132 115 1185 131
rect 1239 165 1292 225
rect 1239 131 1247 165
rect 1281 131 1292 165
rect 1239 115 1292 131
rect 1322 165 1375 225
rect 1322 131 1333 165
rect 1367 131 1375 165
rect 1322 115 1375 131
<< pdiff >>
rect 27 949 80 965
rect 27 677 35 949
rect 69 677 80 949
rect 27 565 80 677
rect 110 949 166 965
rect 110 745 121 949
rect 155 745 166 949
rect 110 565 166 745
rect 196 949 252 965
rect 196 677 207 949
rect 241 677 252 949
rect 196 565 252 677
rect 282 949 338 965
rect 282 677 293 949
rect 327 677 338 949
rect 282 565 338 677
rect 368 565 410 965
rect 440 949 496 965
rect 440 677 451 949
rect 485 677 496 949
rect 440 565 496 677
rect 526 949 582 965
rect 526 677 537 949
rect 571 677 582 949
rect 526 565 582 677
rect 612 949 668 965
rect 612 745 623 949
rect 657 745 668 949
rect 612 565 668 745
rect 698 949 754 965
rect 698 677 709 949
rect 743 677 754 949
rect 698 565 754 677
rect 784 949 840 965
rect 784 677 795 949
rect 829 677 840 949
rect 784 565 840 677
rect 870 565 922 965
rect 952 565 1004 965
rect 1034 949 1102 965
rect 1034 745 1045 949
rect 1079 745 1102 949
rect 1034 713 1102 745
rect 1132 949 1185 965
rect 1132 813 1143 949
rect 1177 813 1185 949
rect 1132 713 1185 813
rect 1239 949 1292 965
rect 1239 813 1247 949
rect 1281 813 1292 949
rect 1239 713 1292 813
rect 1322 949 1375 965
rect 1322 813 1333 949
rect 1367 813 1375 949
rect 1322 713 1375 813
rect 1034 565 1087 713
<< ndiffc >>
rect 35 131 69 228
rect 121 131 155 165
rect 207 131 241 228
rect 293 131 327 228
rect 451 131 485 228
rect 537 131 571 228
rect 623 131 657 165
rect 709 131 743 228
rect 795 131 829 165
rect 1045 131 1079 228
rect 1143 131 1177 165
rect 1247 131 1281 165
rect 1333 131 1367 165
<< pdiffc >>
rect 35 677 69 949
rect 121 745 155 949
rect 207 677 241 949
rect 293 677 327 949
rect 451 677 485 949
rect 537 677 571 949
rect 623 745 657 949
rect 709 677 743 949
rect 795 677 829 949
rect 1045 745 1079 949
rect 1143 813 1177 949
rect 1247 813 1281 949
rect 1333 813 1367 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
rect 979 27 1003 61
rect 1037 27 1061 61
rect 1115 27 1139 61
rect 1173 27 1197 61
rect 1251 27 1275 61
rect 1309 27 1333 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
rect 299 1049 323 1083
rect 357 1049 381 1083
rect 435 1049 459 1083
rect 493 1049 517 1083
rect 571 1049 595 1083
rect 629 1049 653 1083
rect 707 1049 731 1083
rect 765 1049 789 1083
rect 843 1049 867 1083
rect 901 1049 925 1083
rect 979 1049 1003 1083
rect 1037 1049 1061 1083
rect 1115 1049 1139 1083
rect 1173 1049 1197 1083
rect 1251 1049 1275 1083
rect 1309 1049 1333 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
rect 1003 27 1037 61
rect 1139 27 1173 61
rect 1275 27 1309 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
rect 323 1049 357 1083
rect 459 1049 493 1083
rect 595 1049 629 1083
rect 731 1049 765 1083
rect 867 1049 901 1083
rect 1003 1049 1037 1083
rect 1139 1049 1173 1083
rect 1275 1049 1309 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 993
rect 338 965 368 993
rect 410 965 440 991
rect 496 965 526 991
rect 582 965 612 993
rect 668 965 698 993
rect 754 965 784 993
rect 840 965 870 993
rect 922 965 952 993
rect 1004 965 1034 993
rect 1102 965 1132 993
rect 1292 965 1322 993
rect 80 351 110 565
rect 166 533 196 565
rect 152 517 206 533
rect 152 483 162 517
rect 196 483 206 517
rect 152 467 206 483
rect 70 335 124 351
rect 70 301 80 335
rect 114 301 124 335
rect 70 285 124 301
rect 80 243 110 285
rect 166 243 196 467
rect 252 425 282 565
rect 338 467 368 565
rect 410 540 440 565
rect 496 540 526 565
rect 410 510 526 540
rect 338 451 430 467
rect 238 409 292 425
rect 238 375 248 409
rect 282 375 292 409
rect 238 359 292 375
rect 338 417 386 451
rect 420 417 430 451
rect 338 401 430 417
rect 252 243 282 359
rect 338 243 368 401
rect 472 351 502 510
rect 582 362 612 565
rect 668 499 698 565
rect 656 483 710 499
rect 656 449 666 483
rect 700 449 710 483
rect 656 433 710 449
rect 472 335 526 351
rect 472 315 482 335
rect 410 301 482 315
rect 516 301 526 335
rect 410 285 526 301
rect 568 346 622 362
rect 568 312 578 346
rect 612 312 622 346
rect 568 296 622 312
rect 410 243 440 285
rect 496 243 526 285
rect 582 243 612 296
rect 668 243 698 433
rect 754 351 784 565
rect 840 499 870 565
rect 826 483 880 499
rect 826 449 836 483
rect 870 449 880 483
rect 826 433 880 449
rect 922 461 952 565
rect 1004 533 1034 565
rect 1004 503 1048 533
rect 1102 532 1132 713
rect 922 445 976 461
rect 742 335 796 351
rect 742 301 752 335
rect 786 301 796 335
rect 742 285 796 301
rect 754 243 784 285
rect 840 243 870 433
rect 922 411 932 445
rect 966 411 976 445
rect 922 395 976 411
rect 922 243 952 395
rect 1018 351 1048 503
rect 1090 516 1144 532
rect 1292 529 1322 713
rect 1090 482 1100 516
rect 1134 482 1144 516
rect 1090 466 1144 482
rect 1255 513 1322 529
rect 1255 479 1265 513
rect 1299 479 1322 513
rect 1004 335 1058 351
rect 1004 301 1014 335
rect 1048 301 1058 335
rect 1004 285 1058 301
rect 1004 243 1034 285
rect 1102 225 1132 466
rect 1255 463 1322 479
rect 1292 225 1322 463
rect 80 81 110 115
rect 166 82 196 115
rect 252 82 282 115
rect 338 82 368 115
rect 410 82 440 115
rect 496 82 526 115
rect 582 82 612 115
rect 668 82 698 115
rect 754 82 784 115
rect 840 82 870 115
rect 922 82 952 115
rect 1004 82 1034 115
rect 1102 80 1132 115
rect 1292 80 1322 115
<< polycont >>
rect 162 483 196 517
rect 80 301 114 335
rect 248 375 282 409
rect 386 417 420 451
rect 666 449 700 483
rect 482 301 516 335
rect 578 312 612 346
rect 836 449 870 483
rect 752 301 786 335
rect 932 411 966 445
rect 1100 482 1134 516
rect 1265 479 1299 513
rect 1014 301 1048 335
<< locali >>
rect 0 1089 1408 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 323 1089
rect 357 1049 459 1089
rect 493 1049 595 1089
rect 629 1049 731 1089
rect 765 1049 867 1089
rect 901 1049 1003 1089
rect 1037 1049 1139 1089
rect 1173 1049 1275 1089
rect 1309 1049 1408 1089
rect 35 949 69 965
rect 121 949 155 1049
rect 121 729 155 745
rect 207 949 241 965
rect 35 657 69 677
rect 207 657 241 677
rect 35 623 241 657
rect 293 949 327 965
rect 293 590 327 677
rect 451 949 485 1049
rect 451 661 485 677
rect 537 949 571 965
rect 623 949 657 1049
rect 623 729 657 745
rect 709 949 743 965
rect 537 656 571 677
rect 709 656 743 677
rect 537 622 743 656
rect 795 949 829 965
rect 1045 949 1079 1049
rect 1045 729 1079 745
rect 1143 949 1177 965
rect 795 632 829 677
rect 1143 638 1177 813
rect 1247 949 1281 1049
rect 1247 797 1281 813
rect 1333 949 1367 965
rect 795 598 1100 632
rect 293 553 350 590
rect 795 589 829 598
rect 80 483 162 517
rect 196 483 212 517
rect 248 409 282 425
rect 248 359 282 375
rect 64 301 80 335
rect 114 301 130 335
rect 316 318 350 553
rect 752 554 829 589
rect 578 483 612 489
rect 386 451 444 483
rect 420 449 444 451
rect 650 449 666 483
rect 700 449 716 483
rect 386 401 420 417
rect 578 346 612 449
rect 666 409 700 449
rect 752 409 786 554
rect 1066 532 1100 598
rect 1177 604 1202 615
rect 1143 581 1202 604
rect 1066 516 1134 532
rect 1066 485 1100 516
rect 820 449 836 483
rect 870 449 886 483
rect 1089 482 1100 485
rect 1100 466 1134 482
rect 932 445 966 461
rect 932 409 966 411
rect 1168 409 1202 581
rect 1333 557 1367 813
rect 752 375 879 409
rect 1143 375 1202 409
rect 1265 513 1299 529
rect 293 284 350 318
rect 466 301 482 335
rect 516 301 532 335
rect 578 296 612 312
rect 736 301 752 335
rect 786 301 811 335
rect 293 261 327 284
rect 35 228 241 252
rect 69 218 207 228
rect 35 115 69 131
rect 121 165 155 181
rect 121 61 155 131
rect 207 114 241 131
rect 777 261 811 301
rect 293 114 327 131
rect 451 228 485 249
rect 451 61 485 131
rect 537 228 743 252
rect 571 218 709 228
rect 537 114 571 131
rect 623 165 657 181
rect 623 61 657 131
rect 845 181 879 375
rect 998 301 1014 335
rect 1048 301 1064 335
rect 709 114 743 131
rect 795 165 879 181
rect 829 131 879 165
rect 1045 228 1079 249
rect 795 114 829 131
rect 1045 61 1079 131
rect 1143 165 1177 375
rect 1265 261 1299 479
rect 1245 227 1299 261
rect 1143 115 1177 131
rect 1247 165 1281 181
rect 1247 61 1281 131
rect 1333 165 1367 523
rect 1333 115 1367 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 1003 61
rect 1037 21 1139 61
rect 1173 21 1275 61
rect 1309 21 1408 61
rect 0 0 1408 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 323 1083 357 1089
rect 323 1055 357 1083
rect 459 1083 493 1089
rect 459 1055 493 1083
rect 595 1083 629 1089
rect 595 1055 629 1083
rect 731 1083 765 1089
rect 731 1055 765 1083
rect 867 1083 901 1089
rect 867 1055 901 1083
rect 1003 1083 1037 1089
rect 1003 1055 1037 1083
rect 1139 1083 1173 1089
rect 1139 1055 1173 1083
rect 1275 1083 1309 1089
rect 1275 1055 1309 1083
rect 80 449 114 483
rect 248 375 282 409
rect 80 301 114 335
rect 444 449 478 483
rect 578 449 612 483
rect 666 375 700 409
rect 1143 604 1177 638
rect 836 449 870 483
rect 932 375 966 409
rect 482 301 516 335
rect 293 228 327 261
rect 293 227 327 228
rect 777 227 811 261
rect 1014 301 1048 335
rect 1211 227 1245 261
rect 1333 523 1367 557
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
rect 1003 27 1037 55
rect 1003 21 1037 27
rect 1139 27 1173 55
rect 1139 21 1173 27
rect 1275 27 1309 55
rect 1275 21 1309 27
<< metal1 >>
rect 0 1089 1408 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 323 1089
rect 357 1055 459 1089
rect 493 1055 595 1089
rect 629 1055 731 1089
rect 765 1055 867 1089
rect 901 1055 1003 1089
rect 1037 1055 1139 1089
rect 1173 1055 1275 1089
rect 1309 1055 1408 1089
rect 0 1049 1408 1055
rect 1131 638 1189 644
rect 1109 604 1143 638
rect 1177 604 1189 638
rect 1131 598 1189 604
rect 1321 557 1379 563
rect 1299 523 1333 557
rect 1367 523 1379 557
rect 1321 517 1379 523
rect 68 483 126 489
rect 432 483 490 489
rect 566 483 624 489
rect 824 483 882 489
rect 68 449 80 483
rect 114 449 444 483
rect 478 449 578 483
rect 612 450 836 483
rect 612 449 734 450
rect 812 449 836 450
rect 870 449 882 483
rect 68 443 126 449
rect 432 443 490 449
rect 566 443 624 449
rect 824 443 882 449
rect 236 409 294 415
rect 654 409 712 415
rect 920 409 978 415
rect 80 375 248 409
rect 282 375 666 409
rect 700 375 932 409
rect 966 375 978 409
rect 236 369 294 375
rect 654 369 712 375
rect 920 369 978 375
rect 68 335 126 341
rect 470 335 528 341
rect 1002 335 1060 341
rect 68 301 80 335
rect 114 301 482 335
rect 516 301 1014 335
rect 1048 301 1060 335
rect 68 295 126 301
rect 470 295 528 301
rect 1002 295 1060 301
rect 281 261 339 267
rect 765 261 823 267
rect 1199 261 1257 267
rect 281 227 293 261
rect 327 227 777 261
rect 811 227 1211 261
rect 1245 227 1257 261
rect 281 221 339 227
rect 765 221 823 227
rect 1199 221 1257 227
rect 0 55 1408 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 1003 55
rect 1037 21 1139 55
rect 1173 21 1275 55
rect 1309 21 1408 55
rect 0 0 1408 21
<< labels >>
rlabel viali 97 318 97 318 1 A
port 1 n
rlabel viali 265 392 265 392 1 CI
port 2 n
rlabel metal1 129 466 129 466 1 B
port 3 n
rlabel viali 1350 540 1350 540 1 CO
port 5 n
rlabel viali 1160 621 1160 621 1 S
port 6 n
rlabel viali 1228 244 1228 244 1 CON
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
