* File: sky130_osu_sc_18T_hs__aoi22_l.pxi.spice
* Created: Thu Oct 29 17:06:34 2020
* 
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%GND N_GND_M1005_s N_GND_M1007_d N_GND_M1005_b
+ N_GND_c_3_p N_GND_c_26_p N_GND_c_4_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_18T_HS__AOI22_L%GND
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%VDD N_VDD_M1004_d N_VDD_M1004_b N_VDD_c_46_p
+ N_VDD_c_47_p VDD N_VDD_c_48_p N_VDD_c_54_p
+ PM_SKY130_OSU_SC_18T_HS__AOI22_L%VDD
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%A0 N_A0_c_75_n N_A0_c_76_n N_A0_M1005_g
+ N_A0_M1004_g N_A0_c_80_n A0 N_A0_c_82_n N_A0_c_83_n
+ PM_SKY130_OSU_SC_18T_HS__AOI22_L%A0
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%A1 N_A1_M1003_g N_A1_c_113_n N_A1_M1000_g A1
+ N_A1_c_116_n PM_SKY130_OSU_SC_18T_HS__AOI22_L%A1
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%B0 N_B0_M1002_g N_B0_M1001_g N_B0_c_157_n
+ N_B0_c_158_n B0 N_B0_c_160_n PM_SKY130_OSU_SC_18T_HS__AOI22_L%B0
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%B1 N_B1_M1007_g N_B1_M1006_g B1 N_B1_c_203_n
+ N_B1_c_205_n PM_SKY130_OSU_SC_18T_HS__AOI22_L%B1
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%A_27_617# N_A_27_617#_M1004_s
+ N_A_27_617#_M1000_d N_A_27_617#_M1006_d N_A_27_617#_c_223_n
+ N_A_27_617#_c_226_n N_A_27_617#_c_239_n N_A_27_617#_c_228_n
+ N_A_27_617#_c_231_n PM_SKY130_OSU_SC_18T_HS__AOI22_L%A_27_617#
x_PM_SKY130_OSU_SC_18T_HS__AOI22_L%Y N_Y_M1003_d N_Y_M1001_d N_Y_c_284_n
+ N_Y_c_246_n N_Y_c_247_n Y N_Y_c_251_n N_Y_c_252_n N_Y_c_253_n
+ PM_SKY130_OSU_SC_18T_HS__AOI22_L%Y
cc_1 N_GND_M1005_b N_A0_c_75_n 0.0646163f $X=-0.045 $Y=0 $X2=0.295 $Y2=2.63
cc_2 N_GND_M1005_b N_A0_c_76_n 0.0198745f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.69
cc_3 N_GND_c_3_p N_A0_c_76_n 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.69
cc_4 N_GND_c_4_p N_A0_c_76_n 0.00606474f $X=1.825 $Y=0.152 $X2=0.475 $Y2=1.69
cc_5 N_GND_c_5_p N_A0_c_76_n 0.00468827f $X=1.7 $Y=0.17 $X2=0.475 $Y2=1.69
cc_6 N_GND_M1005_b N_A0_c_80_n 0.0324934f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.77
cc_7 N_GND_c_3_p N_A0_c_80_n 0.00534003f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.77
cc_8 N_GND_M1005_b N_A0_c_82_n 0.00438599f $X=-0.045 $Y=0 $X2=0.385 $Y2=2.765
cc_9 N_GND_M1005_b N_A0_c_83_n 0.0421132f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_10 N_GND_M1005_b N_A1_M1003_g 0.0384231f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_11 N_GND_c_4_p N_A1_M1003_g 0.00606474f $X=1.825 $Y=0.152 $X2=0.835 $Y2=1.075
cc_12 N_GND_c_5_p N_A1_M1003_g 0.00468827f $X=1.7 $Y=0.17 $X2=0.835 $Y2=1.075
cc_13 N_GND_M1005_b N_A1_c_113_n 0.0512047f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.57
cc_14 N_GND_M1005_b N_A1_M1000_g 0.0173082f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_15 N_GND_M1005_b A1 0.00204783f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.96
cc_16 N_GND_M1005_b N_A1_c_116_n 0.0119461f $X=-0.045 $Y=0 $X2=0.725 $Y2=2.255
cc_17 N_GND_M1005_b N_B0_M1002_g 0.0194676f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.075
cc_18 N_GND_c_4_p N_B0_M1002_g 0.00606474f $X=1.825 $Y=0.152 $X2=1.335 $Y2=1.075
cc_19 N_GND_c_5_p N_B0_M1002_g 0.00468827f $X=1.7 $Y=0.17 $X2=1.335 $Y2=1.075
cc_20 N_GND_M1005_b N_B0_M1001_g 0.0444247f $X=-0.045 $Y=0 $X2=1.335 $Y2=4.585
cc_21 N_GND_M1005_b N_B0_c_157_n 0.00417976f $X=-0.045 $Y=0 $X2=1.165 $Y2=1.9
cc_22 N_GND_M1005_b N_B0_c_158_n 0.0272094f $X=-0.045 $Y=0 $X2=1.255 $Y2=1.9
cc_23 N_GND_M1005_b B0 0.014652f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.59
cc_24 N_GND_M1005_b N_B0_c_160_n 0.0123234f $X=-0.045 $Y=0 $X2=1.165 $Y2=2.59
cc_25 N_GND_M1005_b N_B1_M1007_g 0.0434394f $X=-0.045 $Y=0 $X2=1.695 $Y2=1.075
cc_26 N_GND_c_26_p N_B1_M1007_g 0.00713292f $X=1.91 $Y=0.825 $X2=1.695 $Y2=1.075
cc_27 N_GND_c_4_p N_B1_M1007_g 0.00606474f $X=1.825 $Y=0.152 $X2=1.695 $Y2=1.075
cc_28 N_GND_c_5_p N_B1_M1007_g 0.00468827f $X=1.7 $Y=0.17 $X2=1.695 $Y2=1.075
cc_29 N_GND_M1005_b N_B1_M1006_g 0.0420537f $X=-0.045 $Y=0 $X2=1.765 $Y2=4.585
cc_30 N_GND_M1005_b B1 0.0102806f $X=-0.045 $Y=0 $X2=1.935 $Y2=2.225
cc_31 N_GND_M1005_b N_B1_c_203_n 0.00958758f $X=-0.045 $Y=0 $X2=1.935 $Y2=2.225
cc_32 N_GND_c_26_p N_B1_c_203_n 0.00412675f $X=1.91 $Y=0.825 $X2=1.935 $Y2=2.225
cc_33 N_GND_M1005_b N_B1_c_205_n 0.0577952f $X=-0.045 $Y=0 $X2=1.765 $Y2=2.205
cc_34 N_GND_c_26_p N_B1_c_205_n 0.00159273f $X=1.91 $Y=0.825 $X2=1.765 $Y2=2.205
cc_35 N_GND_c_26_p N_Y_c_246_n 7.45493e-19 $X=1.91 $Y=0.825 $X2=1.52 $Y2=1.48
cc_36 N_GND_M1005_b N_Y_c_247_n 0.00670877f $X=-0.045 $Y=0 $X2=1.23 $Y2=1.48
cc_37 N_GND_c_3_p N_Y_c_247_n 0.00115996f $X=0.26 $Y=0.825 $X2=1.23 $Y2=1.48
cc_38 N_GND_c_26_p N_Y_c_247_n 6.58722e-19 $X=1.91 $Y=0.825 $X2=1.23 $Y2=1.48
cc_39 N_GND_M1005_b Y 0.00206172f $X=-0.045 $Y=0 $X2=1.605 $Y2=1.7
cc_40 N_GND_M1005_b N_Y_c_251_n 0.00421975f $X=-0.045 $Y=0 $X2=1.595 $Y2=1.85
cc_41 N_GND_M1005_b N_Y_c_252_n 0.0173806f $X=-0.045 $Y=0 $X2=1.595 $Y2=1.85
cc_42 N_GND_M1005_b N_Y_c_253_n 0.00156987f $X=-0.045 $Y=0 $X2=1.085 $Y2=0.825
cc_43 N_GND_c_4_p N_Y_c_253_n 0.00738471f $X=1.825 $Y=0.152 $X2=1.085 $Y2=0.825
cc_44 N_GND_c_5_p N_Y_c_253_n 0.00476747f $X=1.7 $Y=0.17 $X2=1.085 $Y2=0.825
cc_45 N_VDD_M1004_b N_A0_M1004_g 0.0258897f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_46 N_VDD_c_46_p N_A0_M1004_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.475 $Y2=4.585
cc_47 N_VDD_c_47_p N_A0_M1004_g 0.00606474f $X=0.605 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_48 N_VDD_c_48_p N_A0_M1004_g 0.00468827f $X=1.7 $Y=6.49 $X2=0.475 $Y2=4.585
cc_49 N_VDD_M1004_d A0 0.00612249f $X=0.55 $Y=3.085 $X2=0.385 $Y2=3.33
cc_50 N_VDD_M1004_b N_A0_c_82_n 0.00618364f $X=-0.045 $Y=2.905 $X2=0.385
+ $Y2=2.765
cc_51 N_VDD_M1004_b N_A1_M1000_g 0.0189807f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_52 N_VDD_c_46_p N_A1_M1000_g 0.00354579f $X=0.69 $Y=4.475 $X2=0.905 $Y2=4.585
cc_53 N_VDD_c_48_p N_A1_M1000_g 0.00468827f $X=1.7 $Y=6.49 $X2=0.905 $Y2=4.585
cc_54 N_VDD_c_54_p N_A1_M1000_g 0.00606474f $X=1.7 $Y=6.44 $X2=0.905 $Y2=4.585
cc_55 N_VDD_M1004_b A1 0.0104103f $X=-0.045 $Y=2.905 $X2=0.725 $Y2=2.96
cc_56 N_VDD_M1004_b N_A1_c_116_n 0.00527425f $X=-0.045 $Y=2.905 $X2=0.725
+ $Y2=2.255
cc_57 N_VDD_M1004_b N_B0_M1001_g 0.0205564f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=4.585
cc_58 N_VDD_c_48_p N_B0_M1001_g 0.00468827f $X=1.7 $Y=6.49 $X2=1.335 $Y2=4.585
cc_59 N_VDD_c_54_p N_B0_M1001_g 0.0042036f $X=1.7 $Y=6.44 $X2=1.335 $Y2=4.585
cc_60 N_VDD_M1004_b N_B1_M1006_g 0.029191f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=4.585
cc_61 N_VDD_c_48_p N_B1_M1006_g 0.00468827f $X=1.7 $Y=6.49 $X2=1.765 $Y2=4.585
cc_62 N_VDD_c_54_p N_B1_M1006_g 0.0042036f $X=1.7 $Y=6.44 $X2=1.765 $Y2=4.585
cc_63 N_VDD_M1004_b N_A_27_617#_c_223_n 0.00156053f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=4.135
cc_64 N_VDD_c_47_p N_A_27_617#_c_223_n 0.00736239f $X=0.605 $Y=6.507 $X2=0.26
+ $Y2=4.135
cc_65 N_VDD_c_48_p N_A_27_617#_c_223_n 0.00476261f $X=1.7 $Y=6.49 $X2=0.26
+ $Y2=4.135
cc_66 N_VDD_M1004_d N_A_27_617#_c_226_n 0.00743028f $X=0.55 $Y=3.085 $X2=1.035
+ $Y2=3.97
cc_67 N_VDD_c_46_p N_A_27_617#_c_226_n 0.0135055f $X=0.69 $Y=4.475 $X2=1.035
+ $Y2=3.97
cc_68 N_VDD_M1004_b N_A_27_617#_c_228_n 0.00156987f $X=-0.045 $Y=2.905 $X2=1.895
+ $Y2=6
cc_69 N_VDD_c_48_p N_A_27_617#_c_228_n 0.0233834f $X=1.7 $Y=6.49 $X2=1.895 $Y2=6
cc_70 N_VDD_c_54_p N_A_27_617#_c_228_n 0.030762f $X=1.7 $Y=6.44 $X2=1.895 $Y2=6
cc_71 N_VDD_M1004_b N_A_27_617#_c_231_n 0.00155118f $X=-0.045 $Y=2.905 $X2=1.205
+ $Y2=6
cc_72 N_VDD_c_48_p N_A_27_617#_c_231_n 0.0048048f $X=1.7 $Y=6.49 $X2=1.205 $Y2=6
cc_73 N_VDD_c_54_p N_A_27_617#_c_231_n 0.00738333f $X=1.7 $Y=6.44 $X2=1.205
+ $Y2=6
cc_74 N_VDD_M1004_b N_Y_c_252_n 0.00371086f $X=-0.045 $Y=2.905 $X2=1.595
+ $Y2=1.85
cc_75 N_A0_c_75_n N_A1_M1003_g 0.00899556f $X=0.295 $Y=2.63 $X2=0.835 $Y2=1.075
cc_76 N_A0_c_76_n N_A1_M1003_g 0.0857013f $X=0.475 $Y=1.69 $X2=0.835 $Y2=1.075
cc_77 N_A0_c_75_n N_A1_c_113_n 0.0253071f $X=0.295 $Y=2.63 $X2=0.905 $Y2=2.57
cc_78 N_A0_c_75_n N_A1_M1000_g 0.00107789f $X=0.295 $Y=2.63 $X2=0.905 $Y2=4.585
cc_79 A0 N_A1_M1000_g 0.00309207f $X=0.385 $Y=3.33 $X2=0.905 $Y2=4.585
cc_80 N_A0_c_82_n N_A1_M1000_g 0.00277246f $X=0.385 $Y=2.765 $X2=0.905 $Y2=4.585
cc_81 N_A0_c_83_n N_A1_M1000_g 0.0804191f $X=0.475 $Y=2.765 $X2=0.905 $Y2=4.585
cc_82 A0 A1 0.00560453f $X=0.385 $Y=3.33 $X2=0.725 $Y2=2.96
cc_83 N_A0_c_82_n A1 0.00775911f $X=0.385 $Y=2.765 $X2=0.725 $Y2=2.96
cc_84 N_A0_c_83_n A1 0.00417236f $X=0.475 $Y=2.765 $X2=0.725 $Y2=2.96
cc_85 N_A0_c_75_n N_A1_c_116_n 0.00549523f $X=0.295 $Y=2.63 $X2=0.725 $Y2=2.255
cc_86 N_A0_c_82_n N_A1_c_116_n 0.0297299f $X=0.385 $Y=2.765 $X2=0.725 $Y2=2.255
cc_87 N_A0_c_83_n N_A1_c_116_n 0.00281397f $X=0.475 $Y=2.765 $X2=0.725 $Y2=2.255
cc_88 A0 N_A_27_617#_M1004_s 0.0124771f $X=0.385 $Y=3.33 $X2=0.135 $Y2=3.085
cc_89 N_A0_c_82_n N_A_27_617#_M1004_s 0.00882571f $X=0.385 $Y=2.765 $X2=0.135
+ $Y2=3.085
cc_90 N_A0_M1004_g N_A_27_617#_c_226_n 0.0152354f $X=0.475 $Y=4.585 $X2=1.035
+ $Y2=3.97
cc_91 A0 N_A_27_617#_c_226_n 0.00806826f $X=0.385 $Y=3.33 $X2=1.035 $Y2=3.97
cc_92 N_A0_c_82_n N_A_27_617#_c_226_n 0.00155918f $X=0.385 $Y=2.765 $X2=1.035
+ $Y2=3.97
cc_93 A0 N_A_27_617#_c_239_n 0.00366477f $X=0.385 $Y=3.33 $X2=0.345 $Y2=3.97
cc_94 N_A0_c_82_n N_A_27_617#_c_239_n 0.00100283f $X=0.385 $Y=2.765 $X2=0.345
+ $Y2=3.97
cc_95 N_A1_M1003_g N_B0_M1002_g 0.0197201f $X=0.835 $Y=1.075 $X2=1.335 $Y2=1.075
cc_96 N_A1_M1003_g N_B0_M1001_g 0.00961043f $X=0.835 $Y=1.075 $X2=1.335
+ $Y2=4.585
cc_97 N_A1_c_113_n N_B0_M1001_g 0.0772733f $X=0.905 $Y=2.57 $X2=1.335 $Y2=4.585
cc_98 A1 N_B0_M1001_g 0.0011808f $X=0.725 $Y=2.96 $X2=1.335 $Y2=4.585
cc_99 N_A1_M1003_g N_B0_c_157_n 0.00591675f $X=0.835 $Y=1.075 $X2=1.165 $Y2=1.9
cc_100 N_A1_M1003_g N_B0_c_158_n 0.0198874f $X=0.835 $Y=1.075 $X2=1.255 $Y2=1.9
cc_101 N_A1_c_113_n B0 0.0041793f $X=0.905 $Y=2.57 $X2=1.165 $Y2=2.59
cc_102 N_A1_M1000_g B0 0.00301191f $X=0.905 $Y=4.585 $X2=1.165 $Y2=2.59
cc_103 A1 B0 0.00582284f $X=0.725 $Y=2.96 $X2=1.165 $Y2=2.59
cc_104 N_A1_c_116_n B0 0.0073589f $X=0.725 $Y=2.255 $X2=1.165 $Y2=2.59
cc_105 N_A1_M1003_g N_B0_c_160_n 0.0032219f $X=0.835 $Y=1.075 $X2=1.165 $Y2=2.59
cc_106 N_A1_c_113_n N_B0_c_160_n 0.0017522f $X=0.905 $Y=2.57 $X2=1.165 $Y2=2.59
cc_107 N_A1_c_116_n N_B0_c_160_n 0.0272019f $X=0.725 $Y=2.255 $X2=1.165 $Y2=2.59
cc_108 N_A1_M1000_g N_A_27_617#_c_226_n 0.0180368f $X=0.905 $Y=4.585 $X2=1.035
+ $Y2=3.97
cc_109 N_A1_M1003_g N_Y_c_247_n 0.0047962f $X=0.835 $Y=1.075 $X2=1.23 $Y2=1.48
cc_110 A1 N_Y_c_252_n 0.00544969f $X=0.725 $Y=2.96 $X2=1.595 $Y2=1.85
cc_111 N_A1_M1003_g N_Y_c_253_n 0.0103431f $X=0.835 $Y=1.075 $X2=1.085 $Y2=0.825
cc_112 N_B0_M1002_g N_B1_M1007_g 0.0527984f $X=1.335 $Y=1.075 $X2=1.695
+ $Y2=1.075
cc_113 N_B0_c_157_n N_B1_M1007_g 4.28971e-19 $X=1.165 $Y=1.9 $X2=1.695 $Y2=1.075
cc_114 N_B0_M1001_g N_B1_c_205_n 0.0866545f $X=1.335 $Y=4.585 $X2=1.765
+ $Y2=2.205
cc_115 N_B0_c_158_n N_B1_c_205_n 0.0527984f $X=1.255 $Y=1.9 $X2=1.765 $Y2=2.205
cc_116 N_B0_M1001_g N_A_27_617#_c_228_n 0.0130261f $X=1.335 $Y=4.585 $X2=1.895
+ $Y2=6
cc_117 N_B0_M1002_g N_Y_c_246_n 0.0126098f $X=1.335 $Y=1.075 $X2=1.52 $Y2=1.48
cc_118 N_B0_c_157_n N_Y_c_246_n 0.00477495f $X=1.165 $Y=1.9 $X2=1.52 $Y2=1.48
cc_119 N_B0_M1002_g N_Y_c_247_n 7.17871e-19 $X=1.335 $Y=1.075 $X2=1.23 $Y2=1.48
cc_120 N_B0_c_157_n N_Y_c_247_n 0.00568984f $X=1.165 $Y=1.9 $X2=1.23 $Y2=1.48
cc_121 N_B0_c_158_n N_Y_c_247_n 0.00131678f $X=1.255 $Y=1.9 $X2=1.23 $Y2=1.48
cc_122 N_B0_M1002_g Y 0.0019765f $X=1.335 $Y=1.075 $X2=1.605 $Y2=1.7
cc_123 N_B0_c_157_n N_Y_c_251_n 0.00751098f $X=1.165 $Y=1.9 $X2=1.595 $Y2=1.85
cc_124 N_B0_c_158_n N_Y_c_251_n 0.00382225f $X=1.255 $Y=1.9 $X2=1.595 $Y2=1.85
cc_125 N_B0_c_157_n N_Y_c_252_n 0.0201907f $X=1.165 $Y=1.9 $X2=1.595 $Y2=1.85
cc_126 N_B0_c_158_n N_Y_c_252_n 0.0171279f $X=1.255 $Y=1.9 $X2=1.595 $Y2=1.85
cc_127 B0 N_Y_c_252_n 0.00659034f $X=1.165 $Y=2.59 $X2=1.595 $Y2=1.85
cc_128 N_B0_c_160_n N_Y_c_252_n 0.0300971f $X=1.165 $Y=2.59 $X2=1.595 $Y2=1.85
cc_129 N_B0_M1002_g N_Y_c_253_n 0.010214f $X=1.335 $Y=1.075 $X2=1.085 $Y2=0.825
cc_130 N_B0_c_157_n N_Y_c_253_n 0.00420445f $X=1.165 $Y=1.9 $X2=1.085 $Y2=0.825
cc_131 N_B0_c_158_n N_Y_c_253_n 0.00113527f $X=1.255 $Y=1.9 $X2=1.085 $Y2=0.825
cc_132 N_B1_M1006_g N_A_27_617#_c_228_n 0.0135543f $X=1.765 $Y=4.585 $X2=1.895
+ $Y2=6
cc_133 N_B1_M1007_g N_Y_c_246_n 0.0107689f $X=1.695 $Y=1.075 $X2=1.52 $Y2=1.48
cc_134 N_B1_M1007_g Y 0.00642782f $X=1.695 $Y=1.075 $X2=1.605 $Y2=1.7
cc_135 N_B1_M1007_g N_Y_c_251_n 0.0113776f $X=1.695 $Y=1.075 $X2=1.595 $Y2=1.85
cc_136 B1 N_Y_c_251_n 0.00545275f $X=1.935 $Y=2.225 $X2=1.595 $Y2=1.85
cc_137 N_B1_M1007_g N_Y_c_252_n 0.0097422f $X=1.695 $Y=1.075 $X2=1.595 $Y2=1.85
cc_138 B1 N_Y_c_252_n 0.00769441f $X=1.935 $Y=2.225 $X2=1.595 $Y2=1.85
cc_139 N_B1_c_203_n N_Y_c_252_n 0.0209874f $X=1.935 $Y=2.225 $X2=1.595 $Y2=1.85
cc_140 N_B1_c_205_n N_Y_c_252_n 0.0264693f $X=1.765 $Y=2.205 $X2=1.595 $Y2=1.85
cc_141 N_A_27_617#_c_228_n N_Y_M1001_d 0.00376923f $X=1.895 $Y=6 $X2=1.41
+ $Y2=3.085
cc_142 N_A_27_617#_c_228_n N_Y_c_284_n 0.0131604f $X=1.895 $Y=6 $X2=1.55
+ $Y2=4.135
cc_143 N_Y_c_246_n A_282_115# 0.0104934f $X=1.52 $Y=1.48 $X2=1.41 $Y2=0.575
