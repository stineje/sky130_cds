* File: sky130_osu_sc_12T_hs__dffr_1.pex.spice
* Created: Fri Nov 12 15:09:13 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%GND 1 2 3 4 5 6 7 8 9 121 125 127 134
+ 136 143 145 152 154 164 166 176 178 185 187 194 196 203 230 232
c249 194 0 6.51688e-20 $X=7.9 $Y=0.74
c250 176 0 1.71621e-19 $X=6.09 $Y=0.755
c251 152 0 3.07651e-19 $X=2.59 $Y=0.755
c252 134 0 6.24044e-20 $X=1.21 $Y=0.74
c253 121 0 2.41708e-19 $X=-0.05 $Y=0
r254 230 232 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.175 $Y2=0.152
r255 205 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.152
+ $X2=8.85 $Y2=0.152
r256 201 226 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.152
r257 201 203 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.74
r258 196 226 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.152
+ $X2=8.85 $Y2=0.152
r259 192 194 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.74
r260 188 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.152
+ $X2=7.04 $Y2=0.152
r261 183 222 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.152
r262 183 185 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.74
r263 179 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.152
+ $X2=6.09 $Y2=0.152
r264 178 222 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.152
+ $X2=7.04 $Y2=0.152
r265 174 221 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.152
r266 174 176 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.755
r267 166 221 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.152
+ $X2=6.09 $Y2=0.152
r268 162 164 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.34 $Y=0.305
+ $X2=4.34 $Y2=0.74
r269 155 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.152
+ $X2=2.59 $Y2=0.152
r270 150 217 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.152
r271 150 152 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.755
r272 146 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.152
+ $X2=2.07 $Y2=0.152
r273 145 217 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.152
+ $X2=2.59 $Y2=0.152
r274 141 216 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.152
r275 141 143 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.74
r276 137 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.152
+ $X2=1.21 $Y2=0.152
r277 136 216 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.152
+ $X2=2.07 $Y2=0.152
r278 132 215 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.152
r279 132 134 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.74
r280 127 215 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.152
+ $X2=1.21 $Y2=0.152
r281 123 125 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.755
r282 121 232 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=0.19 $X2=9.175 $Y2=0.19
r283 121 230 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=0.19 $X2=0.335 $Y2=0.19
r284 121 192 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r285 121 187 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r286 121 197 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.985 $Y2=0.152
r287 121 162 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.34 $Y2=0.305
r288 121 154 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.255 $Y2=0.152
r289 121 167 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.425 $Y2=0.152
r290 121 123 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r291 121 128 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r292 121 205 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.935 $Y2=0.152
r293 121 196 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.765 $Y2=0.152
r294 121 197 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=7.985 $Y2=0.152
r295 121 187 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r296 121 188 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.125 $Y2=0.152
r297 121 178 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.955 $Y2=0.152
r298 121 179 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.175 $Y2=0.152
r299 121 166 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.005 $Y2=0.152
r300 121 167 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.425 $Y2=0.152
r301 121 154 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=4.255 $Y2=0.152
r302 121 155 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=2.675 $Y2=0.152
r303 121 145 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.505 $Y2=0.152
r304 121 146 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.155 $Y2=0.152
r305 121 136 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.985 $Y2=0.152
r306 121 137 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.295 $Y2=0.152
r307 121 127 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.125 $Y2=0.152
r308 121 128 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r309 9 203 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.575 $X2=8.85 $Y2=0.74
r310 8 194 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.74
r311 7 185 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.575 $X2=7.04 $Y2=0.74
r312 6 176 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.575 $X2=6.09 $Y2=0.755
r313 5 164 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.575 $X2=4.34 $Y2=0.74
r314 4 152 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.575 $X2=2.59 $Y2=0.755
r315 3 143 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.74
r316 2 134 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.74
r317 1 125 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%VDD 1 2 3 4 5 6 7 85 89 91 99 107 109
+ 117 119 127 129 137 139 145 149 164 168
c124 145 0 1.98165e-19 $X=8.85 $Y=3.265
r125 164 168 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=4.287
+ $X2=9.175 $Y2=4.287
r126 153 164 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=4.25 $X2=0.335 $Y2=4.25
r127 149 168 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=4.25 $X2=9.175 $Y2=4.25
r128 147 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=4.287
+ $X2=8.85 $Y2=4.287
r129 147 149 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=8.935 $Y=4.287
+ $X2=9.175 $Y2=4.287
r130 143 162 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.85 $Y=4.135
+ $X2=8.85 $Y2=4.287
r131 143 145 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.85 $Y=4.135
+ $X2=8.85 $Y2=3.265
r132 140 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=4.287
+ $X2=7.83 $Y2=4.287
r133 140 142 21.9153 $w=3.03e-07 $l=5.8e-07 $layer=LI1_cond $X=7.915 $Y=4.287
+ $X2=8.495 $Y2=4.287
r134 139 162 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=4.287
+ $X2=8.85 $Y2=4.287
r135 139 142 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.765 $Y=4.287
+ $X2=8.495 $Y2=4.287
r136 135 161 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.83 $Y=4.135
+ $X2=7.83 $Y2=4.287
r137 135 137 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=7.83 $Y=4.135
+ $X2=7.83 $Y2=3.275
r138 132 134 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.455 $Y=4.287
+ $X2=7.135 $Y2=4.287
r139 130 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.09 $Y2=4.287
r140 130 132 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=4.287
+ $X2=6.455 $Y2=4.287
r141 129 161 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=4.287
+ $X2=7.83 $Y2=4.287
r142 129 134 23.0489 $w=3.03e-07 $l=6.1e-07 $layer=LI1_cond $X=7.745 $Y=4.287
+ $X2=7.135 $Y2=4.287
r143 125 159 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=4.287
r144 125 127 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.09 $Y=4.135
+ $X2=6.09 $Y2=3.21
r145 122 124 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=4.287
+ $X2=5.775 $Y2=4.287
r146 120 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=4.287
+ $X2=4.34 $Y2=4.287
r147 120 122 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.425 $Y=4.287
+ $X2=5.095 $Y2=4.287
r148 119 159 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=6.09 $Y2=4.287
r149 119 124 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=4.287
+ $X2=5.775 $Y2=4.287
r150 115 158 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.34 $Y=4.135
+ $X2=4.34 $Y2=4.287
r151 115 117 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.34 $Y=4.135
+ $X2=4.34 $Y2=3.295
r152 112 114 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=4.287
+ $X2=3.735 $Y2=4.287
r153 110 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=4.287
+ $X2=2.59 $Y2=4.287
r154 110 112 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.675 $Y=4.287
+ $X2=3.055 $Y2=4.287
r155 109 158 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=4.287
+ $X2=4.34 $Y2=4.287
r156 109 114 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=4.255 $Y=4.287
+ $X2=3.735 $Y2=4.287
r157 105 156 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.59 $Y=4.135
+ $X2=2.59 $Y2=4.287
r158 105 107 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.59 $Y=4.135
+ $X2=2.59 $Y2=3.295
r159 102 155 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=4.287
+ $X2=2 $Y2=4.287
r160 102 104 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=2.085 $Y=4.287
+ $X2=2.375 $Y2=4.287
r161 101 156 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=4.287
+ $X2=2.59 $Y2=4.287
r162 101 104 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=4.287
+ $X2=2.375 $Y2=4.287
r163 97 155 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2 $Y=4.135 $X2=2
+ $Y2=4.287
r164 97 99 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2 $Y=4.135 $X2=2
+ $Y2=3.275
r165 94 96 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=4.287
+ $X2=1.695 $Y2=4.287
r166 92 153 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=0.172 $Y2=4.287
r167 92 94 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=4.287
+ $X2=1.015 $Y2=4.287
r168 91 155 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=4.287
+ $X2=2 $Y2=4.287
r169 91 96 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.915 $Y=4.287
+ $X2=1.695 $Y2=4.287
r170 87 153 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.172 $Y2=4.287
r171 87 89 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=3.635
r172 85 149 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=4.135 $X2=9.175 $Y2=4.22
r173 85 142 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=4.135 $X2=8.495 $Y2=4.22
r174 85 161 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=4.135 $X2=7.815 $Y2=4.22
r175 85 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=4.135 $X2=7.135 $Y2=4.22
r176 85 132 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=4.135 $X2=6.455 $Y2=4.22
r177 85 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=4.135 $X2=5.775 $Y2=4.22
r178 85 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=4.135 $X2=5.095 $Y2=4.22
r179 85 158 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=4.135 $X2=4.415 $Y2=4.22
r180 85 114 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=4.135 $X2=3.735 $Y2=4.22
r181 85 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=4.135 $X2=3.055 $Y2=4.22
r182 85 104 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=4.135 $X2=2.375 $Y2=4.22
r183 85 96 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=4.135 $X2=1.695 $Y2=4.22
r184 85 94 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=4.135 $X2=1.015 $Y2=4.22
r185 85 153 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=4.135 $X2=0.335 $Y2=4.22
r186 7 145 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=2.605 $X2=8.85 $Y2=3.265
r187 6 137 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=3.025 $X2=7.83 $Y2=3.275
r188 5 127 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=5.95
+ $Y=2.605 $X2=6.09 $Y2=3.21
r189 4 117 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=2.605 $X2=4.34 $Y2=3.295
r190 3 107 300 $w=1.7e-07 $l=7.499e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.605 $X2=2.59 $Y2=3.295
r191 2 99 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=3.025 $X2=2 $Y2=3.275
r192 1 89 600 $w=1.7e-07 $l=1.09071e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.605 $X2=0.26 $Y2=3.635
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%RN 3 5 7 13 15 21
c38 21 0 7.50258e-20 $X=0.325 $Y=2.85
r39 19 21 0.00301932 $w=2.07e-07 $l=5e-09 $layer=MET1_cond $X=0.32 $Y=2.85
+ $X2=0.325 $Y2=2.85
r40 15 17 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.53 $Y2=1.825
r41 13 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=2.85
+ $X2=0.32 $Y2=2.85
r42 11 15 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=1.99
+ $X2=0.32 $Y2=1.825
r43 11 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=1.99 $X2=0.32
+ $Y2=2.85
r44 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.825 $X2=0.53 $Y2=1.825
r45 5 10 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.53 $Y2=1.825
r46 5 7 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=1.99
+ $X2=0.475 $Y2=3.235
r47 1 10 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.53 $Y2=1.825
r48 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.475 $Y=1.655
+ $X2=0.475 $Y2=0.85
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%A_110_115# 1 3 9 11 14 16 18 20 22 26 32
+ 36 41 42 43 46 51 55 59 60 61 63 65 68
c200 68 0 6.51688e-20 $X=7.89 $Y=1.37
c201 65 0 6.24044e-20 $X=1.22 $Y=1.37
c202 60 0 6.93685e-20 $X=7.805 $Y=1
c203 59 0 4.22339e-21 $X=1.22 $Y=1.255
c204 55 0 1.81152e-19 $X=7.89 $Y=1.27
c205 46 0 7.50258e-20 $X=0.87 $Y=2.26
c206 16 0 3.006e-19 $X=7.615 $Y=1.58
r207 63 68 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=7.89 $Y=1.255
+ $X2=7.89 $Y2=1.37
r208 62 63 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=7.89 $Y=1.085
+ $X2=7.89 $Y2=1.255
r209 60 62 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=7.805 $Y=1
+ $X2=7.89 $Y2=1.085
r210 60 61 6.25874 $w=1.7e-07 $l=6.5e-06 $layer=MET1_cond $X=7.805 $Y=1
+ $X2=1.305 $Y2=1
r211 59 65 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.22 $Y=1.255
+ $X2=1.22 $Y2=1.37
r212 58 61 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.22 $Y=1.085
+ $X2=1.305 $Y2=1
r213 58 59 0.16369 $w=1.7e-07 $l=1.7e-07 $layer=MET1_cond $X=1.22 $Y=1.085
+ $X2=1.22 $Y2=1.255
r214 57 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.89 $Y=1.37
+ $X2=7.89 $Y2=1.37
r215 55 57 4.51852 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=7.89 $Y=1.27 $X2=7.89
+ $Y2=1.37
r216 53 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.22 $Y=1.37
+ $X2=1.22 $Y2=1.37
r217 51 53 5.54545 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=1.26 $Y=1.27 $X2=1.26
+ $Y2=1.37
r218 48 49 8.89069 $w=2.47e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.19
+ $X2=0.87 $Y2=1.19
r219 44 46 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.26
+ $X2=0.87 $Y2=2.26
r220 43 49 5.39411 $w=2.47e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.955 $Y=1.27
+ $X2=0.87 $Y2=1.19
r221 42 51 2.2496 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.135 $Y=1.27
+ $X2=1.26 $Y2=1.27
r222 42 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.135 $Y=1.27
+ $X2=0.955 $Y2=1.27
r223 41 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.175
+ $X2=0.87 $Y2=2.26
r224 40 49 2.92482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=1.355
+ $X2=0.87 $Y2=1.19
r225 40 41 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.87 $Y=1.355
+ $X2=0.87 $Y2=2.175
r226 36 38 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.95
+ $X2=0.69 $Y2=3.63
r227 34 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.26
r228 34 36 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=0.69 $Y=2.345
+ $X2=0.69 $Y2=2.95
r229 30 48 2.92482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=1.19
r230 30 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=0.755
r231 29 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.27 $X2=7.89 $Y2=1.27
r232 24 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.27 $X2=1.22 $Y2=1.27
r233 24 26 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.22 $Y=1.27
+ $X2=1.425 $Y2=1.27
r234 20 29 38.9663 $w=3.64e-07 $l=2.07918e-07 $layer=POLY_cond $X=7.685 $Y=1.105
+ $X2=7.782 $Y2=1.27
r235 20 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.685 $Y=1.105
+ $X2=7.685 $Y2=0.785
r236 16 29 58.1668 $w=3.64e-07 $l=3.84539e-07 $layer=POLY_cond $X=7.615 $Y=1.58
+ $X2=7.782 $Y2=1.27
r237 16 18 956.309 $w=1.5e-07 $l=1.865e-06 $layer=POLY_cond $X=7.615 $Y=1.58
+ $X2=7.615 $Y2=3.445
r238 12 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.435
+ $X2=1.425 $Y2=1.27
r239 12 14 1030.66 $w=1.5e-07 $l=2.01e-06 $layer=POLY_cond $X=1.425 $Y=1.435
+ $X2=1.425 $Y2=3.445
r240 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.105
+ $X2=1.425 $Y2=1.27
r241 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=1.105
+ $X2=1.425 $Y2=0.785
r242 3 38 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=3.63
r243 3 36 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.605 $X2=0.69 $Y2=2.95
r244 1 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%A_342_442# 1 3 11 15 18 22 23 25 26 28
+ 31 36 38
c89 38 0 1.72079e-19 $X=3.365 $Y=0.755
r90 38 40 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=3.365 $Y=0.755
+ $X2=3.465 $Y2=0.755
r91 36 37 15.1353 $w=2.66e-07 $l=3.3e-07 $layer=LI1_cond $X=2.025 $Y=2.375
+ $X2=2.025 $Y2=2.705
r92 31 33 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=3.465 $Y=2.955
+ $X2=3.465 $Y2=3.635
r93 29 31 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=2.79
+ $X2=3.465 $Y2=2.955
r94 27 38 4.99104 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.365 $Y=0.935
+ $X2=3.365 $Y2=0.755
r95 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=0.935
+ $X2=3.365 $Y2=1.2
r96 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=1.285
+ $X2=3.365 $Y2=1.2
r97 25 26 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.28 $Y=1.285
+ $X2=2.2 $Y2=1.285
r98 24 37 3.35683 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.195 $Y=2.705
+ $X2=2.025 $Y2=2.705
r99 23 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.295 $Y=2.705
+ $X2=3.465 $Y2=2.79
r100 23 24 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.295 $Y=2.705
+ $X2=2.195 $Y2=2.705
r101 22 36 9.15133 $w=2.66e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.11 $Y=2.21
+ $X2=2.025 $Y2=2.375
r102 21 26 6.81649 $w=1.7e-07 $l=2.25555e-07 $layer=LI1_cond $X=2.11 $Y=1.47
+ $X2=2.2 $Y2=1.285
r103 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.11 $Y=1.47
+ $X2=2.11 $Y2=2.21
r104 18 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.375 $X2=1.94 $Y2=2.375
r105 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.375
+ $X2=1.892 $Y2=2.54
r106 18 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.375
+ $X2=1.892 $Y2=2.21
r107 15 19 730.691 $w=1.5e-07 $l=1.425e-06 $layer=POLY_cond $X=1.855 $Y=0.785
+ $X2=1.855 $Y2=2.21
r108 11 20 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.785 $Y=3.445
+ $X2=1.785 $Y2=2.54
r109 3 33 400 $w=1.7e-07 $l=1.13695e-06 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.605 $X2=3.465 $Y2=3.635
r110 3 31 400 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=2.605 $X2=3.465 $Y2=2.955
r111 1 40 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.575 $X2=3.465 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%D 3 7 10 14 19
c42 19 0 1.36979e-19 $X=2.865 $Y=1.74
c43 10 0 1.98306e-19 $X=2.865 $Y=1.74
r44 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.74
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.74 $X2=2.865 $Y2=1.74
r46 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.905
r47 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.74
+ $X2=2.865 $Y2=1.575
r48 7 12 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=2.805 $Y=3.235
+ $X2=2.805 $Y2=1.905
r49 3 11 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=2.805 $Y=0.85
+ $X2=2.805 $Y2=1.575
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%CK 3 7 10 13 15 17 18 20 23 25 29 30 33
+ 34 37 42 46 50 54 56 57 59 65 69 72 73 74 75 82
c250 75 0 1.48522e-19 $X=5.6 $Y=2.11
c251 73 0 1.48522e-19 $X=3.37 $Y=2.11
c252 72 0 1.89675e-19 $X=5.31 $Y=2.11
c253 59 0 3.12771e-20 $X=6.45 $Y=2.11
c254 57 0 6.91727e-20 $X=5.06 $Y=2.11
c255 56 0 8.3306e-20 $X=5.34 $Y=2.11
c256 50 0 3.67809e-19 $X=3.705 $Y=1.4
c257 46 0 1.89329e-19 $X=3.62 $Y=2.11
c258 37 0 1.16696e-19 $X=5.425 $Y=2.285
c259 25 0 1.36979e-19 $X=3.255 $Y=2.285
c260 18 0 1.37092e-19 $X=6.305 $Y=2.45
r261 75 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=2.11
+ $X2=5.455 $Y2=2.11
r262 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.305 $Y=2.11
+ $X2=6.45 $Y2=2.11
r263 74 75 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.305 $Y=2.11
+ $X2=5.6 $Y2=2.11
r264 73 77 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.37 $Y=2.11
+ $X2=3.225 $Y2=2.11
r265 72 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.31 $Y=2.11
+ $X2=5.455 $Y2=2.11
r266 72 73 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.31 $Y=2.11
+ $X2=3.37 $Y2=2.11
r267 69 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=2.11
+ $X2=5.455 $Y2=2.11
r268 69 71 11.7308 $w=1.82e-07 $l=1.75e-07 $layer=LI1_cond $X=5.44 $Y=2.11
+ $X2=5.44 $Y2=2.285
r269 65 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.225 $Y=2.11
+ $X2=3.225 $Y2=2.11
r270 65 67 11.7308 $w=1.82e-07 $l=1.75e-07 $layer=LI1_cond $X=3.24 $Y=2.11
+ $X2=3.24 $Y2=2.285
r271 59 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.45 $Y=2.11
+ $X2=6.45 $Y2=2.11
r272 59 62 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.45 $Y=2.11
+ $X2=6.45 $Y2=2.285
r273 56 69 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.34 $Y=2.11 $X2=5.44
+ $Y2=2.11
r274 56 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.34 $Y=2.11
+ $X2=5.06 $Y2=2.11
r275 52 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=2.025
+ $X2=5.06 $Y2=2.11
r276 52 54 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.975 $Y=2.025
+ $X2=4.975 $Y2=1.4
r277 48 50 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.705 $Y=2.025
+ $X2=3.705 $Y2=1.4
r278 47 65 1.129 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.34 $Y=2.11 $X2=3.24
+ $Y2=2.11
r279 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.11
+ $X2=3.705 $Y2=2.025
r280 46 47 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.62 $Y=2.11
+ $X2=3.34 $Y2=2.11
r281 45 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=2.285 $X2=6.45 $Y2=2.285
r282 40 42 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=6.305 $Y=1.28
+ $X2=6.385 $Y2=1.28
r283 37 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.425
+ $Y=2.285 $X2=5.425 $Y2=2.285
r284 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.425 $Y=2.285
+ $X2=5.425 $Y2=2.45
r285 33 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.4 $X2=4.975 $Y2=1.4
r286 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.4
+ $X2=4.975 $Y2=1.235
r287 29 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.4 $X2=3.705 $Y2=1.4
r288 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.4
+ $X2=3.705 $Y2=1.235
r289 25 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.255
+ $Y=2.285 $X2=3.255 $Y2=2.285
r290 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=2.285
+ $X2=3.255 $Y2=2.45
r291 23 45 38.571 $w=3.25e-07 $l=1.75656e-07 $layer=POLY_cond $X=6.385 $Y=2.12
+ $X2=6.407 $Y2=2.285
r292 22 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.385 $Y=1.355
+ $X2=6.385 $Y2=1.28
r293 22 23 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.385 $Y=1.355
+ $X2=6.385 $Y2=2.12
r294 18 45 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.305 $Y=2.45
+ $X2=6.407 $Y2=2.285
r295 18 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.305 $Y=2.45
+ $X2=6.305 $Y2=3.235
r296 15 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=1.28
r297 15 17 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.305 $Y=1.205
+ $X2=6.305 $Y2=0.85
r298 13 39 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.515 $Y=3.235
+ $X2=5.515 $Y2=2.45
r299 10 34 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.915 $Y=0.85
+ $X2=4.915 $Y2=1.235
r300 7 30 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.765 $Y=0.85
+ $X2=3.765 $Y2=1.235
r301 3 27 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.165 $Y=3.235
+ $X2=3.165 $Y2=2.45
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%A_217_605# 1 3 11 15 17 18 21 22 27 31
+ 35 37 38 41 44 47 50 56 57 62 64
c147 64 0 7.97351e-20 $X=4.205 $Y=1.37
c148 57 0 1.35571e-19 $X=4.06 $Y=1.37
c149 50 0 7.35919e-20 $X=1.65 $Y=1.37
c150 47 0 1.5821e-19 $X=4.295 $Y=2.285
c151 31 0 6.36774e-20 $X=4.555 $Y=3.235
c152 22 0 1.89329e-19 $X=4.2 $Y=2.285
c153 21 0 6.91727e-20 $X=4.48 $Y=2.285
c154 15 0 6.36774e-20 $X=4.125 $Y=3.235
r155 60 62 0.0994534 $w=2.35e-07 $l=1.4e-07 $layer=MET1_cond $X=1.65 $Y=1.367
+ $X2=1.79 $Y2=1.367
r156 57 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.37
+ $X2=4.205 $Y2=1.37
r157 57 62 2.18574 $w=1.7e-07 $l=2.27e-06 $layer=MET1_cond $X=4.06 $Y=1.37
+ $X2=1.79 $Y2=1.37
r158 54 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=1.37
+ $X2=4.205 $Y2=1.37
r159 54 56 5.43564 $w=2.02e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=1.345
+ $X2=4.295 $Y2=1.345
r160 50 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.65 $Y=1.37
+ $X2=1.65 $Y2=1.37
r161 50 52 7.13264 $w=1.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.645 $Y=1.37
+ $X2=1.645 $Y2=1.485
r162 50 51 7.44072 $w=1.78e-07 $l=1.2e-07 $layer=LI1_cond $X=1.645 $Y=1.37
+ $X2=1.645 $Y2=1.25
r163 45 56 1.74864 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.295 $Y=1.455
+ $X2=4.295 $Y2=1.345
r164 45 47 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.295 $Y=1.455
+ $X2=4.295 $Y2=2.285
r165 44 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.64 $Y=1.725
+ $X2=1.64 $Y2=1.485
r166 41 51 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.64 $Y=0.74
+ $X2=1.64 $Y2=1.25
r167 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.64 $Y2=1.725
r168 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.295 $Y2=1.81
r169 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.895
+ $X2=1.295 $Y2=1.81
r170 33 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.21 $Y=1.895
+ $X2=1.21 $Y2=3.275
r171 29 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.555 $Y=2.42
+ $X2=4.555 $Y2=3.235
r172 25 27 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.555 $Y=1.265
+ $X2=4.555 $Y2=0.85
r173 24 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=2.285 $X2=4.295 $Y2=2.285
r174 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=2.285
+ $X2=4.295 $Y2=2.285
r175 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=2.285
+ $X2=4.555 $Y2=2.42
r176 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=2.285
+ $X2=4.295 $Y2=2.285
r177 20 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.4 $X2=4.295 $Y2=1.4
r178 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=1.4
+ $X2=4.295 $Y2=1.4
r179 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.48 $Y=1.4
+ $X2=4.555 $Y2=1.265
r180 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=1.4
+ $X2=4.295 $Y2=1.4
r181 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=2.42
+ $X2=4.2 $Y2=2.285
r182 13 15 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.125 $Y=2.42
+ $X2=4.125 $Y2=3.235
r183 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=1.265
+ $X2=4.2 $Y2=1.4
r184 9 11 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.125 $Y=1.265
+ $X2=4.125 $Y2=0.85
r185 3 35 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=3.025 $X2=1.21 $Y2=3.275
r186 1 41 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%A_618_89# 1 3 9 11 13 14 15 18 20 24 26
+ 30 34 36 37 39 44 51 55 60 63 67 69 70 75
c199 75 0 1.37092e-19 $X=6.36 $Y=1.74
c200 70 0 4.17962e-19 $X=5.6 $Y=1.74
c201 69 0 2.9867e-19 $X=6.215 $Y=1.74
c202 51 0 5.69161e-20 $X=6.52 $Y=0.755
c203 44 0 1.89675e-19 $X=5.455 $Y=1.725
c204 34 0 1.69503e-19 $X=3.285 $Y=1.28
c205 24 0 1.48522e-19 $X=4.915 $Y=3.235
c206 18 0 1.48522e-19 $X=3.765 $Y=3.235
r207 70 72 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=1.74
+ $X2=5.455 $Y2=1.74
r208 69 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.215 $Y=1.74
+ $X2=6.36 $Y2=1.74
r209 69 70 0.592173 $w=1.7e-07 $l=6.15e-07 $layer=MET1_cond $X=6.215 $Y=1.74
+ $X2=5.6 $Y2=1.74
r210 65 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=2.705
+ $X2=6.795 $Y2=2.705
r211 63 64 17.474 $w=1.92e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=1.725
+ $X2=6.795 $Y2=1.725
r212 62 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.36 $Y=1.74
+ $X2=6.36 $Y2=1.74
r213 62 63 10.1667 $w=1.92e-07 $l=1.6e-07 $layer=LI1_cond $X=6.36 $Y=1.725
+ $X2=6.52 $Y2=1.725
r214 60 67 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.62
+ $X2=6.795 $Y2=2.705
r215 59 64 1.10697 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=6.795 $Y=1.825
+ $X2=6.795 $Y2=1.725
r216 59 60 48.9848 $w=1.78e-07 $l=7.95e-07 $layer=LI1_cond $X=6.795 $Y=1.825
+ $X2=6.795 $Y2=2.62
r217 55 57 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.52 $Y=2.955
+ $X2=6.52 $Y2=3.635
r218 53 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.79
+ $X2=6.52 $Y2=2.705
r219 53 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=2.79
+ $X2=6.52 $Y2=2.955
r220 49 63 1.44825 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.52 $Y=1.625 $X2=6.52
+ $Y2=1.725
r221 49 51 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.52 $Y=1.625
+ $X2=6.52 $Y2=0.755
r222 47 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=1.74
+ $X2=5.455 $Y2=1.74
r223 44 47 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.455 $Y=1.725
+ $X2=5.455 $Y2=1.74
r224 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.725 $X2=5.455 $Y2=1.725
r225 39 41 24.9945 $w=3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.47 $Y=1.725
+ $X2=5.47 $Y2=1.85
r226 39 40 55.9777 $w=3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.47 $Y=1.725
+ $X2=5.47 $Y2=1.52
r227 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.165 $Y=1.28
+ $X2=3.285 $Y2=1.28
r228 30 40 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.515 $Y=0.85
+ $X2=5.515 $Y2=1.52
r229 27 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.99 $Y=1.85
+ $X2=4.915 $Y2=1.85
r230 26 41 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.32 $Y=1.85
+ $X2=5.47 $Y2=1.85
r231 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.32 $Y=1.85
+ $X2=4.99 $Y2=1.85
r232 22 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.915 $Y=1.925
+ $X2=4.915 $Y2=1.85
r233 22 24 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=4.915 $Y=1.925
+ $X2=4.915 $Y2=3.235
r234 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.85
+ $X2=3.765 $Y2=1.85
r235 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=1.85
+ $X2=4.915 $Y2=1.85
r236 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.84 $Y=1.85 $X2=3.84
+ $Y2=1.85
r237 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.925
+ $X2=3.765 $Y2=1.85
r238 16 18 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=3.765 $Y=1.925
+ $X2=3.765 $Y2=3.235
r239 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=1.85
+ $X2=3.765 $Y2=1.85
r240 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.69 $Y=1.85
+ $X2=3.36 $Y2=1.85
r241 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.285 $Y=1.775
+ $X2=3.36 $Y2=1.85
r242 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.355
+ $X2=3.285 $Y2=1.28
r243 12 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.285 $Y=1.355
+ $X2=3.285 $Y2=1.775
r244 9 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.205
+ $X2=3.165 $Y2=1.28
r245 9 11 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=3.165 $Y=1.205
+ $X2=3.165 $Y2=0.85
r246 3 57 400 $w=1.7e-07 $l=1.09777e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=3.635
r247 3 55 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.605 $X2=6.52 $Y2=2.955
r248 1 51 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%A_1160_89# 1 3 11 14 26 29 30 31 32 33
+ 35 36 39 40 42 43 44 45 46 48 52 54 55 58 61 64 69 70 71 73 75 80 81
c210 44 0 8.77106e-20 $X=8.61 $Y=2.375
c211 40 0 1.81152e-19 $X=8.522 $Y=1.575
c212 39 0 3.51237e-19 $X=8.52 $Y=1.74
c213 36 0 1.31857e-19 $X=5.965 $Y=1.605
c214 35 0 2.19969e-19 $X=5.965 $Y=1.77
c215 33 0 1.50225e-19 $X=5.89 $Y=2.255
c216 31 0 2.82071e-19 $X=5.89 $Y=1.365
r217 80 81 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.52 $Y=1.74
+ $X2=8.375 $Y2=1.74
r218 75 81 1.32143 $w=1.75e-07 $l=1.46e-06 $layer=MET1_cond $X=6.915 $Y=1.737
+ $X2=8.375 $Y2=1.737
r219 72 75 0.0698591 $w=1.75e-07 $l=1.2657e-07 $layer=MET1_cond $X=6.825
+ $Y=1.825 $X2=6.915 $Y2=1.737
r220 72 73 0.501568 $w=1.8e-07 $l=5.7e-07 $layer=MET1_cond $X=6.825 $Y=1.825
+ $X2=6.825 $Y2=2.395
r221 71 77 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=2.48
+ $X2=5.935 $Y2=2.48
r222 70 73 0.0699153 $w=1.7e-07 $l=1.25499e-07 $layer=MET1_cond $X=6.735 $Y=2.48
+ $X2=6.825 $Y2=2.395
r223 70 71 0.630688 $w=1.7e-07 $l=6.55e-07 $layer=MET1_cond $X=6.735 $Y=2.48
+ $X2=6.08 $Y2=2.48
r224 64 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.52 $Y=1.74
+ $X2=8.52 $Y2=1.74
r225 62 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=1.74
+ $X2=7.47 $Y2=1.74
r226 62 64 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.555 $Y=1.74
+ $X2=8.52 $Y2=1.74
r227 60 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.825
+ $X2=7.47 $Y2=1.74
r228 60 61 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=7.47 $Y=1.825
+ $X2=7.47 $Y2=2.96
r229 56 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.655
+ $X2=7.47 $Y2=1.74
r230 56 58 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.47 $Y=1.655
+ $X2=7.47 $Y2=0.74
r231 54 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=3.045
+ $X2=7.47 $Y2=2.96
r232 54 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.385 $Y=3.045
+ $X2=7.125 $Y2=3.045
r233 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=3.13
+ $X2=7.125 $Y2=3.045
r234 50 52 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.04 $Y=3.13
+ $X2=7.04 $Y2=3.275
r235 48 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.935 $Y=2.48
+ $X2=5.935 $Y2=2.48
r236 46 68 17.1635 $w=1.82e-07 $l=2.62393e-07 $layer=LI1_cond $X=5.935 $Y=2.025
+ $X2=5.95 $Y2=1.77
r237 46 48 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.935 $Y=2.025
+ $X2=5.935 $Y2=2.48
r238 44 45 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=2.375
+ $X2=8.61 $Y2=2.525
r239 42 43 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=1.2 $X2=8.61
+ $Y2=1.35
r240 41 44 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=8.585 $Y=1.905
+ $X2=8.585 $Y2=2.375
r241 40 43 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.585 $Y=1.575
+ $X2=8.585 $Y2=1.35
r242 39 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.52
+ $Y=1.74 $X2=8.52 $Y2=1.74
r243 39 41 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.74
+ $X2=8.522 $Y2=1.905
r244 39 40 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=1.74
+ $X2=8.522 $Y2=1.575
r245 35 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.965
+ $Y=1.77 $X2=5.965 $Y2=1.77
r246 35 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=1.77
+ $X2=5.965 $Y2=1.935
r247 35 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=1.77
+ $X2=5.965 $Y2=1.605
r248 32 33 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.89 $Y=2.105
+ $X2=5.89 $Y2=2.255
r249 32 37 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.905 $Y=2.105
+ $X2=5.905 $Y2=1.935
r250 31 36 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.905 $Y=1.365
+ $X2=5.905 $Y2=1.605
r251 30 31 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=5.89 $Y=1.205
+ $X2=5.89 $Y2=1.365
r252 29 45 228.147 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=8.635 $Y=3.235
+ $X2=8.635 $Y2=2.525
r253 26 42 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=8.635 $Y=0.85
+ $X2=8.635 $Y2=1.2
r254 14 33 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=5.875 $Y=3.235
+ $X2=5.875 $Y2=2.255
r255 11 30 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=5.875 $Y=0.85
+ $X2=5.875 $Y2=1.205
r256 3 52 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=3.025 $X2=7.04 $Y2=3.275
r257 1 58 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.575 $X2=7.47 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%A_998_115# 1 3 11 15 18 23 25 26 29 33
+ 36 41 44 45 46 47 54
c146 47 0 2.65484e-19 $X=5.44 $Y=1.37
c147 46 0 3.12771e-20 $X=6.985 $Y=1.37
c148 45 0 1.5821e-19 $X=4.78 $Y=1.37
c149 41 0 1.71621e-19 $X=5.215 $Y=0.755
c150 36 0 1.69973e-19 $X=7.13 $Y=1.37
c151 33 0 1.66794e-19 $X=5.315 $Y=1.37
c152 23 0 1.57671e-19 $X=4.635 $Y=1.37
r153 47 52 0.0905432 $w=2.3e-07 $l=1.25e-07 $layer=MET1_cond $X=5.44 $Y=1.37
+ $X2=5.315 $Y2=1.37
r154 46 54 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=1.37
+ $X2=7.13 $Y2=1.37
r155 46 47 1.48765 $w=1.7e-07 $l=1.545e-06 $layer=MET1_cond $X=6.985 $Y=1.37
+ $X2=5.44 $Y2=1.37
r156 45 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.78 $Y=1.37
+ $X2=4.635 $Y2=1.37
r157 44 52 0.0969593 $w=2.3e-07 $l=1.35e-07 $layer=MET1_cond $X=5.18 $Y=1.37
+ $X2=5.315 $Y2=1.37
r158 44 45 0.385153 $w=1.7e-07 $l=4e-07 $layer=MET1_cond $X=5.18 $Y=1.37
+ $X2=4.78 $Y2=1.37
r159 41 43 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=5.222 $Y=0.755
+ $X2=5.222 $Y2=1.035
r160 36 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=1.37
+ $X2=7.13 $Y2=1.37
r161 33 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=1.37
+ $X2=5.315 $Y2=1.37
r162 33 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.315 $Y=1.37
+ $X2=5.315 $Y2=1.035
r163 27 29 17.1172 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=5.215 $Y=2.79
+ $X2=5.215 $Y2=3.295
r164 25 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=2.705
+ $X2=5.215 $Y2=2.79
r165 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=2.705
+ $X2=4.72 $Y2=2.705
r166 23 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.37
+ $X2=4.635 $Y2=1.37
r167 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=2.62
+ $X2=4.72 $Y2=2.705
r168 21 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.635 $Y=2.62
+ $X2=4.635 $Y2=1.37
r169 18 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.37 $X2=7.13 $Y2=1.37
r170 18 20 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=7.162 $Y=1.37
+ $X2=7.162 $Y2=1.535
r171 18 19 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=7.162 $Y=1.37
+ $X2=7.162 $Y2=1.205
r172 15 20 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=7.255 $Y=3.445
+ $X2=7.255 $Y2=1.535
r173 11 19 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=7.255 $Y=0.785
+ $X2=7.255 $Y2=1.205
r174 3 29 300 $w=1.7e-07 $l=7.94575e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.605 $X2=5.215 $Y2=3.295
r175 1 41 182 $w=1.7e-07 $l=3.01869e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.575 $X2=5.215 $Y2=0.755
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%QN 1 3 11 15 18 23 27 31 32 33 34 38 42
c85 42 0 8.77106e-20 $X=8.425 $Y=2.48
c86 33 0 1.02575e-19 $X=8.92 $Y=2.285
c87 31 0 1.18035e-19 $X=8.92 $Y=1.37
c88 18 0 1.98165e-19 $X=9.005 $Y=1.915
r89 40 42 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=8.42 $Y=2.48
+ $X2=8.425 $Y2=2.48
r90 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.005 $Y=2.2
+ $X2=9.005 $Y2=1.915
r91 35 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.005 $Y=1.455
+ $X2=9.005 $Y2=1.915
r92 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=2.285
+ $X2=9.005 $Y2=2.2
r93 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=2.285
+ $X2=8.505 $Y2=2.285
r94 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=1.37
+ $X2=9.005 $Y2=1.455
r95 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=1.37
+ $X2=8.505 $Y2=1.37
r96 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.48
r97 27 29 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=3.265
r98 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=2.37
+ $X2=8.505 $Y2=2.285
r99 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.42 $Y=2.37
+ $X2=8.42 $Y2=2.48
r100 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=1.285
+ $X2=8.505 $Y2=1.37
r101 21 23 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.42 $Y=1.285
+ $X2=8.42 $Y2=0.74
r102 18 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=1.915 $X2=9.005 $Y2=1.915
r103 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.915
+ $X2=9.005 $Y2=2.08
r104 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.915
+ $X2=9.005 $Y2=1.75
r105 15 20 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.065 $Y=3.235
+ $X2=9.065 $Y2=2.08
r106 11 19 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=9.065 $Y=0.85
+ $X2=9.065 $Y2=1.75
r107 3 29 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=2.605 $X2=8.42 $Y2=3.265
r108 1 23 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.575 $X2=8.42 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_HS__DFFR_1%Q 1 3 11 15 18 21 25 28
r19 25 26 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=2.807
+ $X2=9.395 $Y2=2.807
r20 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=2.85
+ $X2=9.275 $Y2=2.85
r21 24 25 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=9.275 $Y=2.807
+ $X2=9.28 $Y2=2.807
r22 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=1.035
+ $X2=9.395 $Y2=1.035
r23 18 26 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.395 $Y=2.68
+ $X2=9.395 $Y2=2.807
r24 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.12
+ $X2=9.395 $Y2=1.035
r25 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=9.395 $Y=1.12
+ $X2=9.395 $Y2=2.68
r26 13 25 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.28 $Y=2.935
+ $X2=9.28 $Y2=2.807
r27 13 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.28 $Y=2.935
+ $X2=9.28 $Y2=3.265
r28 9 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=0.95 $X2=9.28
+ $Y2=1.035
r29 9 11 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.28 $Y=0.95 $X2=9.28
+ $Y2=0.74
r30 3 15 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=2.605 $X2=9.28 $Y2=3.265
r31 1 11 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.575 $X2=9.28 $Y2=0.74
.ends

