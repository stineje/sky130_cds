* File: sky130_osu_sc_15T_ls__xor2_l.spice
* Created: Fri Nov 12 15:00:53 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__xor2_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__xor2_l  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1000 A_196_115# N_A_27_115#_M1000_g N_GND_M1002_d N_GND_M1002_b NSHORT L=0.15
+ W=0.74 AD=0.0777 AS=0.1036 PD=0.95 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A_238_89#_M1011_g A_196_115# N_GND_M1002_b NSHORT L=0.15
+ W=0.74 AD=0.1665 AS=0.0777 PD=1.19 PS=0.95 NRD=13.776 NRS=8.1 M=1 R=4.93333
+ SA=75001 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 A_388_115# N_A_M1007_g N_Y_M1011_d N_GND_M1002_b NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.1665 PD=0.95 PS=1.19 NRD=8.1 NRS=13.776 M=1 R=4.93333
+ SA=75001.6 SB=75001 A=0.111 P=1.78 MULT=1
MM1008 N_GND_M1008_d N_B_M1008_g A_388_115# N_GND_M1002_b NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.0777 PD=1.02 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75001.9
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1003 N_A_238_89#_M1003_d N_B_M1003_g N_GND_M1008_d N_GND_M1002_b NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75002.4 A=0.3 P=4.3 MULT=1
MM1005 A_196_565# N_A_M1005_g N_VDD_M1001_d N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.21 AS=0.28 PD=2.21 PS=2.28 NRD=4.9053 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75001.9 A=0.3 P=4.3 MULT=1
MM1006 N_Y_M1006_d N_A_238_89#_M1006_g A_196_565# N_VDD_M1001_b PHIGHVT L=0.15
+ W=2 AD=0.45 AS=0.21 PD=2.45 PS=2.21 NRD=8.3528 NRS=4.9053 M=1 R=13.3333
+ SA=75001 SB=75001.6 A=0.3 P=4.3 MULT=1
MM1010 A_388_565# N_A_27_115#_M1010_g N_Y_M1006_d N_VDD_M1001_b PHIGHVT L=0.15
+ W=2 AD=0.21 AS=0.45 PD=2.21 PS=2.45 NRD=4.9053 NRS=8.3528 M=1 R=13.3333
+ SA=75001.6 SB=75001 A=0.3 P=4.3 MULT=1
MM1009 N_VDD_M1009_d N_B_M1009_g A_388_565# N_VDD_M1001_b PHIGHVT L=0.15 W=2
+ AD=0.28 AS=0.21 PD=2.28 PS=2.21 NRD=0 NRS=4.9053 M=1 R=13.3333 SA=75001.9
+ SB=75000.6 A=0.3 P=4.3 MULT=1
MM1004 N_A_238_89#_M1004_d N_B_M1004_g N_VDD_M1009_d N_VDD_M1001_b PHIGHVT
+ L=0.15 W=2 AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75002.4 SB=75000.2 A=0.3 P=4.3 MULT=1
DX12_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=9.54325 P=12.37
pX13_noxref noxref_12 A A PROBETYPE=1
pX14_noxref noxref_13 Y Y PROBETYPE=1
pX15_noxref noxref_14 B B PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__xor2_l.pxi.spice"
*
.ends
*
*
