magic
tech sky130A
magscale 1 2
timestamp 1606864599
<< checkpaint >>
rect -1209 -1243 2161 2575
<< nwell >>
rect -9 581 990 1341
<< nmos >>
rect 80 115 110 315
rect 166 115 196 315
rect 252 115 282 315
rect 338 115 368 315
rect 424 115 454 315
rect 510 115 540 315
rect 596 115 626 315
rect 682 115 712 315
rect 768 115 798 315
rect 854 115 884 315
<< pmoshvt >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
rect 338 617 368 1217
rect 424 617 454 1217
rect 510 617 540 1217
rect 596 617 626 1217
rect 682 617 712 1217
rect 768 617 798 1217
rect 854 617 884 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 267 166 315
rect 110 131 121 267
rect 155 131 166 267
rect 110 115 166 131
rect 196 267 252 315
rect 196 131 207 267
rect 241 131 252 267
rect 196 115 252 131
rect 282 267 338 315
rect 282 131 293 267
rect 327 131 338 267
rect 282 115 338 131
rect 368 267 424 315
rect 368 131 379 267
rect 413 131 424 267
rect 368 115 424 131
rect 454 267 510 315
rect 454 131 465 267
rect 499 131 510 267
rect 454 115 510 131
rect 540 267 596 315
rect 540 131 551 267
rect 585 131 596 267
rect 540 115 596 131
rect 626 267 682 315
rect 626 131 637 267
rect 671 131 682 267
rect 626 115 682 131
rect 712 267 768 315
rect 712 131 723 267
rect 757 131 768 267
rect 712 115 768 131
rect 798 267 854 315
rect 798 131 809 267
rect 843 131 854 267
rect 798 115 854 131
rect 884 267 937 315
rect 884 131 895 267
rect 929 131 937 267
rect 884 115 937 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 725 35 1201
rect 69 725 80 1201
rect 27 617 80 725
rect 110 617 166 1217
rect 196 1201 252 1217
rect 196 793 207 1201
rect 241 793 252 1201
rect 196 617 252 793
rect 282 1201 338 1217
rect 282 657 293 1201
rect 327 657 338 1201
rect 282 617 338 657
rect 368 1201 424 1217
rect 368 657 379 1201
rect 413 657 424 1201
rect 368 617 424 657
rect 454 1201 510 1217
rect 454 657 465 1201
rect 499 657 510 1201
rect 454 617 510 657
rect 540 1201 596 1217
rect 540 657 551 1201
rect 585 657 596 1201
rect 540 617 596 657
rect 626 1201 682 1217
rect 626 657 637 1201
rect 671 657 682 1201
rect 626 617 682 657
rect 712 1201 768 1217
rect 712 657 723 1201
rect 757 657 768 1201
rect 712 617 768 657
rect 798 1201 854 1217
rect 798 657 809 1201
rect 843 657 854 1201
rect 798 617 854 657
rect 884 1201 937 1217
rect 884 657 895 1201
rect 929 657 937 1201
rect 884 617 937 657
<< ndiffc >>
rect 35 131 69 267
rect 121 131 155 267
rect 207 131 241 267
rect 293 131 327 267
rect 379 131 413 267
rect 465 131 499 267
rect 551 131 585 267
rect 637 131 671 267
rect 723 131 757 267
rect 809 131 843 267
rect 895 131 929 267
<< pdiffc >>
rect 35 725 69 1201
rect 207 793 241 1201
rect 293 657 327 1201
rect 379 657 413 1201
rect 465 657 499 1201
rect 551 657 585 1201
rect 637 657 671 1201
rect 723 657 757 1201
rect 809 657 843 1201
rect 895 657 929 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
rect 299 27 323 61
rect 357 27 381 61
rect 435 27 459 61
rect 493 27 517 61
rect 571 27 595 61
rect 629 27 653 61
rect 707 27 731 61
rect 765 27 789 61
rect 843 27 867 61
rect 901 27 925 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
rect 299 1271 323 1305
rect 357 1271 381 1305
rect 435 1271 459 1305
rect 493 1271 517 1305
rect 571 1271 595 1305
rect 629 1271 653 1305
rect 707 1271 731 1305
rect 765 1271 789 1305
rect 843 1271 867 1305
rect 901 1271 925 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
rect 323 27 357 61
rect 459 27 493 61
rect 595 27 629 61
rect 731 27 765 61
rect 867 27 901 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
rect 323 1271 357 1305
rect 459 1271 493 1305
rect 595 1271 629 1305
rect 731 1271 765 1305
rect 867 1271 901 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 338 1217 368 1244
rect 424 1217 454 1243
rect 510 1217 540 1243
rect 596 1217 626 1243
rect 682 1217 712 1243
rect 768 1217 798 1243
rect 854 1217 884 1243
rect 80 568 110 617
rect 27 552 110 568
rect 27 518 37 552
rect 71 518 110 552
rect 27 502 110 518
rect 166 510 196 617
rect 252 592 282 617
rect 338 592 368 617
rect 424 592 454 617
rect 510 592 540 617
rect 596 592 626 617
rect 682 592 712 617
rect 768 592 798 617
rect 854 592 884 617
rect 252 562 884 592
rect 80 315 110 502
rect 163 494 217 510
rect 163 460 173 494
rect 207 460 217 494
rect 163 444 217 460
rect 166 315 196 444
rect 259 420 289 562
rect 259 404 313 420
rect 259 384 269 404
rect 252 370 269 384
rect 303 384 313 404
rect 596 384 626 562
rect 303 370 884 384
rect 252 354 884 370
rect 252 315 282 354
rect 338 315 368 354
rect 424 315 454 354
rect 510 315 540 354
rect 596 315 626 354
rect 682 315 712 354
rect 768 315 798 354
rect 854 315 884 354
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
rect 338 89 368 115
rect 424 89 454 115
rect 510 89 540 115
rect 596 89 626 115
rect 682 89 712 115
rect 768 89 798 115
rect 854 89 884 115
<< polycont >>
rect 37 518 71 552
rect 173 460 207 494
rect 269 370 303 404
<< locali >>
rect 0 1311 990 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 323 1311
rect 357 1271 459 1311
rect 493 1271 595 1311
rect 629 1271 731 1311
rect 765 1271 867 1311
rect 901 1271 990 1311
rect 35 1201 69 1217
rect 207 1201 241 1271
rect 207 777 241 793
rect 293 1201 327 1217
rect 69 725 139 743
rect 35 709 139 725
rect 37 552 71 575
rect 37 502 71 518
rect 105 404 139 709
rect 173 494 207 649
rect 293 535 327 657
rect 379 1201 413 1271
rect 379 641 413 657
rect 465 1201 499 1217
rect 465 535 499 657
rect 551 1201 585 1271
rect 551 641 585 657
rect 637 1201 671 1217
rect 637 535 671 657
rect 723 1201 757 1271
rect 723 641 757 657
rect 809 1201 843 1217
rect 809 535 843 657
rect 895 1201 929 1271
rect 895 641 929 657
rect 173 444 207 460
rect 105 370 269 404
rect 303 370 319 404
rect 35 267 69 283
rect 35 61 69 131
rect 121 267 155 370
rect 121 115 155 131
rect 207 267 241 283
rect 207 61 241 131
rect 293 267 327 279
rect 293 115 327 131
rect 379 267 413 283
rect 379 61 413 131
rect 465 267 499 279
rect 465 115 499 131
rect 551 267 585 283
rect 551 61 585 131
rect 637 267 671 279
rect 637 115 671 131
rect 723 267 757 283
rect 723 61 757 131
rect 809 267 843 279
rect 809 115 843 131
rect 895 267 929 283
rect 895 61 929 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 323 61
rect 357 21 459 61
rect 493 21 595 61
rect 629 21 731 61
rect 765 21 867 61
rect 901 21 990 61
rect 0 0 990 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 323 1305 357 1311
rect 323 1277 357 1305
rect 459 1305 493 1311
rect 459 1277 493 1305
rect 595 1305 629 1311
rect 595 1277 629 1305
rect 731 1305 765 1311
rect 731 1277 765 1305
rect 867 1305 901 1311
rect 867 1277 901 1305
rect 37 575 71 609
rect 173 649 207 683
rect 293 501 327 535
rect 465 501 499 535
rect 637 501 671 535
rect 809 501 843 535
rect 293 279 327 313
rect 465 279 499 313
rect 637 279 671 313
rect 809 279 843 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
rect 323 27 357 55
rect 323 21 357 27
rect 459 27 493 55
rect 459 21 493 27
rect 595 27 629 55
rect 595 21 629 27
rect 731 27 765 55
rect 731 21 765 27
rect 867 27 901 55
rect 867 21 901 27
<< metal1 >>
rect 0 1311 990 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 323 1311
rect 357 1277 459 1311
rect 493 1277 595 1311
rect 629 1277 731 1311
rect 765 1277 867 1311
rect 901 1277 990 1311
rect 0 1271 990 1277
rect 161 683 219 689
rect 140 649 173 683
rect 207 649 219 683
rect 161 643 219 649
rect 25 609 83 615
rect 25 575 37 609
rect 71 575 105 609
rect 25 569 83 575
rect 281 535 339 541
rect 453 535 511 541
rect 625 535 683 541
rect 797 535 855 541
rect 281 501 293 535
rect 327 501 465 535
rect 499 501 637 535
rect 671 501 809 535
rect 843 501 855 535
rect 281 495 339 501
rect 453 495 511 501
rect 625 495 683 501
rect 797 495 855 501
rect 293 319 327 495
rect 465 319 499 495
rect 637 319 671 495
rect 809 319 843 495
rect 281 313 339 319
rect 453 313 511 319
rect 625 313 683 319
rect 797 313 855 319
rect 281 279 293 313
rect 327 279 465 313
rect 499 279 637 313
rect 671 279 683 313
rect 712 279 809 313
rect 843 279 855 313
rect 281 273 339 279
rect 453 273 511 279
rect 625 273 683 279
rect 797 273 855 279
rect 0 55 990 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 323 55
rect 357 21 459 55
rect 493 21 595 55
rect 629 21 731 55
rect 765 21 867 55
rect 901 21 990 55
rect 0 0 990 21
<< labels >>
rlabel metal1 311 444 311 444 1 Y
port 1 n
rlabel metal1 190 666 190 666 1 A
port 2 n
rlabel metal1 54 592 54 592 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
