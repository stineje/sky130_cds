* File: sky130_osu_sc_18T_ls__inv_l.pxi.spice
* Created: Thu Oct 29 17:36:54 2020
* 
x_PM_SKY130_OSU_SC_18T_LS__INV_L%GND N_GND_M1000_s N_GND_M1000_b N_GND_c_2_p GND
+ PM_SKY130_OSU_SC_18T_LS__INV_L%GND
x_PM_SKY130_OSU_SC_18T_LS__INV_L%VDD N_VDD_M1001_s N_VDD_M1001_b N_VDD_c_16_p
+ VDD N_VDD_c_18_p PM_SKY130_OSU_SC_18T_LS__INV_L%VDD
x_PM_SKY130_OSU_SC_18T_LS__INV_L%A N_A_M1000_g N_A_M1001_g N_A_c_29_n N_A_c_30_n
+ N_A_c_31_n A N_A_c_32_n PM_SKY130_OSU_SC_18T_LS__INV_L%A
x_PM_SKY130_OSU_SC_18T_LS__INV_L%Y N_Y_M1000_d N_Y_M1001_d Y N_Y_c_60_n
+ N_Y_c_61_n N_Y_c_62_n N_Y_c_63_n PM_SKY130_OSU_SC_18T_LS__INV_L%Y
cc_1 N_GND_M1000_b N_A_M1000_g 0.0996027f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.945
cc_2 N_GND_c_2_p N_A_M1000_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=0.945
cc_3 GND N_A_M1000_g 0.00468827f $X=0.34 $Y=0.22 $X2=0.475 $Y2=0.945
cc_4 N_GND_M1000_b N_A_M1001_g 0.0337175f $X=-0.045 $Y=0 $X2=0.475 $Y2=5.085
cc_5 N_GND_M1000_b N_A_c_29_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.305
cc_6 N_GND_M1000_b N_A_c_30_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_7 N_GND_M1000_b N_A_c_31_n 0.0393936f $X=-0.045 $Y=0 $X2=0.535 $Y2=2.305
cc_8 N_GND_M1000_b N_A_c_32_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=3.33
cc_9 N_GND_M1000_b Y 0.0587019f $X=-0.045 $Y=0 $X2=0.755 $Y2=2.205
cc_10 N_GND_M1000_b N_Y_c_60_n 0.0161674f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.48
cc_11 N_GND_M1000_b N_Y_c_61_n 0.00507896f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_12 N_GND_M1000_b N_Y_c_62_n 0.00237997f $X=-0.045 $Y=0 $X2=0.69 $Y2=2.96
cc_13 N_GND_M1000_b N_Y_c_63_n 0.0198055f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.825
cc_14 GND N_Y_c_63_n 0.00476261f $X=0.34 $Y=0.22 $X2=0.69 $Y2=0.825
cc_15 N_VDD_M1001_b N_A_M1001_g 0.108718f $X=-0.045 $Y=2.905 $X2=0.475 $Y2=5.085
cc_16 N_VDD_c_16_p N_A_M1001_g 0.00713292f $X=0.26 $Y=4.815 $X2=0.475 $Y2=5.085
cc_17 VDD N_A_M1001_g 0.00468827f $X=0.34 $Y=6.44 $X2=0.475 $Y2=5.085
cc_18 N_VDD_c_18_p N_A_M1001_g 0.00606474f $X=0.34 $Y=6.49 $X2=0.475 $Y2=5.085
cc_19 N_VDD_M1001_b A 0.0221642f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=3.33
cc_20 N_VDD_M1001_b N_A_c_32_n 0.0153337f $X=-0.045 $Y=2.905 $X2=0.32 $Y2=3.33
cc_21 N_VDD_M1001_b N_Y_c_61_n 0.00914195f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_22 N_VDD_M1001_b N_Y_c_62_n 0.0539944f $X=-0.045 $Y=2.905 $X2=0.69 $Y2=2.96
cc_23 VDD N_Y_c_62_n 0.00476261f $X=0.34 $Y=6.44 $X2=0.69 $Y2=2.96
cc_24 N_VDD_c_18_p N_Y_c_62_n 0.00757793f $X=0.34 $Y=6.49 $X2=0.69 $Y2=2.96
cc_25 N_A_M1000_g Y 0.0127139f $X=0.475 $Y=0.945 $X2=0.755 $Y2=2.205
cc_26 N_A_M1001_g Y 0.00874077f $X=0.475 $Y=5.085 $X2=0.755 $Y2=2.205
cc_27 N_A_c_30_n Y 0.0178517f $X=0.535 $Y=2.305 $X2=0.755 $Y2=2.205
cc_28 N_A_c_31_n Y 0.00719822f $X=0.535 $Y=2.305 $X2=0.755 $Y2=2.205
cc_29 N_A_c_32_n Y 0.0183799f $X=0.32 $Y=3.33 $X2=0.755 $Y2=2.205
cc_30 N_A_M1000_g N_Y_c_60_n 0.0119993f $X=0.475 $Y=0.945 $X2=0.69 $Y2=1.48
cc_31 N_A_c_31_n N_Y_c_60_n 0.0011424f $X=0.535 $Y=2.305 $X2=0.69 $Y2=1.48
cc_32 N_A_M1001_g N_Y_c_61_n 0.00478745f $X=0.475 $Y=5.085 $X2=0.69 $Y2=2.96
cc_33 N_A_c_30_n N_Y_c_61_n 0.00194461f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_34 N_A_c_31_n N_Y_c_61_n 0.00126139f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_35 A N_Y_c_61_n 0.00827053f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_36 N_A_c_32_n N_Y_c_61_n 0.00640429f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_37 N_A_M1001_g N_Y_c_62_n 0.0481998f $X=0.475 $Y=5.085 $X2=0.69 $Y2=2.96
cc_38 N_A_c_30_n N_Y_c_62_n 0.00202105f $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_39 N_A_c_31_n N_Y_c_62_n 8.13098e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=2.96
cc_40 A N_Y_c_62_n 0.0149533f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_41 N_A_c_32_n N_Y_c_62_n 0.0305887f $X=0.32 $Y=3.33 $X2=0.69 $Y2=2.96
cc_42 N_A_M1000_g N_Y_c_63_n 0.0152627f $X=0.475 $Y=0.945 $X2=0.69 $Y2=0.825
cc_43 N_A_c_30_n N_Y_c_63_n 0.00124107f $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
cc_44 N_A_c_31_n N_Y_c_63_n 6.24081e-19 $X=0.535 $Y=2.305 $X2=0.69 $Y2=0.825
