* File: sky130_osu_sc_15T_ls__buf_l.pxi.spice
* Created: Fri Nov 12 14:55:23 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__BUF_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_15T_LS__BUF_L%GND
x_PM_SKY130_OSU_SC_15T_LS__BUF_L%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_27_p
+ N_VDD_c_28_p N_VDD_c_34_p VDD N_VDD_c_29_p PM_SKY130_OSU_SC_15T_LS__BUF_L%VDD
x_PM_SKY130_OSU_SC_15T_LS__BUF_L%A N_A_M1002_g N_A_M1001_g N_A_c_49_n N_A_c_50_n
+ A PM_SKY130_OSU_SC_15T_LS__BUF_L%A
x_PM_SKY130_OSU_SC_15T_LS__BUF_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_M1003_g N_A_27_115#_c_83_n
+ N_A_27_115#_c_84_n N_A_27_115#_c_85_n N_A_27_115#_c_86_n N_A_27_115#_c_89_n
+ N_A_27_115#_c_90_n N_A_27_115#_c_91_n N_A_27_115#_c_92_n
+ PM_SKY130_OSU_SC_15T_LS__BUF_L%A_27_115#
x_PM_SKY130_OSU_SC_15T_LS__BUF_L%Y N_Y_M1000_d N_Y_M1003_d N_Y_c_133_n
+ N_Y_c_138_n Y N_Y_c_136_n N_Y_c_137_n PM_SKY130_OSU_SC_15T_LS__BUF_L%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.0712812f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.835
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.835
cc_3 N_GND_c_3_p N_A_M1002_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.835
cc_4 N_GND_c_4_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.835
cc_5 N_GND_M1002_b N_A_M1001_g 0.0156812f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.195
cc_6 N_GND_M1002_b N_A_c_49_n 0.040771f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.22
cc_7 N_GND_M1002_b N_A_c_50_n 0.00595324f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.22
cc_8 N_GND_M1002_b N_A_27_115#_M1000_g 0.0488034f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.835
cc_9 N_GND_c_3_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905
+ $Y2=0.835
cc_10 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=0.835
cc_11 N_GND_M1002_b N_A_27_115#_c_83_n 0.0597491f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.6
cc_12 N_GND_M1002_b N_A_27_115#_c_84_n 0.0562401f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=1.675
cc_13 N_GND_M1002_b N_A_27_115#_c_85_n 0.0168393f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.675
cc_14 N_GND_M1002_b N_A_27_115#_c_86_n 0.0251493f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_15 N_GND_c_2_p N_A_27_115#_c_86_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_16 N_GND_c_4_p N_A_27_115#_c_86_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_17 N_GND_M1002_b N_A_27_115#_c_89_n 0.0412202f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=4.28
cc_18 N_GND_M1002_b N_A_27_115#_c_90_n 0.0172272f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.675
cc_19 N_GND_M1002_b N_A_27_115#_c_91_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.675
cc_20 N_GND_M1002_b N_A_27_115#_c_92_n 0.00663593f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.675
cc_21 N_GND_M1002_b N_Y_c_133_n 0.0178338f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.74
cc_22 N_GND_c_4_p N_Y_c_133_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.12 $Y2=0.74
cc_23 N_GND_M1002_b Y 0.0164841f $X=-0.045 $Y=0 $X2=1.07 $Y2=2
cc_24 N_GND_M1002_b N_Y_c_136_n 0.014537f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.22
cc_25 N_GND_M1002_b N_Y_c_137_n 0.00501078f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.7
cc_26 N_VDD_M1001_b N_A_M1001_g 0.0675162f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=4.195
cc_27 N_VDD_c_27_p N_A_M1001_g 0.00496961f $X=0.605 $Y=5.397 $X2=0.475 $Y2=4.195
cc_28 N_VDD_c_28_p N_A_M1001_g 0.00316701f $X=0.69 $Y=4.28 $X2=0.475 $Y2=4.195
cc_29 N_VDD_c_29_p N_A_M1001_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=4.195
cc_30 N_VDD_M1001_b N_A_c_50_n 0.011209f $X=-0.045 $Y=2.645 $X2=0.635 $Y2=2.22
cc_31 N_VDD_M1001_b A 0.0157561f $X=-0.045 $Y=2.645 $X2=0.635 $Y2=3.07
cc_32 N_VDD_M1001_b N_A_27_115#_M1003_g 0.0614257f $X=-0.045 $Y=2.645 $X2=0.905
+ $Y2=4.195
cc_33 N_VDD_c_28_p N_A_27_115#_M1003_g 0.00316701f $X=0.69 $Y=4.28 $X2=0.905
+ $Y2=4.195
cc_34 N_VDD_c_34_p N_A_27_115#_M1003_g 0.00496961f $X=1.02 $Y=5.33 $X2=0.905
+ $Y2=4.195
cc_35 N_VDD_c_29_p N_A_27_115#_M1003_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.905
+ $Y2=4.195
cc_36 N_VDD_M1001_b N_A_27_115#_c_85_n 0.0187682f $X=-0.045 $Y=2.645 $X2=1.18
+ $Y2=2.675
cc_37 N_VDD_M1001_b N_A_27_115#_c_89_n 0.0455808f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=4.28
cc_38 N_VDD_c_27_p N_A_27_115#_c_89_n 0.00452684f $X=0.605 $Y=5.397 $X2=0.26
+ $Y2=4.28
cc_39 N_VDD_c_29_p N_A_27_115#_c_89_n 0.00435496f $X=1.02 $Y=5.36 $X2=0.26
+ $Y2=4.28
cc_40 N_VDD_M1001_b N_Y_c_138_n 0.038618f $X=-0.045 $Y=2.645 $X2=1.12 $Y2=2.7
cc_41 N_VDD_c_34_p N_Y_c_138_n 0.00452684f $X=1.02 $Y=5.33 $X2=1.12 $Y2=2.7
cc_42 N_VDD_c_29_p N_Y_c_138_n 0.00435496f $X=1.02 $Y=5.36 $X2=1.12 $Y2=2.7
cc_43 N_VDD_M1001_b N_Y_c_137_n 0.0107503f $X=-0.045 $Y=2.645 $X2=1.12 $Y2=2.7
cc_44 N_A_M1002_g N_A_27_115#_M1000_g 0.0439177f $X=0.475 $Y=0.835 $X2=0.905
+ $Y2=0.835
cc_45 A N_A_27_115#_M1003_g 0.00419145f $X=0.635 $Y=3.07 $X2=0.905 $Y2=4.195
cc_46 N_A_M1002_g N_A_27_115#_c_83_n 0.00260138f $X=0.475 $Y=0.835 $X2=1.18
+ $Y2=2.6
cc_47 N_A_M1001_g N_A_27_115#_c_83_n 0.00209773f $X=0.475 $Y=4.195 $X2=1.18
+ $Y2=2.6
cc_48 N_A_c_49_n N_A_27_115#_c_83_n 0.0139096f $X=0.635 $Y=2.22 $X2=1.18 $Y2=2.6
cc_49 N_A_c_50_n N_A_27_115#_c_83_n 0.00361737f $X=0.635 $Y=2.22 $X2=1.18
+ $Y2=2.6
cc_50 N_A_M1001_g N_A_27_115#_c_85_n 0.0653954f $X=0.475 $Y=4.195 $X2=1.18
+ $Y2=2.675
cc_51 N_A_c_50_n N_A_27_115#_c_85_n 0.00468272f $X=0.635 $Y=2.22 $X2=1.18
+ $Y2=2.675
cc_52 N_A_M1002_g N_A_27_115#_c_86_n 0.0212724f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=0.74
cc_53 N_A_M1002_g N_A_27_115#_c_89_n 0.0620725f $X=0.475 $Y=0.835 $X2=0.26
+ $Y2=4.28
cc_54 N_A_c_50_n N_A_27_115#_c_89_n 0.0696932f $X=0.635 $Y=2.22 $X2=0.26
+ $Y2=4.28
cc_55 A N_A_27_115#_c_89_n 0.0155137f $X=0.635 $Y=3.07 $X2=0.26 $Y2=4.28
cc_56 N_A_M1002_g N_A_27_115#_c_90_n 0.0207696f $X=0.475 $Y=0.835 $X2=0.88
+ $Y2=1.675
cc_57 N_A_c_49_n N_A_27_115#_c_90_n 0.00273049f $X=0.635 $Y=2.22 $X2=0.88
+ $Y2=1.675
cc_58 N_A_c_50_n N_A_27_115#_c_90_n 0.00886797f $X=0.635 $Y=2.22 $X2=0.88
+ $Y2=1.675
cc_59 N_A_M1002_g N_A_27_115#_c_92_n 6.59135e-19 $X=0.475 $Y=0.835 $X2=0.965
+ $Y2=1.675
cc_60 N_A_c_50_n N_Y_c_138_n 0.0203054f $X=0.635 $Y=2.22 $X2=1.12 $Y2=2.7
cc_61 A N_Y_c_138_n 0.00731851f $X=0.635 $Y=3.07 $X2=1.12 $Y2=2.7
cc_62 N_A_M1002_g Y 0.00310306f $X=0.475 $Y=0.835 $X2=1.07 $Y2=2
cc_63 N_A_c_49_n Y 0.00441844f $X=0.635 $Y=2.22 $X2=1.07 $Y2=2
cc_64 N_A_c_50_n Y 0.0200396f $X=0.635 $Y=2.22 $X2=1.07 $Y2=2
cc_65 N_A_M1002_g N_Y_c_136_n 0.00102215f $X=0.475 $Y=0.835 $X2=1.12 $Y2=1.22
cc_66 N_A_c_50_n N_Y_c_137_n 0.00609526f $X=0.635 $Y=2.22 $X2=1.12 $Y2=2.7
cc_67 N_A_27_115#_M1000_g N_Y_c_133_n 0.0100708f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=0.74
cc_68 N_A_27_115#_c_84_n N_Y_c_133_n 0.00477112f $X=1.18 $Y=1.675 $X2=1.12
+ $Y2=0.74
cc_69 N_A_27_115#_c_92_n N_Y_c_133_n 7.50437e-19 $X=0.965 $Y=1.675 $X2=1.12
+ $Y2=0.74
cc_70 N_A_27_115#_M1003_g N_Y_c_138_n 0.0355152f $X=0.905 $Y=4.195 $X2=1.12
+ $Y2=2.7
cc_71 N_A_27_115#_c_85_n N_Y_c_138_n 0.0134943f $X=1.18 $Y=2.675 $X2=1.12
+ $Y2=2.7
cc_72 N_A_27_115#_M1000_g Y 0.00406656f $X=0.905 $Y=0.835 $X2=1.07 $Y2=2
cc_73 N_A_27_115#_c_83_n Y 0.0310322f $X=1.18 $Y=2.6 $X2=1.07 $Y2=2
cc_74 N_A_27_115#_c_84_n Y 0.0161039f $X=1.18 $Y=1.675 $X2=1.07 $Y2=2
cc_75 N_A_27_115#_c_90_n Y 8.73078e-19 $X=0.88 $Y=1.675 $X2=1.07 $Y2=2
cc_76 N_A_27_115#_c_92_n Y 0.0121742f $X=0.965 $Y=1.675 $X2=1.07 $Y2=2
cc_77 N_A_27_115#_M1000_g N_Y_c_136_n 0.00714414f $X=0.905 $Y=0.835 $X2=1.12
+ $Y2=1.22
cc_78 N_A_27_115#_c_84_n N_Y_c_136_n 0.0014753f $X=1.18 $Y=1.675 $X2=1.12
+ $Y2=1.22
cc_79 N_A_27_115#_c_92_n N_Y_c_136_n 0.00278861f $X=0.965 $Y=1.675 $X2=1.12
+ $Y2=1.22
cc_80 N_A_27_115#_M1003_g N_Y_c_137_n 0.0015856f $X=0.905 $Y=4.195 $X2=1.12
+ $Y2=2.7
cc_81 N_A_27_115#_c_83_n N_Y_c_137_n 0.00226191f $X=1.18 $Y=2.6 $X2=1.12 $Y2=2.7
cc_82 N_A_27_115#_c_85_n N_Y_c_137_n 0.00513726f $X=1.18 $Y=2.675 $X2=1.12
+ $Y2=2.7
