* File: sky130_osu_sc_18T_ls__and2_4.pxi.spice
* Created: Fri Nov 12 13:39:14 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__AND2_4%GND N_GND_M1001_d N_GND_M1008_s N_GND_M1011_s
+ N_GND_M1005_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p N_GND_c_22_p N_GND_c_30_p
+ N_GND_c_36_p GND N_GND_c_3_p PM_SKY130_OSU_SC_18T_LS__AND2_4%GND
x_PM_SKY130_OSU_SC_18T_LS__AND2_4%VDD N_VDD_M1004_s N_VDD_M1010_d N_VDD_M1003_d
+ N_VDD_M1007_d N_VDD_M1004_b N_VDD_c_75_p N_VDD_c_76_p N_VDD_c_87_p
+ N_VDD_c_94_p N_VDD_c_100_p N_VDD_c_106_p N_VDD_c_111_p VDD N_VDD_c_77_p
+ PM_SKY130_OSU_SC_18T_LS__AND2_4%VDD
x_PM_SKY130_OSU_SC_18T_LS__AND2_4%A N_A_M1005_g N_A_M1004_g N_A_c_130_n
+ N_A_c_131_n A PM_SKY130_OSU_SC_18T_LS__AND2_4%A
x_PM_SKY130_OSU_SC_18T_LS__AND2_4%B N_B_M1001_g N_B_M1010_g N_B_c_164_n
+ N_B_c_165_n B PM_SKY130_OSU_SC_18T_LS__AND2_4%B
x_PM_SKY130_OSU_SC_18T_LS__AND2_4%A_27_115# N_A_27_115#_M1005_s
+ N_A_27_115#_M1004_d N_A_27_115#_M1000_g N_A_27_115#_c_237_n
+ N_A_27_115#_M1002_g N_A_27_115#_c_204_n N_A_27_115#_c_205_n
+ N_A_27_115#_M1008_g N_A_27_115#_c_242_n N_A_27_115#_M1003_g
+ N_A_27_115#_c_210_n N_A_27_115#_c_212_n N_A_27_115#_c_213_n
+ N_A_27_115#_M1009_g N_A_27_115#_c_249_n N_A_27_115#_M1006_g
+ N_A_27_115#_c_218_n N_A_27_115#_c_219_n N_A_27_115#_M1011_g
+ N_A_27_115#_c_254_n N_A_27_115#_M1007_g N_A_27_115#_c_224_n
+ N_A_27_115#_c_225_n N_A_27_115#_c_226_n N_A_27_115#_c_227_n
+ N_A_27_115#_c_228_n N_A_27_115#_c_231_n N_A_27_115#_c_232_n
+ N_A_27_115#_c_261_n N_A_27_115#_c_233_n N_A_27_115#_c_235_n
+ N_A_27_115#_c_236_n N_A_27_115#_c_277_n
+ PM_SKY130_OSU_SC_18T_LS__AND2_4%A_27_115#
x_PM_SKY130_OSU_SC_18T_LS__AND2_4%Y N_Y_M1000_d N_Y_M1009_d N_Y_M1002_s
+ N_Y_M1006_s N_Y_c_335_n N_Y_c_340_n N_Y_c_341_n N_Y_c_345_n N_Y_c_346_n
+ N_Y_c_349_n Y N_Y_c_351_n N_Y_c_353_n N_Y_c_354_n N_Y_c_357_n
+ PM_SKY130_OSU_SC_18T_LS__AND2_4%Y
cc_1 N_GND_M1005_b N_A_M1005_g 0.0806078f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_A_M1005_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_A_M1005_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=1.075
cc_4 N_GND_M1005_b N_A_c_130_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.765
cc_5 N_GND_M1005_b N_A_c_131_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.765
cc_6 N_GND_M1005_b N_B_M1001_g 0.0460664f $X=-0.045 $Y=0 $X2=0.835 $Y2=1.075
cc_7 N_GND_c_2_p N_B_M1001_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=1.075
cc_8 N_GND_c_8_p N_B_M1001_g 0.00376152f $X=1.05 $Y=0.825 $X2=0.835 $Y2=1.075
cc_9 N_GND_c_3_p N_B_M1001_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.835 $Y2=1.075
cc_10 N_GND_M1005_b N_B_M1010_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_11 N_GND_M1005_b N_B_c_164_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_12 N_GND_M1005_b N_B_c_165_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.425
cc_13 N_GND_M1005_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.96
cc_14 N_GND_M1005_b N_A_27_115#_M1000_g 0.0215719f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_15 N_GND_c_8_p N_A_27_115#_M1000_g 0.0103278f $X=1.05 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_16 N_GND_c_16_p N_A_27_115#_M1000_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_c_3_p N_A_27_115#_M1000_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.335
+ $Y2=1.075
cc_18 N_GND_M1005_b N_A_27_115#_c_204_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.81
cc_19 N_GND_M1005_b N_A_27_115#_c_205_n 0.00954592f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.885
cc_20 N_GND_M1005_b N_A_27_115#_M1008_g 0.0202142f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_21 N_GND_c_16_p N_A_27_115#_M1008_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=1.075
cc_22 N_GND_c_22_p N_A_27_115#_M1008_g 0.00356864f $X=1.98 $Y=0.825 $X2=1.765
+ $Y2=1.075
cc_23 N_GND_c_3_p N_A_27_115#_M1008_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.765
+ $Y2=1.075
cc_24 N_GND_M1005_b N_A_27_115#_c_210_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.845
cc_25 N_GND_c_22_p N_A_27_115#_c_210_n 0.00256938f $X=1.98 $Y=0.825 $X2=2.12
+ $Y2=1.845
cc_26 N_GND_M1005_b N_A_27_115#_c_212_n 0.0448266f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.845
cc_27 N_GND_M1005_b N_A_27_115#_c_213_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.885
cc_28 N_GND_M1005_b N_A_27_115#_M1009_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.075
cc_29 N_GND_c_22_p N_A_27_115#_M1009_g 0.00356864f $X=1.98 $Y=0.825 $X2=2.195
+ $Y2=1.075
cc_30 N_GND_c_30_p N_A_27_115#_M1009_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=1.075
cc_31 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.195
+ $Y2=1.075
cc_32 N_GND_M1005_b N_A_27_115#_c_218_n 0.0369419f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.845
cc_33 N_GND_M1005_b N_A_27_115#_c_219_n 0.0268552f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.885
cc_34 N_GND_M1005_b N_A_27_115#_M1011_g 0.0264941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.075
cc_35 N_GND_c_30_p N_A_27_115#_M1011_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=1.075
cc_36 N_GND_c_36_p N_A_27_115#_M1011_g 0.00713292f $X=2.84 $Y=0.825 $X2=2.625
+ $Y2=1.075
cc_37 N_GND_c_3_p N_A_27_115#_M1011_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.625
+ $Y2=1.075
cc_38 N_GND_M1005_b N_A_27_115#_c_224_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.885
cc_39 N_GND_M1005_b N_A_27_115#_c_225_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.885
cc_40 N_GND_M1005_b N_A_27_115#_c_226_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.845
cc_41 N_GND_M1005_b N_A_27_115#_c_227_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.885
cc_42 N_GND_M1005_b N_A_27_115#_c_228_n 0.0143389f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.825
cc_43 N_GND_c_2_p N_A_27_115#_c_228_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.825
cc_44 N_GND_c_3_p N_A_27_115#_c_228_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.825
cc_45 N_GND_M1005_b N_A_27_115#_c_231_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.935
cc_46 N_GND_M1005_b N_A_27_115#_c_232_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.935
cc_47 N_GND_M1005_b N_A_27_115#_c_233_n 0.0230268f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_48 N_GND_c_8_p N_A_27_115#_c_233_n 0.00704977f $X=1.05 $Y=0.825 $X2=1.43
+ $Y2=1.935
cc_49 N_GND_M1005_b N_A_27_115#_c_235_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.935
cc_50 N_GND_M1005_b N_A_27_115#_c_236_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.545
cc_51 N_GND_M1005_b N_Y_c_335_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_52 N_GND_c_8_p N_Y_c_335_n 0.0187614f $X=1.05 $Y=0.825 $X2=1.55 $Y2=0.825
cc_53 N_GND_c_16_p N_Y_c_335_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.825
cc_54 N_GND_c_22_p N_Y_c_335_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=0.825
cc_55 N_GND_c_3_p N_Y_c_335_n 0.00475776f $X=2.38 $Y=0.19 $X2=1.55 $Y2=0.825
cc_56 N_GND_M1005_b N_Y_c_340_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_57 N_GND_M1005_b N_Y_c_341_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.825
cc_58 N_GND_c_22_p N_Y_c_341_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=0.825
cc_59 N_GND_c_30_p N_Y_c_341_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.825
cc_60 N_GND_c_3_p N_Y_c_341_n 0.00475776f $X=2.38 $Y=0.19 $X2=2.41 $Y2=0.825
cc_61 N_GND_M1005_b N_Y_c_345_n 0.0152877f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.59
cc_62 N_GND_M1005_b N_Y_c_346_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.595
cc_63 N_GND_c_8_p N_Y_c_346_n 0.00127231f $X=1.05 $Y=0.825 $X2=1.55 $Y2=1.595
cc_64 N_GND_c_22_p N_Y_c_346_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=1.595
cc_65 N_GND_M1005_b N_Y_c_349_n 0.00463624f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.475
cc_66 N_GND_M1005_b Y 0.0306813f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_67 N_GND_M1008_s N_Y_c_351_n 0.0127884f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.48
cc_68 N_GND_c_22_p N_Y_c_351_n 0.0142303f $X=1.98 $Y=0.825 $X2=2.265 $Y2=1.48
cc_69 N_GND_M1005_b N_Y_c_353_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.59
cc_70 N_GND_M1005_b N_Y_c_354_n 0.00409378f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.595
cc_71 N_GND_c_22_p N_Y_c_354_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=1.595
cc_72 N_GND_c_36_p N_Y_c_354_n 0.00134236f $X=2.84 $Y=0.825 $X2=2.41 $Y2=1.595
cc_73 N_GND_M1005_b N_Y_c_357_n 0.06145f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.475
cc_74 N_VDD_M1004_b N_A_M1004_g 0.0189471f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_75 N_VDD_c_75_p N_A_M1004_g 0.00713292f $X=0.26 $Y=4.135 $X2=0.475 $Y2=4.585
cc_76 N_VDD_c_76_p N_A_M1004_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=4.585
cc_77 N_VDD_c_77_p N_A_M1004_g 0.00468827f $X=2.38 $Y=6.47 $X2=0.475 $Y2=4.585
cc_78 N_VDD_M1004_b N_A_c_130_n 0.0111025f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=2.765
cc_79 N_VDD_M1004_s N_A_c_131_n 0.0127298f $X=0.135 $Y=3.085 $X2=0.27 $Y2=2.765
cc_80 N_VDD_M1004_b N_A_c_131_n 0.00612103f $X=-0.045 $Y=2.905 $X2=0.27
+ $Y2=2.765
cc_81 N_VDD_c_75_p N_A_c_131_n 0.00370742f $X=0.26 $Y=4.135 $X2=0.27 $Y2=2.765
cc_82 N_VDD_M1004_s A 0.00742066f $X=0.135 $Y=3.085 $X2=0.275 $Y2=3.33
cc_83 N_VDD_M1004_b A 0.00970321f $X=-0.045 $Y=2.905 $X2=0.275 $Y2=3.33
cc_84 N_VDD_c_75_p A 0.00434783f $X=0.26 $Y=4.135 $X2=0.275 $Y2=3.33
cc_85 N_VDD_M1004_b N_B_M1010_g 0.0187476f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_86 N_VDD_c_76_p N_B_M1010_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=4.585
cc_87 N_VDD_c_87_p N_B_M1010_g 0.00354579f $X=1.12 $Y=3.795 $X2=0.905 $Y2=4.585
cc_88 N_VDD_c_77_p N_B_M1010_g 0.00468827f $X=2.38 $Y=6.47 $X2=0.905 $Y2=4.585
cc_89 N_VDD_M1004_b N_B_c_165_n 0.00170274f $X=-0.045 $Y=2.905 $X2=0.95
+ $Y2=2.425
cc_90 N_VDD_M1004_b B 0.00856863f $X=-0.045 $Y=2.905 $X2=0.955 $Y2=2.96
cc_91 N_VDD_c_87_p B 0.00240671f $X=1.12 $Y=3.795 $X2=0.955 $Y2=2.96
cc_92 N_VDD_M1004_b N_A_27_115#_c_237_n 0.017104f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.96
cc_93 N_VDD_c_87_p N_A_27_115#_c_237_n 0.00354579f $X=1.12 $Y=3.795 $X2=1.335
+ $Y2=2.96
cc_94 N_VDD_c_94_p N_A_27_115#_c_237_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.335
+ $Y2=2.96
cc_95 N_VDD_c_77_p N_A_27_115#_c_237_n 0.00468827f $X=2.38 $Y=6.47 $X2=1.335
+ $Y2=2.96
cc_96 N_VDD_M1004_b N_A_27_115#_c_205_n 0.00428234f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.885
cc_97 N_VDD_M1004_b N_A_27_115#_c_242_n 0.017006f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.96
cc_98 N_VDD_c_87_p N_A_27_115#_c_242_n 3.67508e-19 $X=1.12 $Y=3.795 $X2=1.765
+ $Y2=2.96
cc_99 N_VDD_c_94_p N_A_27_115#_c_242_n 0.00610567f $X=1.895 $Y=6.507 $X2=1.765
+ $Y2=2.96
cc_100 N_VDD_c_100_p N_A_27_115#_c_242_n 0.00373985f $X=1.98 $Y=3.455 $X2=1.765
+ $Y2=2.96
cc_101 N_VDD_c_77_p N_A_27_115#_c_242_n 0.00470215f $X=2.38 $Y=6.47 $X2=1.765
+ $Y2=2.96
cc_102 N_VDD_M1004_b N_A_27_115#_c_213_n 0.00396043f $X=-0.045 $Y=2.905 $X2=2.12
+ $Y2=2.885
cc_103 N_VDD_c_100_p N_A_27_115#_c_213_n 0.00379272f $X=1.98 $Y=3.455 $X2=2.12
+ $Y2=2.885
cc_104 N_VDD_M1004_b N_A_27_115#_c_249_n 0.0166898f $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.96
cc_105 N_VDD_c_100_p N_A_27_115#_c_249_n 0.00354579f $X=1.98 $Y=3.455 $X2=2.195
+ $Y2=2.96
cc_106 N_VDD_c_106_p N_A_27_115#_c_249_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.195
+ $Y2=2.96
cc_107 N_VDD_c_77_p N_A_27_115#_c_249_n 0.00468827f $X=2.38 $Y=6.47 $X2=2.195
+ $Y2=2.96
cc_108 N_VDD_M1004_b N_A_27_115#_c_219_n 0.00840215f $X=-0.045 $Y=2.905 $X2=2.55
+ $Y2=2.885
cc_109 N_VDD_M1004_b N_A_27_115#_c_254_n 0.0209036f $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=2.96
cc_110 N_VDD_c_106_p N_A_27_115#_c_254_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.625
+ $Y2=2.96
cc_111 N_VDD_c_111_p N_A_27_115#_c_254_n 0.00713292f $X=2.84 $Y=3.455 $X2=2.625
+ $Y2=2.96
cc_112 N_VDD_c_77_p N_A_27_115#_c_254_n 0.00468827f $X=2.38 $Y=6.47 $X2=2.625
+ $Y2=2.96
cc_113 N_VDD_M1004_b N_A_27_115#_c_224_n 0.0021704f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.885
cc_114 N_VDD_M1004_b N_A_27_115#_c_225_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.885
cc_115 N_VDD_M1004_b N_A_27_115#_c_227_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.885
cc_116 N_VDD_M1004_b N_A_27_115#_c_261_n 0.00155118f $X=-0.045 $Y=2.905 $X2=0.69
+ $Y2=3.795
cc_117 N_VDD_c_76_p N_A_27_115#_c_261_n 0.0075556f $X=1.035 $Y=6.507 $X2=0.69
+ $Y2=3.795
cc_118 N_VDD_c_77_p N_A_27_115#_c_261_n 0.00475776f $X=2.38 $Y=6.47 $X2=0.69
+ $Y2=3.795
cc_119 N_VDD_M1004_b N_A_27_115#_c_236_n 8.22047e-19 $X=-0.045 $Y=2.905 $X2=0.65
+ $Y2=3.545
cc_120 N_VDD_M1004_b N_Y_c_340_n 0.00344954f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=2.59
cc_121 N_VDD_c_94_p N_Y_c_340_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55 $Y2=2.59
cc_122 N_VDD_c_77_p N_Y_c_340_n 0.00475776f $X=2.38 $Y=6.47 $X2=1.55 $Y2=2.59
cc_123 N_VDD_M1004_b N_Y_c_345_n 0.00380347f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.59
cc_124 N_VDD_c_106_p N_Y_c_345_n 0.00734006f $X=2.755 $Y=6.507 $X2=2.41 $Y2=2.59
cc_125 N_VDD_c_77_p N_Y_c_345_n 0.00475776f $X=2.38 $Y=6.47 $X2=2.41 $Y2=2.59
cc_126 N_VDD_c_100_p N_Y_c_353_n 0.00634153f $X=1.98 $Y=3.455 $X2=2.265 $Y2=2.59
cc_127 N_A_M1005_g N_B_M1001_g 0.129148f $X=0.475 $Y=1.075 $X2=0.835 $Y2=1.075
cc_128 N_A_M1005_g N_B_M1010_g 0.0498038f $X=0.475 $Y=1.075 $X2=0.905 $Y2=4.585
cc_129 N_A_M1005_g N_B_c_165_n 7.8234e-19 $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.425
cc_130 N_A_M1005_g N_A_27_115#_c_228_n 0.0158058f $X=0.475 $Y=1.075 $X2=0.26
+ $Y2=0.825
cc_131 N_A_M1005_g N_A_27_115#_c_231_n 0.0160984f $X=0.475 $Y=1.075 $X2=0.525
+ $Y2=1.935
cc_132 N_A_c_130_n N_A_27_115#_c_231_n 0.00117122f $X=0.475 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_133 N_A_c_131_n N_A_27_115#_c_231_n 2.65873e-19 $X=0.27 $Y=2.765 $X2=0.525
+ $Y2=1.935
cc_134 N_A_c_130_n N_A_27_115#_c_232_n 0.00133457f $X=0.475 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_135 N_A_c_131_n N_A_27_115#_c_232_n 0.0055861f $X=0.27 $Y=2.765 $X2=0.345
+ $Y2=1.935
cc_136 N_A_M1005_g N_A_27_115#_c_235_n 0.00322084f $X=0.475 $Y=1.075 $X2=0.61
+ $Y2=1.935
cc_137 N_A_M1005_g N_A_27_115#_c_236_n 0.0265302f $X=0.475 $Y=1.075 $X2=0.65
+ $Y2=3.545
cc_138 N_A_M1004_g N_A_27_115#_c_236_n 0.0140172f $X=0.475 $Y=4.585 $X2=0.65
+ $Y2=3.545
cc_139 N_A_c_130_n N_A_27_115#_c_236_n 0.00766302f $X=0.475 $Y=2.765 $X2=0.65
+ $Y2=3.545
cc_140 N_A_c_131_n N_A_27_115#_c_236_n 0.0456533f $X=0.27 $Y=2.765 $X2=0.65
+ $Y2=3.545
cc_141 A N_A_27_115#_c_236_n 0.00758489f $X=0.275 $Y=3.33 $X2=0.65 $Y2=3.545
cc_142 N_A_M1004_g N_A_27_115#_c_277_n 0.00884152f $X=0.475 $Y=4.585 $X2=0.65
+ $Y2=3.715
cc_143 N_B_M1001_g N_A_27_115#_M1000_g 0.0349978f $X=0.835 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_144 N_B_M1010_g N_A_27_115#_c_204_n 0.00773101f $X=0.905 $Y=4.585 $X2=1.37
+ $Y2=2.81
cc_145 N_B_c_164_n N_A_27_115#_c_204_n 0.0206104f $X=0.95 $Y=2.425 $X2=1.37
+ $Y2=2.81
cc_146 N_B_c_165_n N_A_27_115#_c_204_n 0.0033451f $X=0.95 $Y=2.425 $X2=1.37
+ $Y2=2.81
cc_147 N_B_M1001_g N_A_27_115#_c_212_n 0.0104742f $X=0.835 $Y=1.075 $X2=1.84
+ $Y2=1.845
cc_148 N_B_M1010_g N_A_27_115#_c_224_n 0.0401773f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.885
cc_149 N_B_c_165_n N_A_27_115#_c_224_n 0.00173699f $X=0.95 $Y=2.425 $X2=1.352
+ $Y2=2.885
cc_150 B N_A_27_115#_c_224_n 0.00389258f $X=0.955 $Y=2.96 $X2=1.352 $Y2=2.885
cc_151 N_B_M1001_g N_A_27_115#_c_233_n 0.0182215f $X=0.835 $Y=1.075 $X2=1.43
+ $Y2=1.935
cc_152 N_B_c_164_n N_A_27_115#_c_233_n 0.00258465f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_153 N_B_c_165_n N_A_27_115#_c_233_n 0.0101796f $X=0.95 $Y=2.425 $X2=1.43
+ $Y2=1.935
cc_154 N_B_M1001_g N_A_27_115#_c_236_n 0.00755919f $X=0.835 $Y=1.075 $X2=0.65
+ $Y2=3.545
cc_155 N_B_M1010_g N_A_27_115#_c_236_n 0.0133197f $X=0.905 $Y=4.585 $X2=0.65
+ $Y2=3.545
cc_156 N_B_c_165_n N_A_27_115#_c_236_n 0.0541375f $X=0.95 $Y=2.425 $X2=0.65
+ $Y2=3.545
cc_157 B N_A_27_115#_c_236_n 0.00866797f $X=0.955 $Y=2.96 $X2=0.65 $Y2=3.545
cc_158 B N_A_27_115#_c_277_n 0.00286715f $X=0.955 $Y=2.96 $X2=0.65 $Y2=3.715
cc_159 N_B_c_165_n N_Y_c_340_n 0.0149875f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.59
cc_160 B N_Y_c_340_n 0.00649253f $X=0.955 $Y=2.96 $X2=1.55 $Y2=2.59
cc_161 N_B_M1001_g N_Y_c_346_n 8.18972e-19 $X=0.835 $Y=1.075 $X2=1.55 $Y2=1.595
cc_162 N_B_c_164_n N_Y_c_349_n 5.85867e-19 $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.475
cc_163 N_B_c_165_n N_Y_c_349_n 0.00592261f $X=0.95 $Y=2.425 $X2=1.55 $Y2=2.475
cc_164 N_B_M1001_g Y 6.71108e-19 $X=0.835 $Y=1.075 $X2=1.555 $Y2=2.22
cc_165 N_B_c_165_n Y 0.00695761f $X=0.95 $Y=2.425 $X2=1.555 $Y2=2.22
cc_166 N_A_27_115#_M1000_g N_Y_c_335_n 0.00233629f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_167 N_A_27_115#_M1008_g N_Y_c_335_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_168 N_A_27_115#_c_212_n N_Y_c_335_n 0.00171364f $X=1.84 $Y=1.845 $X2=1.55
+ $Y2=0.825
cc_169 N_A_27_115#_c_233_n N_Y_c_335_n 0.00500271f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_170 N_A_27_115#_c_237_n N_Y_c_340_n 0.00278785f $X=1.335 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_171 N_A_27_115#_c_204_n N_Y_c_340_n 0.00744772f $X=1.37 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_172 N_A_27_115#_c_205_n N_Y_c_340_n 0.0167599f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.59
cc_173 N_A_27_115#_c_242_n N_Y_c_340_n 0.00392729f $X=1.765 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_174 N_A_27_115#_c_212_n N_Y_c_340_n 0.0013767f $X=1.84 $Y=1.845 $X2=1.55
+ $Y2=2.59
cc_175 N_A_27_115#_c_233_n N_Y_c_340_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_176 N_A_27_115#_M1009_g N_Y_c_341_n 0.00231637f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_177 N_A_27_115#_c_218_n N_Y_c_341_n 0.00280419f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=0.825
cc_178 N_A_27_115#_M1011_g N_Y_c_341_n 0.00231637f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_179 N_A_27_115#_c_249_n N_Y_c_345_n 0.00392729f $X=2.195 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_180 N_A_27_115#_c_218_n N_Y_c_345_n 0.00250559f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.59
cc_181 N_A_27_115#_c_219_n N_Y_c_345_n 0.0206674f $X=2.55 $Y=2.885 $X2=2.41
+ $Y2=2.59
cc_182 N_A_27_115#_c_254_n N_Y_c_345_n 0.00392729f $X=2.625 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_183 N_A_27_115#_M1000_g N_Y_c_346_n 0.00554705f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_184 N_A_27_115#_M1008_g N_Y_c_346_n 0.00259902f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_185 N_A_27_115#_c_233_n N_Y_c_346_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.595
cc_186 N_A_27_115#_c_204_n N_Y_c_349_n 0.00821104f $X=1.37 $Y=2.81 $X2=1.55
+ $Y2=2.475
cc_187 N_A_27_115#_c_205_n N_Y_c_349_n 0.00229755f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.475
cc_188 N_A_27_115#_c_212_n N_Y_c_349_n 0.00174847f $X=1.84 $Y=1.845 $X2=1.55
+ $Y2=2.475
cc_189 N_A_27_115#_c_233_n N_Y_c_349_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.475
cc_190 N_A_27_115#_M1000_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_191 N_A_27_115#_c_204_n Y 0.00892438f $X=1.37 $Y=2.81 $X2=1.555 $Y2=2.22
cc_192 N_A_27_115#_M1008_g Y 0.00251111f $X=1.765 $Y=1.075 $X2=1.555 $Y2=2.22
cc_193 N_A_27_115#_c_212_n Y 0.0128645f $X=1.84 $Y=1.845 $X2=1.555 $Y2=2.22
cc_194 N_A_27_115#_c_233_n Y 0.0148238f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_195 N_A_27_115#_M1008_g N_Y_c_351_n 0.0130095f $X=1.765 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_196 N_A_27_115#_c_210_n N_Y_c_351_n 0.00213861f $X=2.12 $Y=1.845 $X2=2.265
+ $Y2=1.48
cc_197 N_A_27_115#_M1009_g N_Y_c_351_n 0.0130095f $X=2.195 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_198 N_A_27_115#_c_212_n N_Y_c_353_n 0.0121767f $X=1.84 $Y=1.845 $X2=2.265
+ $Y2=2.59
cc_199 N_A_27_115#_c_225_n N_Y_c_353_n 0.0158479f $X=1.765 $Y=2.885 $X2=2.265
+ $Y2=2.59
cc_200 N_A_27_115#_M1009_g N_Y_c_354_n 0.00259902f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=1.595
cc_201 N_A_27_115#_M1011_g N_Y_c_354_n 0.00939545f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=1.595
cc_202 N_A_27_115#_M1009_g N_Y_c_357_n 0.00251111f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_203 N_A_27_115#_c_218_n N_Y_c_357_n 0.0184054f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.475
cc_204 N_A_27_115#_M1011_g N_Y_c_357_n 0.00251111f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_205 N_A_27_115#_c_226_n N_Y_c_357_n 0.00140336f $X=2.195 $Y=1.845 $X2=2.41
+ $Y2=2.475
cc_206 N_A_27_115#_c_227_n N_Y_c_357_n 0.00372651f $X=2.195 $Y=2.885 $X2=2.41
+ $Y2=2.475
