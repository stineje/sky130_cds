* File: sky130_osu_sc_12T_ms__inv_4.pxi.spice
* Created: Fri Nov 12 15:24:30 2021
* 
x_PM_SKY130_OSU_SC_12T_MS__INV_4%GND N_GND_M1000_d N_GND_M1001_d N_GND_M1007_d
+ N_GND_M1000_b N_GND_c_2_p N_GND_c_3_p N_GND_c_10_p N_GND_c_17_p N_GND_c_23_p
+ GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_MS__INV_4%GND
x_PM_SKY130_OSU_SC_12T_MS__INV_4%VDD N_VDD_M1002_s N_VDD_M1004_s N_VDD_M1006_s
+ N_VDD_M1002_b N_VDD_c_59_p N_VDD_c_60_p N_VDD_c_65_p N_VDD_c_71_p N_VDD_c_76_p
+ VDD N_VDD_c_61_p PM_SKY130_OSU_SC_12T_MS__INV_4%VDD
x_PM_SKY130_OSU_SC_12T_MS__INV_4%A N_A_c_97_n N_A_M1000_g N_A_c_101_n
+ N_A_c_132_n N_A_M1002_g N_A_c_102_n N_A_c_103_n N_A_c_104_n N_A_M1001_g
+ N_A_c_137_n N_A_M1004_g N_A_c_108_n N_A_c_110_n N_A_c_111_n N_A_M1003_g
+ N_A_c_143_n N_A_M1005_g N_A_c_115_n N_A_c_116_n N_A_c_117_n N_A_M1007_g
+ N_A_c_148_n N_A_M1006_g N_A_c_121_n N_A_c_122_n N_A_c_123_n N_A_c_124_n
+ N_A_c_125_n N_A_c_126_n N_A_c_127_n N_A_c_128_n N_A_c_129_n N_A_c_130_n
+ N_A_c_131_n A PM_SKY130_OSU_SC_12T_MS__INV_4%A
x_PM_SKY130_OSU_SC_12T_MS__INV_4%Y N_Y_M1000_s N_Y_M1003_s N_Y_M1002_d
+ N_Y_M1005_d N_Y_c_217_n N_Y_c_239_n N_Y_c_221_n N_Y_c_242_n N_Y_c_225_n
+ N_Y_c_245_n Y N_Y_c_230_n N_Y_c_246_n N_Y_c_234_n N_Y_c_238_n
+ PM_SKY130_OSU_SC_12T_MS__INV_4%Y
cc_1 N_GND_M1000_b N_A_c_97_n 0.0208613f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.22
cc_2 N_GND_c_2_p N_A_c_97_n 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=1.22
cc_3 N_GND_c_3_p N_A_c_97_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.22
cc_4 N_GND_c_4_p N_A_c_97_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.475 $Y2=1.22
cc_5 N_GND_M1000_b N_A_c_101_n 0.0262237f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.33
cc_6 N_GND_M1000_b N_A_c_102_n 0.0162043f $X=-0.045 $Y=0 $X2=0.83 $Y2=1.295
cc_7 N_GND_M1000_b N_A_c_103_n 0.0114349f $X=-0.045 $Y=0 $X2=0.83 $Y2=2.405
cc_8 N_GND_M1000_b N_A_c_104_n 0.0166526f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.22
cc_9 N_GND_c_3_p N_A_c_104_n 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.22
cc_10 N_GND_c_10_p N_A_c_104_n 0.00311745f $X=1.12 $Y=0.755 $X2=0.905 $Y2=1.22
cc_11 N_GND_c_4_p N_A_c_104_n 0.00468827f $X=1.7 $Y=0.19 $X2=0.905 $Y2=1.22
cc_12 N_GND_M1000_b N_A_c_108_n 0.0213783f $X=-0.045 $Y=0 $X2=1.26 $Y2=1.295
cc_13 N_GND_c_10_p N_A_c_108_n 0.00283047f $X=1.12 $Y=0.755 $X2=1.26 $Y2=1.295
cc_14 N_GND_M1000_b N_A_c_110_n 0.0173499f $X=-0.045 $Y=0 $X2=1.26 $Y2=2.405
cc_15 N_GND_M1000_b N_A_c_111_n 0.0166526f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.22
cc_16 N_GND_c_10_p N_A_c_111_n 0.00311745f $X=1.12 $Y=0.755 $X2=1.335 $Y2=1.22
cc_17 N_GND_c_17_p N_A_c_111_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.335 $Y2=1.22
cc_18 N_GND_c_4_p N_A_c_111_n 0.00468827f $X=1.7 $Y=0.19 $X2=1.335 $Y2=1.22
cc_19 N_GND_M1000_b N_A_c_115_n 0.0385034f $X=-0.045 $Y=0 $X2=1.69 $Y2=1.295
cc_20 N_GND_M1000_b N_A_c_116_n 0.0295863f $X=-0.045 $Y=0 $X2=1.69 $Y2=2.405
cc_21 N_GND_M1000_b N_A_c_117_n 0.0208613f $X=-0.045 $Y=0 $X2=1.765 $Y2=1.22
cc_22 N_GND_c_17_p N_A_c_117_n 0.00606474f $X=1.895 $Y=0.152 $X2=1.765 $Y2=1.22
cc_23 N_GND_c_23_p N_A_c_117_n 0.00502587f $X=1.98 $Y=0.755 $X2=1.765 $Y2=1.22
cc_24 N_GND_c_4_p N_A_c_117_n 0.00468827f $X=1.7 $Y=0.19 $X2=1.765 $Y2=1.22
cc_25 N_GND_M1000_b N_A_c_121_n 0.0106787f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.295
cc_26 N_GND_M1000_b N_A_c_122_n 0.0348407f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_27 N_GND_M1000_b N_A_c_123_n 0.0276572f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.66
cc_28 N_GND_M1000_b N_A_c_124_n 0.00422354f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.405
cc_29 N_GND_M1000_b N_A_c_125_n 0.0106787f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.295
cc_30 N_GND_M1000_b N_A_c_126_n 0.00980309f $X=-0.045 $Y=0 $X2=0.905 $Y2=2.405
cc_31 N_GND_M1000_b N_A_c_127_n 0.0106787f $X=-0.045 $Y=0 $X2=1.335 $Y2=1.295
cc_32 N_GND_M1000_b N_A_c_128_n 0.00980309f $X=-0.045 $Y=0 $X2=1.335 $Y2=2.405
cc_33 N_GND_M1000_b N_A_c_129_n 0.0176577f $X=-0.045 $Y=0 $X2=0.32 $Y2=2.85
cc_34 N_GND_M1000_b N_A_c_130_n 0.0132529f $X=-0.045 $Y=0 $X2=0.405 $Y2=1.825
cc_35 N_GND_M1000_b N_A_c_131_n 0.00267654f $X=-0.045 $Y=0 $X2=0.535 $Y2=1.825
cc_36 N_GND_M1000_b N_Y_c_217_n 0.00154299f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.755
cc_37 N_GND_c_3_p N_Y_c_217_n 0.00740081f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.755
cc_38 N_GND_c_10_p N_Y_c_217_n 8.14297e-19 $X=1.12 $Y=0.755 $X2=0.69 $Y2=0.755
cc_39 N_GND_c_4_p N_Y_c_217_n 0.0047139f $X=1.7 $Y=0.19 $X2=0.69 $Y2=0.755
cc_40 N_GND_M1000_b N_Y_c_221_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_41 N_GND_c_10_p N_Y_c_221_n 8.14297e-19 $X=1.12 $Y=0.755 $X2=1.55 $Y2=0.755
cc_42 N_GND_c_17_p N_Y_c_221_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_43 N_GND_c_4_p N_Y_c_221_n 0.0047139f $X=1.7 $Y=0.19 $X2=1.55 $Y2=0.755
cc_44 N_GND_M1000_b N_Y_c_225_n 0.00294733f $X=-0.045 $Y=0 $X2=0.69 $Y2=1.115
cc_45 N_GND_c_2_p N_Y_c_225_n 0.00134236f $X=0.26 $Y=0.755 $X2=0.69 $Y2=1.115
cc_46 N_GND_c_3_p N_Y_c_225_n 0.00245319f $X=1.035 $Y=0.152 $X2=0.69 $Y2=1.115
cc_47 N_GND_c_10_p N_Y_c_225_n 7.53951e-19 $X=1.12 $Y=0.755 $X2=0.69 $Y2=1.115
cc_48 N_GND_M1000_b Y 0.0456345f $X=-0.045 $Y=0 $X2=0.76 $Y2=1.72
cc_49 N_GND_M1001_d N_Y_c_230_n 0.0100144f $X=0.98 $Y=0.575 $X2=1.405 $Y2=1
cc_50 N_GND_c_3_p N_Y_c_230_n 0.0028844f $X=1.035 $Y=0.152 $X2=1.405 $Y2=1
cc_51 N_GND_c_10_p N_Y_c_230_n 0.0142303f $X=1.12 $Y=0.755 $X2=1.405 $Y2=1
cc_52 N_GND_c_17_p N_Y_c_230_n 0.0028844f $X=1.895 $Y=0.152 $X2=1.405 $Y2=1
cc_53 N_GND_M1000_b N_Y_c_234_n 0.00409378f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.115
cc_54 N_GND_c_10_p N_Y_c_234_n 7.53951e-19 $X=1.12 $Y=0.755 $X2=1.55 $Y2=1.115
cc_55 N_GND_c_17_p N_Y_c_234_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.55 $Y2=1.115
cc_56 N_GND_c_23_p N_Y_c_234_n 0.00134236f $X=1.98 $Y=0.755 $X2=1.55 $Y2=1.115
cc_57 N_GND_M1000_b N_Y_c_238_n 0.0754129f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.365
cc_58 N_VDD_M1002_b N_A_c_132_n 0.0181616f $X=-0.045 $Y=2.425 $X2=0.475 $Y2=2.48
cc_59 N_VDD_c_59_p N_A_c_132_n 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=2.48
cc_60 N_VDD_c_60_p N_A_c_132_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=2.48
cc_61 N_VDD_c_61_p N_A_c_132_n 0.00468827f $X=1.7 $Y=4.25 $X2=0.475 $Y2=2.48
cc_62 N_VDD_M1002_b N_A_c_103_n 0.00448664f $X=-0.045 $Y=2.425 $X2=0.83
+ $Y2=2.405
cc_63 N_VDD_M1002_b N_A_c_137_n 0.0159283f $X=-0.045 $Y=2.425 $X2=0.905 $Y2=2.48
cc_64 N_VDD_c_60_p N_A_c_137_n 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=2.48
cc_65 N_VDD_c_65_p N_A_c_137_n 0.00337744f $X=1.12 $Y=2.955 $X2=0.905 $Y2=2.48
cc_66 N_VDD_c_61_p N_A_c_137_n 0.00468827f $X=1.7 $Y=4.25 $X2=0.905 $Y2=2.48
cc_67 N_VDD_M1002_b N_A_c_110_n 0.00500158f $X=-0.045 $Y=2.425 $X2=1.26
+ $Y2=2.405
cc_68 N_VDD_c_65_p N_A_c_110_n 0.00341318f $X=1.12 $Y=2.955 $X2=1.26 $Y2=2.405
cc_69 N_VDD_M1002_b N_A_c_143_n 0.0159283f $X=-0.045 $Y=2.425 $X2=1.335 $Y2=2.48
cc_70 N_VDD_c_65_p N_A_c_143_n 0.00337744f $X=1.12 $Y=2.955 $X2=1.335 $Y2=2.48
cc_71 N_VDD_c_71_p N_A_c_143_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335 $Y2=2.48
cc_72 N_VDD_c_61_p N_A_c_143_n 0.00468827f $X=1.7 $Y=4.25 $X2=1.335 $Y2=2.48
cc_73 N_VDD_M1002_b N_A_c_116_n 0.00840215f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_74 N_VDD_M1002_b N_A_c_148_n 0.0204783f $X=-0.045 $Y=2.425 $X2=1.765 $Y2=2.48
cc_75 N_VDD_c_71_p N_A_c_148_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.765 $Y2=2.48
cc_76 N_VDD_c_76_p N_A_c_148_n 0.00636672f $X=1.98 $Y=2.955 $X2=1.765 $Y2=2.48
cc_77 N_VDD_c_61_p N_A_c_148_n 0.00468827f $X=1.7 $Y=4.25 $X2=1.765 $Y2=2.48
cc_78 N_VDD_M1002_b N_A_c_124_n 0.00244521f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.405
cc_79 N_VDD_M1002_b N_A_c_126_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=2.405
cc_80 N_VDD_M1002_b N_A_c_128_n 8.75564e-19 $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.405
cc_81 N_VDD_M1002_s N_A_c_129_n 0.00953431f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.85
cc_82 N_VDD_M1002_b N_A_c_129_n 0.00618364f $X=-0.045 $Y=2.425 $X2=0.32 $Y2=2.85
cc_83 N_VDD_c_59_p N_A_c_129_n 0.00252874f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.85
cc_84 N_VDD_M1002_s A 0.0162774f $X=0.135 $Y=2.605 $X2=0.32 $Y2=2.845
cc_85 N_VDD_c_59_p A 0.00522047f $X=0.26 $Y=3.635 $X2=0.32 $Y2=2.845
cc_86 N_VDD_c_65_p A 9.09141e-19 $X=1.12 $Y=2.955 $X2=0.32 $Y2=2.845
cc_87 N_VDD_M1002_b N_Y_c_239_n 0.00361433f $X=-0.045 $Y=2.425 $X2=0.69 $Y2=2.48
cc_88 N_VDD_c_60_p N_Y_c_239_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69 $Y2=2.48
cc_89 N_VDD_c_61_p N_Y_c_239_n 0.00475776f $X=1.7 $Y=4.25 $X2=0.69 $Y2=2.48
cc_90 N_VDD_M1002_b N_Y_c_242_n 0.00465961f $X=-0.045 $Y=2.425 $X2=1.55 $Y2=2.48
cc_91 N_VDD_c_71_p N_Y_c_242_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.48
cc_92 N_VDD_c_61_p N_Y_c_242_n 0.00475776f $X=1.7 $Y=4.25 $X2=1.55 $Y2=2.48
cc_93 N_VDD_M1002_b N_Y_c_245_n 0.00248543f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=2.365
cc_94 N_VDD_M1002_b N_Y_c_246_n 0.00520877f $X=-0.045 $Y=2.425 $X2=1.405
+ $Y2=2.48
cc_95 N_VDD_c_65_p N_Y_c_246_n 0.0090257f $X=1.12 $Y=2.955 $X2=1.405 $Y2=2.48
cc_96 N_VDD_M1002_b N_Y_c_238_n 0.00409378f $X=-0.045 $Y=2.425 $X2=1.55
+ $Y2=2.365
cc_97 A N_Y_M1002_d 0.00250716f $X=0.32 $Y=2.845 $X2=0.55 $Y2=2.605
cc_98 N_A_c_97_n N_Y_c_217_n 0.00182852f $X=0.475 $Y=1.22 $X2=0.69 $Y2=0.755
cc_99 N_A_c_102_n N_Y_c_217_n 0.00251439f $X=0.83 $Y=1.295 $X2=0.69 $Y2=0.755
cc_100 N_A_c_104_n N_Y_c_217_n 0.00182852f $X=0.905 $Y=1.22 $X2=0.69 $Y2=0.755
cc_101 N_A_c_131_n N_Y_c_217_n 0.00109947f $X=0.535 $Y=1.825 $X2=0.69 $Y2=0.755
cc_102 N_A_c_132_n N_Y_c_239_n 0.00183112f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.48
cc_103 N_A_c_103_n N_Y_c_239_n 0.00869502f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.48
cc_104 N_A_c_137_n N_Y_c_239_n 0.00335296f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.48
cc_105 N_A_c_122_n N_Y_c_239_n 2.38128e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_106 N_A_c_129_n N_Y_c_239_n 0.0226156f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.48
cc_107 N_A_c_131_n N_Y_c_239_n 0.00165526f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.48
cc_108 A N_Y_c_239_n 0.00938699f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.48
cc_109 N_A_c_111_n N_Y_c_221_n 0.00182852f $X=1.335 $Y=1.22 $X2=1.55 $Y2=0.755
cc_110 N_A_c_115_n N_Y_c_221_n 0.00310013f $X=1.69 $Y=1.295 $X2=1.55 $Y2=0.755
cc_111 N_A_c_117_n N_Y_c_221_n 0.00182852f $X=1.765 $Y=1.22 $X2=1.55 $Y2=0.755
cc_112 N_A_c_143_n N_Y_c_242_n 0.00335296f $X=1.335 $Y=2.48 $X2=1.55 $Y2=2.48
cc_113 N_A_c_116_n N_Y_c_242_n 0.0105836f $X=1.69 $Y=2.405 $X2=1.55 $Y2=2.48
cc_114 N_A_c_148_n N_Y_c_242_n 0.00335296f $X=1.765 $Y=2.48 $X2=1.55 $Y2=2.48
cc_115 N_A_c_97_n N_Y_c_225_n 0.00880716f $X=0.475 $Y=1.22 $X2=0.69 $Y2=1.115
cc_116 N_A_c_104_n N_Y_c_225_n 0.00198464f $X=0.905 $Y=1.22 $X2=0.69 $Y2=1.115
cc_117 N_A_c_122_n N_Y_c_225_n 6.32153e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=1.115
cc_118 N_A_c_132_n N_Y_c_245_n 0.00169643f $X=0.475 $Y=2.48 $X2=0.69 $Y2=2.365
cc_119 N_A_c_103_n N_Y_c_245_n 0.00259868f $X=0.83 $Y=2.405 $X2=0.69 $Y2=2.365
cc_120 N_A_c_137_n N_Y_c_245_n 0.00144225f $X=0.905 $Y=2.48 $X2=0.69 $Y2=2.365
cc_121 N_A_c_122_n N_Y_c_245_n 2.98633e-19 $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.365
cc_122 N_A_c_124_n N_Y_c_245_n 0.00102602f $X=0.475 $Y=2.405 $X2=0.69 $Y2=2.365
cc_123 N_A_c_126_n N_Y_c_245_n 0.00150284f $X=0.905 $Y=2.405 $X2=0.69 $Y2=2.365
cc_124 N_A_c_129_n N_Y_c_245_n 0.0071561f $X=0.32 $Y=2.85 $X2=0.69 $Y2=2.365
cc_125 N_A_c_131_n N_Y_c_245_n 0.00173027f $X=0.535 $Y=1.825 $X2=0.69 $Y2=2.365
cc_126 A N_Y_c_245_n 0.00805971f $X=0.32 $Y=2.845 $X2=0.69 $Y2=2.365
cc_127 N_A_c_97_n Y 0.00150089f $X=0.475 $Y=1.22 $X2=0.76 $Y2=1.72
cc_128 N_A_c_101_n Y 0.00792324f $X=0.475 $Y=2.33 $X2=0.76 $Y2=1.72
cc_129 N_A_c_102_n Y 0.0163225f $X=0.83 $Y=1.295 $X2=0.76 $Y2=1.72
cc_130 N_A_c_103_n Y 0.0038871f $X=0.83 $Y=2.405 $X2=0.76 $Y2=1.72
cc_131 N_A_c_104_n Y 0.00150089f $X=0.905 $Y=1.22 $X2=0.76 $Y2=1.72
cc_132 N_A_c_122_n Y 0.00610708f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_133 N_A_c_123_n Y 0.00675469f $X=0.535 $Y=1.66 $X2=0.76 $Y2=1.72
cc_134 N_A_c_129_n Y 0.0182346f $X=0.32 $Y=2.85 $X2=0.76 $Y2=1.72
cc_135 N_A_c_131_n Y 0.0178517f $X=0.535 $Y=1.825 $X2=0.76 $Y2=1.72
cc_136 N_A_c_104_n N_Y_c_230_n 0.00869047f $X=0.905 $Y=1.22 $X2=1.405 $Y2=1
cc_137 N_A_c_108_n N_Y_c_230_n 0.0022289f $X=1.26 $Y=1.295 $X2=1.405 $Y2=1
cc_138 N_A_c_111_n N_Y_c_230_n 0.00869047f $X=1.335 $Y=1.22 $X2=1.405 $Y2=1
cc_139 N_A_c_137_n N_Y_c_246_n 0.00693713f $X=0.905 $Y=2.48 $X2=1.405 $Y2=2.48
cc_140 N_A_c_110_n N_Y_c_246_n 0.0120397f $X=1.26 $Y=2.405 $X2=1.405 $Y2=2.48
cc_141 N_A_c_143_n N_Y_c_246_n 0.00693713f $X=1.335 $Y=2.48 $X2=1.405 $Y2=2.48
cc_142 N_A_c_126_n N_Y_c_246_n 0.00560085f $X=0.905 $Y=2.405 $X2=1.405 $Y2=2.48
cc_143 N_A_c_128_n N_Y_c_246_n 0.00560085f $X=1.335 $Y=2.405 $X2=1.405 $Y2=2.48
cc_144 N_A_c_111_n N_Y_c_234_n 0.00198464f $X=1.335 $Y=1.22 $X2=1.55 $Y2=1.115
cc_145 N_A_c_117_n N_Y_c_234_n 0.00878106f $X=1.765 $Y=1.22 $X2=1.55 $Y2=1.115
cc_146 N_A_c_111_n N_Y_c_238_n 0.00150089f $X=1.335 $Y=1.22 $X2=1.55 $Y2=2.365
cc_147 N_A_c_143_n N_Y_c_238_n 0.00144225f $X=1.335 $Y=2.48 $X2=1.55 $Y2=2.365
cc_148 N_A_c_115_n N_Y_c_238_n 0.0169795f $X=1.69 $Y=1.295 $X2=1.55 $Y2=2.365
cc_149 N_A_c_116_n N_Y_c_238_n 0.0141541f $X=1.69 $Y=2.405 $X2=1.55 $Y2=2.365
cc_150 N_A_c_117_n N_Y_c_238_n 0.00150089f $X=1.765 $Y=1.22 $X2=1.55 $Y2=2.365
cc_151 N_A_c_148_n N_Y_c_238_n 0.00541616f $X=1.765 $Y=2.48 $X2=1.55 $Y2=2.365
cc_152 N_A_c_128_n N_Y_c_238_n 0.00150284f $X=1.335 $Y=2.405 $X2=1.55 $Y2=2.365
