* File: sky130_osu_sc_18T_ls__or2_1.pxi.spice
* Created: Fri Nov 12 14:19:09 2021
* 
x_PM_SKY130_OSU_SC_18T_LS__OR2_1%GND N_GND_M1003_s N_GND_M1000_d N_GND_M1003_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_LS__OR2_1%GND
x_PM_SKY130_OSU_SC_18T_LS__OR2_1%VDD N_VDD_M1005_d N_VDD_M1002_b N_VDD_c_39_p
+ N_VDD_c_45_p N_VDD_c_52_p VDD N_VDD_c_40_p PM_SKY130_OSU_SC_18T_LS__OR2_1%VDD
x_PM_SKY130_OSU_SC_18T_LS__OR2_1%B N_B_M1003_g N_B_M1002_g N_B_c_66_n N_B_c_67_n
+ B PM_SKY130_OSU_SC_18T_LS__OR2_1%B
x_PM_SKY130_OSU_SC_18T_LS__OR2_1%A N_A_M1000_g N_A_M1005_g N_A_c_94_n N_A_c_95_n
+ A PM_SKY130_OSU_SC_18T_LS__OR2_1%A
x_PM_SKY130_OSU_SC_18T_LS__OR2_1%A_27_617# N_A_27_617#_M1003_d
+ N_A_27_617#_M1002_s N_A_27_617#_M1001_g N_A_27_617#_M1004_g
+ N_A_27_617#_c_137_n N_A_27_617#_c_138_n N_A_27_617#_c_139_n
+ N_A_27_617#_c_151_n N_A_27_617#_c_155_n N_A_27_617#_c_157_n
+ N_A_27_617#_c_140_n N_A_27_617#_c_141_n N_A_27_617#_c_144_n
+ N_A_27_617#_c_146_n PM_SKY130_OSU_SC_18T_LS__OR2_1%A_27_617#
x_PM_SKY130_OSU_SC_18T_LS__OR2_1%Y N_Y_M1001_d N_Y_M1004_d N_Y_c_206_n
+ N_Y_c_209_n Y N_Y_c_211_n N_Y_c_213_n PM_SKY130_OSU_SC_18T_LS__OR2_1%Y
cc_1 N_GND_M1003_b N_B_M1003_g 0.083817f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_B_M1003_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_B_M1003_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_B_M1003_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.075
cc_5 N_GND_M1003_b N_B_M1002_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_6 N_GND_M1003_b N_B_c_66_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.675
cc_7 N_GND_M1003_b N_B_c_67_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.675
cc_8 N_GND_M1003_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.96
cc_9 N_GND_M1003_b N_A_M1000_g 0.0440597f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.075
cc_10 N_GND_c_3_p N_A_M1000_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.075
cc_11 N_GND_c_11_p N_A_M1000_g 0.00354579f $X=1.12 $Y=0.825 $X2=0.905 $Y2=1.075
cc_12 N_GND_c_4_p N_A_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=1.075
cc_13 N_GND_M1003_b N_A_M1005_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_14 N_GND_M1003_b N_A_c_94_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.385
cc_15 N_GND_M1003_b N_A_c_95_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.385
cc_16 N_GND_M1003_b N_A_27_617#_M1001_g 0.0277213f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_c_11_p N_A_27_617#_M1001_g 0.00354579f $X=1.12 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_18 N_GND_c_18_p N_A_27_617#_M1001_g 0.00606474f $X=1.12 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_19 N_GND_c_4_p N_A_27_617#_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335
+ $Y2=1.075
cc_20 N_GND_M1003_b N_A_27_617#_c_137_n 0.0364586f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.1
cc_21 N_GND_M1003_b N_A_27_617#_c_138_n 0.0466273f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.81
cc_22 N_GND_M1003_b N_A_27_617#_c_139_n 0.0076653f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.96
cc_23 N_GND_M1003_b N_A_27_617#_c_140_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.545
cc_24 N_GND_M1003_b N_A_27_617#_c_141_n 0.00710171f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.825
cc_25 N_GND_c_3_p N_A_27_617#_c_141_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.825
cc_26 N_GND_c_4_p N_A_27_617#_c_141_n 0.00475776f $X=1.02 $Y=0.19 $X2=0.69
+ $Y2=0.825
cc_27 N_GND_M1003_b N_A_27_617#_c_144_n 0.0200876f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_28 N_GND_c_11_p N_A_27_617#_c_144_n 0.00702738f $X=1.12 $Y=0.825 $X2=1.43
+ $Y2=1.935
cc_29 N_GND_M1003_b N_A_27_617#_c_146_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.935
cc_30 N_GND_M1003_b N_Y_c_206_n 0.00156053f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_31 N_GND_c_18_p N_Y_c_206_n 0.00757793f $X=1.12 $Y=0.152 $X2=1.55 $Y2=0.825
cc_32 N_GND_c_4_p N_Y_c_206_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.825
cc_33 N_GND_M1003_b N_Y_c_209_n 0.016457f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_34 N_GND_M1003_b Y 0.039938f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_35 N_GND_M1003_b N_Y_c_211_n 0.0121687f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.48
cc_36 N_GND_c_11_p N_Y_c_211_n 0.00125659f $X=1.12 $Y=0.825 $X2=1.55 $Y2=1.48
cc_37 N_GND_M1003_b N_Y_c_213_n 0.0141689f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_38 N_VDD_M1002_b N_B_M1002_g 0.0260091f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_39 N_VDD_c_39_p N_B_M1002_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475 $Y2=4.585
cc_40 N_VDD_c_40_p N_B_M1002_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.475 $Y2=4.585
cc_41 N_VDD_M1002_b N_B_c_67_n 0.00375034f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.675
cc_42 N_VDD_M1002_b B 0.0108395f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.96
cc_43 N_VDD_M1002_b N_A_M1005_g 0.0195137f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_44 N_VDD_c_39_p N_A_M1005_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905 $Y2=4.585
cc_45 N_VDD_c_45_p N_A_M1005_g 0.00354579f $X=1.12 $Y=4.135 $X2=0.905 $Y2=4.585
cc_46 N_VDD_c_40_p N_A_M1005_g 0.00468827f $X=1.02 $Y=6.47 $X2=0.905 $Y2=4.585
cc_47 N_VDD_M1002_b N_A_c_95_n 0.00153494f $X=-0.045 $Y=2.905 $X2=0.95 $Y2=2.385
cc_48 N_VDD_M1005_d A 0.0077995f $X=0.98 $Y=3.085 $X2=0.95 $Y2=3.33
cc_49 N_VDD_c_45_p A 0.00247404f $X=1.12 $Y=4.135 $X2=0.95 $Y2=3.33
cc_50 N_VDD_M1002_b N_A_27_617#_c_139_n 0.0267159f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.96
cc_51 N_VDD_c_45_p N_A_27_617#_c_139_n 0.00354579f $X=1.12 $Y=4.135 $X2=1.352
+ $Y2=2.96
cc_52 N_VDD_c_52_p N_A_27_617#_c_139_n 0.00606474f $X=1.12 $Y=6.507 $X2=1.352
+ $Y2=2.96
cc_53 N_VDD_c_40_p N_A_27_617#_c_139_n 0.00468827f $X=1.02 $Y=6.47 $X2=1.352
+ $Y2=2.96
cc_54 N_VDD_M1002_b N_A_27_617#_c_151_n 0.00156053f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.795
cc_55 N_VDD_c_39_p N_A_27_617#_c_151_n 0.00736239f $X=1.035 $Y=6.507 $X2=0.26
+ $Y2=3.795
cc_56 N_VDD_c_40_p N_A_27_617#_c_151_n 0.00476261f $X=1.02 $Y=6.47 $X2=0.26
+ $Y2=3.795
cc_57 N_VDD_M1002_b N_A_27_617#_c_140_n 0.00106577f $X=-0.045 $Y=2.905 $X2=0.61
+ $Y2=3.545
cc_58 N_VDD_M1002_b N_Y_c_209_n 0.010295f $X=-0.045 $Y=2.905 $X2=1.55 $Y2=2.59
cc_59 N_VDD_c_52_p N_Y_c_209_n 0.00757793f $X=1.12 $Y=6.507 $X2=1.55 $Y2=2.59
cc_60 N_VDD_c_40_p N_Y_c_209_n 0.00476261f $X=1.02 $Y=6.47 $X2=1.55 $Y2=2.59
cc_61 N_B_M1003_g N_A_M1000_g 0.0402111f $X=0.475 $Y=1.075 $X2=0.905 $Y2=1.075
cc_62 N_B_c_66_n N_A_M1005_g 0.154838f $X=0.475 $Y=2.675 $X2=0.905 $Y2=4.585
cc_63 N_B_M1003_g N_A_c_94_n 0.0148656f $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.385
cc_64 N_B_M1003_g N_A_c_95_n 0.00121111f $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.385
cc_65 N_B_M1002_g N_A_27_617#_c_155_n 0.0140282f $X=0.475 $Y=4.585 $X2=0.525
+ $Y2=3.63
cc_66 B N_A_27_617#_c_155_n 0.00520961f $X=0.27 $Y=2.96 $X2=0.525 $Y2=3.63
cc_67 N_B_c_67_n N_A_27_617#_c_157_n 0.00369517f $X=0.27 $Y=2.675 $X2=0.345
+ $Y2=3.63
cc_68 B N_A_27_617#_c_157_n 0.00431991f $X=0.27 $Y=2.96 $X2=0.345 $Y2=3.63
cc_69 N_B_M1003_g N_A_27_617#_c_140_n 0.0231435f $X=0.475 $Y=1.075 $X2=0.61
+ $Y2=3.545
cc_70 N_B_M1002_g N_A_27_617#_c_140_n 0.026563f $X=0.475 $Y=4.585 $X2=0.61
+ $Y2=3.545
cc_71 N_B_c_66_n N_A_27_617#_c_140_n 0.00764878f $X=0.475 $Y=2.675 $X2=0.61
+ $Y2=3.545
cc_72 N_B_c_67_n N_A_27_617#_c_140_n 0.0350086f $X=0.27 $Y=2.675 $X2=0.61
+ $Y2=3.545
cc_73 B N_A_27_617#_c_140_n 0.00758489f $X=0.27 $Y=2.96 $X2=0.61 $Y2=3.545
cc_74 N_B_M1003_g N_A_27_617#_c_141_n 0.00765999f $X=0.475 $Y=1.075 $X2=0.69
+ $Y2=0.825
cc_75 N_B_M1003_g N_A_27_617#_c_146_n 0.0113001f $X=0.475 $Y=1.075 $X2=0.65
+ $Y2=1.935
cc_76 N_A_M1000_g N_A_27_617#_M1001_g 0.030724f $X=0.905 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_77 N_A_M1000_g N_A_27_617#_c_137_n 0.0119161f $X=0.905 $Y=1.075 $X2=1.37
+ $Y2=2.1
cc_78 N_A_M1005_g N_A_27_617#_c_138_n 0.00914307f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.81
cc_79 N_A_c_94_n N_A_27_617#_c_138_n 0.0204279f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.81
cc_80 N_A_c_95_n N_A_27_617#_c_138_n 0.00375034f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.81
cc_81 N_A_M1005_g N_A_27_617#_c_139_n 0.0540618f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.96
cc_82 N_A_c_95_n N_A_27_617#_c_139_n 0.00341181f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.96
cc_83 A N_A_27_617#_c_139_n 0.00374181f $X=0.95 $Y=3.33 $X2=1.352 $Y2=2.96
cc_84 N_A_M1005_g N_A_27_617#_c_155_n 0.00457566f $X=0.905 $Y=4.585 $X2=0.525
+ $Y2=3.63
cc_85 N_A_M1000_g N_A_27_617#_c_140_n 0.00429604f $X=0.905 $Y=1.075 $X2=0.61
+ $Y2=3.545
cc_86 N_A_M1005_g N_A_27_617#_c_140_n 0.00776428f $X=0.905 $Y=4.585 $X2=0.61
+ $Y2=3.545
cc_87 N_A_c_94_n N_A_27_617#_c_140_n 0.0021255f $X=0.95 $Y=2.385 $X2=0.61
+ $Y2=3.545
cc_88 N_A_c_95_n N_A_27_617#_c_140_n 0.0822139f $X=0.95 $Y=2.385 $X2=0.61
+ $Y2=3.545
cc_89 A N_A_27_617#_c_140_n 0.00866797f $X=0.95 $Y=3.33 $X2=0.61 $Y2=3.545
cc_90 N_A_M1000_g N_A_27_617#_c_141_n 0.00765999f $X=0.905 $Y=1.075 $X2=0.69
+ $Y2=0.825
cc_91 N_A_M1000_g N_A_27_617#_c_144_n 0.0163305f $X=0.905 $Y=1.075 $X2=1.43
+ $Y2=1.935
cc_92 N_A_c_94_n N_A_27_617#_c_144_n 0.00276813f $X=0.95 $Y=2.385 $X2=1.43
+ $Y2=1.935
cc_93 N_A_c_95_n N_A_27_617#_c_144_n 0.0114342f $X=0.95 $Y=2.385 $X2=1.43
+ $Y2=1.935
cc_94 A A_110_617# 0.0123256f $X=0.95 $Y=3.33 $X2=0.55 $Y2=3.085
cc_95 N_A_c_95_n N_Y_c_209_n 0.0212254f $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_96 A N_Y_c_209_n 0.00659455f $X=0.95 $Y=3.33 $X2=1.55 $Y2=2.59
cc_97 N_A_M1000_g Y 6.73508e-19 $X=0.905 $Y=1.075 $X2=1.555 $Y2=2.22
cc_98 N_A_c_95_n Y 0.00825539f $X=0.95 $Y=2.385 $X2=1.555 $Y2=2.22
cc_99 N_A_M1000_g N_Y_c_211_n 7.99941e-19 $X=0.905 $Y=1.075 $X2=1.55 $Y2=1.48
cc_100 N_A_c_94_n N_Y_c_213_n 3.65268e-19 $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_101 N_A_c_95_n N_Y_c_213_n 0.00535705f $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_102 N_A_27_617#_c_155_n A_110_617# 0.00613297f $X=0.525 $Y=3.63 $X2=0.55
+ $Y2=3.085
cc_103 N_A_27_617#_c_140_n A_110_617# 0.00377193f $X=0.61 $Y=3.545 $X2=0.55
+ $Y2=3.085
cc_104 N_A_27_617#_M1001_g N_Y_c_206_n 0.0057847f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_105 N_A_27_617#_c_137_n N_Y_c_206_n 0.00168f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=0.825
cc_106 N_A_27_617#_c_144_n N_Y_c_206_n 0.00510008f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_107 N_A_27_617#_c_137_n N_Y_c_209_n 0.00125776f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_108 N_A_27_617#_c_138_n N_Y_c_209_n 0.0115869f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_109 N_A_27_617#_c_139_n N_Y_c_209_n 0.00755607f $X=1.352 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_110 N_A_27_617#_c_144_n N_Y_c_209_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_111 N_A_27_617#_M1001_g Y 0.00406656f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_112 N_A_27_617#_c_137_n Y 0.00704613f $X=1.37 $Y=2.1 $X2=1.555 $Y2=2.22
cc_113 N_A_27_617#_c_138_n Y 0.00892438f $X=1.352 $Y=2.81 $X2=1.555 $Y2=2.22
cc_114 N_A_27_617#_c_144_n Y 0.0151477f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_115 N_A_27_617#_M1001_g N_Y_c_211_n 0.00669813f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.48
cc_116 N_A_27_617#_c_137_n N_Y_c_211_n 0.00154864f $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=1.48
cc_117 N_A_27_617#_c_144_n N_Y_c_211_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.48
cc_118 N_A_27_617#_c_137_n N_Y_c_213_n 4.58687e-19 $X=1.37 $Y=2.1 $X2=1.55
+ $Y2=2.59
cc_119 N_A_27_617#_c_138_n N_Y_c_213_n 0.00721849f $X=1.352 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_120 N_A_27_617#_c_144_n N_Y_c_213_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
