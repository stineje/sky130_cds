* File: sky130_osu_sc_18T_ls__dffs_l.pex.spice
* Created: Fri Nov 12 14:16:14 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%GND 1 2 3 4 5 6 97 99 107 113 115 125
+ 127 137 139 149 151 158 180 182
c192 137 0 1.67294e-19 $X=5.14 $Y=0.825
c193 113 0 3.07193e-19 $X=1.64 $Y=0.825
c194 97 0 1.27355e-19 $X=-0.05 $Y=0
r195 180 182 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=7.815 $Y2=0.152
r196 156 158 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.825
r197 152 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=0.152
+ $X2=6.88 $Y2=0.152
r198 147 172 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.152
r199 147 149 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.88 $Y=0.305
+ $X2=6.88 $Y2=0.825
r200 139 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=0.152
+ $X2=6.88 $Y2=0.152
r201 135 137 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.14 $Y=0.305
+ $X2=5.14 $Y2=0.825
r202 128 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.152
+ $X2=3.39 $Y2=0.152
r203 123 168 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.152
r204 123 125 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=0.305
+ $X2=3.39 $Y2=0.825
r205 115 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.152
+ $X2=3.39 $Y2=0.152
r206 111 113 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.64 $Y=0.305
+ $X2=1.64 $Y2=0.825
r207 109 110 15.8697 $w=3.03e-07 $l=4.2e-07 $layer=LI1_cond $X=1.555 $Y=0.152
+ $X2=1.135 $Y2=0.152
r208 105 107 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.825
r209 97 182 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=0.19
+ $X2=7.815 $Y2=0.19
r210 97 180 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=0.19
+ $X2=0.335 $Y2=0.19
r211 97 156 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r212 97 151 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r213 97 135 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.14 $Y2=0.305
r214 97 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.055 $Y2=0.152
r215 97 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.152
+ $X2=5.225 $Y2=0.152
r216 97 111 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.64 $Y2=0.305
r217 97 109 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.555 $Y2=0.152
r218 97 116 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.152
+ $X2=1.725 $Y2=0.152
r219 97 105 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r220 97 99 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r221 97 110 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r222 97 151 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r223 97 152 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=6.965 $Y2=0.152
r224 97 139 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.795 $Y2=0.152
r225 97 140 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=5.225 $Y2=0.152
r226 97 127 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=4.415 $Y=0.152
+ $X2=5.055 $Y2=0.152
r227 97 128 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=3.475 $Y2=0.152
r228 97 115 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=3.305 $Y2=0.152
r229 97 116 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=1.725 $Y2=0.152
r230 97 99 23.8046 $w=3.03e-07 $l=6.3e-07 $layer=LI1_cond $X=0.335 $Y=0.152
+ $X2=0.965 $Y2=0.152
r231 6 158 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.825
r232 5 149 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.575 $X2=6.88 $Y2=0.825
r233 4 137 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5
+ $Y=0.575 $X2=5.14 $Y2=0.825
r234 3 125 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.575 $X2=3.39 $Y2=0.825
r235 2 113 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.575 $X2=1.64 $Y2=0.825
r236 1 107 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%VDD 1 2 3 4 5 6 7 8 81 85 89 95 103 107
+ 115 119 127 131 137 141 147 151 157 175 178 182
r105 178 182 3.4836 $w=3.05e-07 $l=7.48e-06 $layer=MET1_cond $X=0.335 $Y=6.507
+ $X2=7.815 $Y2=6.507
r106 175 182 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=7.815 $Y=6.47
+ $X2=7.815 $Y2=6.47
r107 164 178 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.335 $Y=6.47
+ $X2=0.335 $Y2=6.47
r108 157 160 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.9 $Y=4.475
+ $X2=7.9 $Y2=5.835
r109 155 175 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=6.507
r110 155 160 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=6.355
+ $X2=7.9 $Y2=5.835
r111 152 173 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.035 $Y=6.507
+ $X2=6.95 $Y2=6.507
r112 152 154 3.7785 $w=3.03e-07 $l=1e-07 $layer=LI1_cond $X=7.035 $Y=6.507
+ $X2=7.135 $Y2=6.507
r113 151 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.9 $Y2=6.507
r114 151 154 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.815 $Y=6.507
+ $X2=7.135 $Y2=6.507
r115 147 150 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.95 $Y=4.815
+ $X2=6.95 $Y2=5.835
r116 145 173 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.95 $Y=6.355
+ $X2=6.95 $Y2=6.507
r117 145 150 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.95 $Y=6.355
+ $X2=6.95 $Y2=5.835
r118 142 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.09 $Y2=6.507
r119 142 144 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.455 $Y2=6.507
r120 141 173 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=6.507
+ $X2=6.95 $Y2=6.507
r121 141 144 15.4919 $w=3.03e-07 $l=4.1e-07 $layer=LI1_cond $X=6.865 $Y=6.507
+ $X2=6.455 $Y2=6.507
r122 137 140 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.09 $Y=4.815
+ $X2=6.09 $Y2=5.835
r123 135 172 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=6.507
r124 135 140 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=5.835
r125 132 171 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.14 $Y2=6.507
r126 132 134 20.7818 $w=3.03e-07 $l=5.5e-07 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.775 $Y2=6.507
r127 131 172 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=6.09 $Y2=6.507
r128 131 134 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=5.775 $Y2=6.507
r129 127 130 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.14 $Y=3.455
+ $X2=5.14 $Y2=5.835
r130 125 171 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.14 $Y=6.355
+ $X2=5.14 $Y2=6.507
r131 125 130 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.14 $Y=6.355
+ $X2=5.14 $Y2=5.835
r132 122 124 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=6.507
+ $X2=4.415 $Y2=6.507
r133 120 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=6.507
+ $X2=3.39 $Y2=6.507
r134 120 122 9.8241 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=3.475 $Y=6.507
+ $X2=3.735 $Y2=6.507
r135 119 171 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=6.507
+ $X2=5.14 $Y2=6.507
r136 119 124 24.1824 $w=3.03e-07 $l=6.4e-07 $layer=LI1_cond $X=5.055 $Y=6.507
+ $X2=4.415 $Y2=6.507
r137 115 118 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=3.39 $Y=3.795
+ $X2=3.39 $Y2=5.835
r138 113 169 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.39 $Y=6.355
+ $X2=3.39 $Y2=6.507
r139 113 118 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=6.355
+ $X2=3.39 $Y2=5.835
r140 110 112 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.375 $Y=6.507
+ $X2=3.055 $Y2=6.507
r141 108 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=6.507
+ $X2=1.64 $Y2=6.507
r142 108 110 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=1.725 $Y=6.507
+ $X2=2.375 $Y2=6.507
r143 107 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=6.507
+ $X2=3.39 $Y2=6.507
r144 107 112 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.305 $Y=6.507
+ $X2=3.055 $Y2=6.507
r145 103 106 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.64 $Y=3.795
+ $X2=1.64 $Y2=5.835
r146 101 168 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.64 $Y=6.355
+ $X2=1.64 $Y2=6.507
r147 101 106 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.64 $Y=6.355
+ $X2=1.64 $Y2=5.835
r148 100 166 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=6.507
+ $X2=1.12 $Y2=6.507
r149 99 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=6.507
+ $X2=1.64 $Y2=6.507
r150 99 100 13.2248 $w=3.03e-07 $l=3.5e-07 $layer=LI1_cond $X=1.555 $Y=6.507
+ $X2=1.205 $Y2=6.507
r151 95 98 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=4.815
+ $X2=1.12 $Y2=5.835
r152 93 166 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=6.507
r153 93 98 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=6.355
+ $X2=1.12 $Y2=5.835
r154 90 164 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r155 90 92 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.015 $Y2=6.507
r156 89 166 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.12 $Y2=6.507
r157 89 92 0.7557 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=1.035 $Y=6.507
+ $X2=1.015 $Y2=6.507
r158 85 88 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=4.815
+ $X2=0.26 $Y2=5.835
r159 83 164 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r160 83 88 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r161 81 175 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=6.355 $X2=7.815 $Y2=6.44
r162 81 154 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=6.355 $X2=7.135 $Y2=6.44
r163 81 144 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=6.355 $X2=6.455 $Y2=6.44
r164 81 134 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=6.355 $X2=5.775 $Y2=6.44
r165 81 171 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=6.355 $X2=5.095 $Y2=6.44
r166 81 124 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=6.355 $X2=4.415 $Y2=6.44
r167 81 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=6.355 $X2=3.735 $Y2=6.44
r168 81 112 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=6.355 $X2=3.055 $Y2=6.44
r169 81 110 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=6.355 $X2=2.375 $Y2=6.44
r170 81 168 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=6.355 $X2=1.695 $Y2=6.44
r171 81 92 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=6.355 $X2=1.015 $Y2=6.44
r172 81 164 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=6.355 $X2=0.335 $Y2=6.44
r173 8 160 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=4.085 $X2=7.9 $Y2=5.835
r174 8 157 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=4.085 $X2=7.9 $Y2=4.475
r175 7 150 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=4.085 $X2=6.95 $Y2=5.835
r176 7 147 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=4.085 $X2=6.95 $Y2=4.815
r177 6 140 300 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=5.965
+ $Y=4.085 $X2=6.09 $Y2=5.835
r178 6 137 300 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=2 $X=5.965
+ $Y=4.085 $X2=6.09 $Y2=4.815
r179 5 130 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5
+ $Y=3.085 $X2=5.14 $Y2=5.835
r180 5 127 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5
+ $Y=3.085 $X2=5.14 $Y2=3.455
r181 4 118 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=3.25 $Y=3.085 $X2=3.39 $Y2=5.835
r182 4 115 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=3.25 $Y=3.085 $X2=3.39 $Y2=3.795
r183 3 106 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=1.515 $Y=3.085 $X2=1.64 $Y2=5.835
r184 3 103 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=1.515 $Y=3.085 $X2=1.64 $Y2=3.795
r185 2 98 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=5.835
r186 2 95 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=4.085 $X2=1.12 $Y2=4.815
r187 1 88 300 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=5.835
r188 1 85 300 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=4.085 $X2=0.26 $Y2=4.815
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%SN 3 7 9 11 14 17 21 25 31 36 37 39 44
r130 37 39 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.465 $Y=1.48
+ $X2=0.32 $Y2=1.48
r131 36 44 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.715 $Y=1.48
+ $X2=6.86 $Y2=1.48
r132 36 37 6.01801 $w=1.7e-07 $l=6.25e-06 $layer=MET1_cond $X=6.715 $Y=1.48
+ $X2=0.465 $Y2=1.48
r133 31 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.86 $Y=1.48
+ $X2=6.86 $Y2=1.48
r134 31 34 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.86 $Y=1.48
+ $X2=6.86 $Y2=1.59
r135 25 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=1.48
+ $X2=0.32 $Y2=1.48
r136 25 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.48
+ $X2=0.32 $Y2=1.85
r137 23 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.59 $X2=6.86 $Y2=1.59
r138 21 23 19.0665 $w=3.16e-07 $l=1.25e-07 $layer=POLY_cond $X=6.735 $Y=1.59
+ $X2=6.86 $Y2=1.59
r139 20 21 10.6772 $w=3.16e-07 $l=7e-08 $layer=POLY_cond $X=6.665 $Y=1.59
+ $X2=6.735 $Y2=1.59
r140 17 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.85 $X2=0.32 $Y2=1.85
r141 17 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.85
+ $X2=0.367 $Y2=2.015
r142 17 18 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.85
+ $X2=0.367 $Y2=1.685
r143 12 21 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.755
+ $X2=6.735 $Y2=1.59
r144 12 14 1707.51 $w=1.5e-07 $l=3.33e-06 $layer=POLY_cond $X=6.735 $Y=1.755
+ $X2=6.735 $Y2=5.085
r145 9 20 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.665 $Y=1.425
+ $X2=6.665 $Y2=1.59
r146 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.665 $Y=1.425
+ $X2=6.665 $Y2=0.945
r147 7 19 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=0.475 $Y=5.085
+ $X2=0.475 $Y2=2.015
r148 3 18 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.475 $Y=0.945
+ $X2=0.475 $Y2=1.685
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%A_152_89# 1 3 11 15 21 26 27 28 29 30 32
+ 35 39 44
c86 44 0 1.71621e-19 $X=2.507 $Y=1.415
c87 27 0 1.29912e-19 $X=2.33 $Y=1.765
r88 43 44 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.507 $Y=1.245
+ $X2=2.507 $Y2=1.415
r89 39 41 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=2.515 $Y=3.455
+ $X2=2.515 $Y2=5.835
r90 37 39 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=2.515 $Y=3.27
+ $X2=2.515 $Y2=3.455
r91 35 43 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=2.515 $Y=0.825
+ $X2=2.515 $Y2=1.245
r92 32 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.415 $Y=1.68
+ $X2=2.415 $Y2=1.415
r93 29 37 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.345 $Y=3.185
+ $X2=2.515 $Y2=3.27
r94 29 30 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.345 $Y=3.185
+ $X2=1.115 $Y2=3.185
r95 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=1.765
+ $X2=2.415 $Y2=1.68
r96 27 28 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.33 $Y=1.765
+ $X2=1.115 $Y2=1.765
r97 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=3.1
+ $X2=1.115 $Y2=3.185
r98 24 26 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.03 $Y=3.1
+ $X2=1.03 $Y2=2.305
r99 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=1.85
+ $X2=1.115 $Y2=1.765
r100 23 26 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.03 $Y=1.85
+ $X2=1.03 $Y2=2.305
r101 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=2.305 $X2=1.03 $Y2=2.305
r102 19 21 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.905 $Y=2.305
+ $X2=1.03 $Y2=2.305
r103 17 19 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.835 $Y=2.305
+ $X2=0.905 $Y2=2.305
r104 13 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.47
+ $X2=0.905 $Y2=2.305
r105 13 15 1340.88 $w=1.5e-07 $l=2.615e-06 $layer=POLY_cond $X=0.905 $Y=2.47
+ $X2=0.905 $Y2=5.085
r106 9 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=2.14
+ $X2=0.835 $Y2=2.305
r107 9 11 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.835 $Y=2.14
+ $X2=0.835 $Y2=0.945
r108 3 41 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=2.29
+ $Y=3.085 $X2=2.515 $Y2=5.835
r109 3 39 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=2.29
+ $Y=3.085 $X2=2.515 $Y2=3.455
r110 1 35 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.575 $X2=2.515 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%D 3 7 10 14 19
c41 19 0 1.41836e-19 $X=1.915 $Y=2.22
c42 10 0 1.12321e-19 $X=1.915 $Y=2.22
r43 14 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.915 $Y=2.22
+ $X2=1.915 $Y2=2.22
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=2.22 $X2=1.915 $Y2=2.22
r45 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=2.22
+ $X2=1.915 $Y2=2.385
r46 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=2.22
+ $X2=1.915 $Y2=2.055
r47 7 12 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=1.855 $Y=4.585
+ $X2=1.855 $Y2=2.385
r48 3 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.855 $Y=1.075
+ $X2=1.855 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%CK 3 7 10 13 17 18 20 23 25 29 30 33 34
+ 37 40 41 44 48 52 54 55 57 63 70 74 75 76 77 84
c218 55 0 6.79641e-20 $X=4.11 $Y=2.59
c219 48 0 1.98654e-19 $X=2.755 $Y=1.85
c220 44 0 1.86602e-19 $X=2.67 $Y=2.59
c221 30 0 1.29912e-19 $X=2.755 $Y=1.685
c222 25 0 1.41836e-19 $X=2.275 $Y=2.765
r223 77 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.65 $Y=2.59
+ $X2=4.505 $Y2=2.59
r224 76 84 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.355 $Y=2.59
+ $X2=5.5 $Y2=2.59
r225 76 77 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=5.355 $Y=2.59
+ $X2=4.65 $Y2=2.59
r226 75 79 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.42 $Y=2.59
+ $X2=2.275 $Y2=2.59
r227 74 82 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.36 $Y=2.59
+ $X2=4.505 $Y2=2.59
r228 74 75 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=4.36 $Y=2.59
+ $X2=2.42 $Y2=2.59
r229 70 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.505 $Y=2.59
+ $X2=4.505 $Y2=2.59
r230 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.505 $Y=2.59
+ $X2=4.505 $Y2=2.765
r231 63 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.275 $Y=2.59
+ $X2=2.275 $Y2=2.59
r232 63 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.275 $Y=2.59
+ $X2=2.275 $Y2=2.765
r233 57 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.5 $Y=2.59 $X2=5.5
+ $Y2=2.59
r234 57 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.5 $Y=2.59
+ $X2=5.5 $Y2=2.765
r235 54 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.59
+ $X2=4.505 $Y2=2.59
r236 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.42 $Y=2.59
+ $X2=4.11 $Y2=2.59
r237 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=2.505
+ $X2=4.11 $Y2=2.59
r238 50 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.025 $Y=2.505
+ $X2=4.025 $Y2=1.85
r239 46 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.755 $Y=2.505
+ $X2=2.755 $Y2=1.85
r240 45 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.59
+ $X2=2.275 $Y2=2.59
r241 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.67 $Y=2.59
+ $X2=2.755 $Y2=2.505
r242 44 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.67 $Y=2.59
+ $X2=2.36 $Y2=2.59
r243 43 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=2.765 $X2=5.5 $Y2=2.765
r244 40 41 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=5.382 $Y=1.685
+ $X2=5.382 $Y2=1.835
r245 37 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=2.765 $X2=4.505 $Y2=2.765
r246 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=2.765
+ $X2=4.505 $Y2=2.93
r247 33 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.85 $X2=4.025 $Y2=1.85
r248 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.85
+ $X2=4.025 $Y2=1.685
r249 29 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.85 $X2=2.755 $Y2=1.85
r250 29 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.85
+ $X2=2.755 $Y2=1.685
r251 25 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=2.765 $X2=2.275 $Y2=2.765
r252 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=2.765
+ $X2=2.275 $Y2=2.93
r253 23 43 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=5.41 $Y=2.6
+ $X2=5.457 $Y2=2.765
r254 23 41 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=5.41 $Y=2.6
+ $X2=5.41 $Y2=1.835
r255 18 43 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=5.355 $Y=2.93
+ $X2=5.457 $Y2=2.765
r256 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.355 $Y=2.93
+ $X2=5.355 $Y2=4.585
r257 17 40 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.355 $Y=1.075
+ $X2=5.355 $Y2=1.685
r258 13 39 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=4.565 $Y=4.585
+ $X2=4.565 $Y2=2.93
r259 10 34 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.965 $Y=1.075
+ $X2=3.965 $Y2=1.685
r260 7 30 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.815 $Y=1.075
+ $X2=2.815 $Y2=1.685
r261 3 27 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.215 $Y=4.585
+ $X2=2.215 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%A_27_115# 1 3 11 15 17 18 21 22 27 31 35
+ 37 38 41 49 54 55 56 61
c127 55 0 1.35571e-19 $X=3.11 $Y=1.85
c128 49 0 1.5821e-19 $X=3.345 $Y=2.765
c129 31 0 6.36774e-20 $X=3.605 $Y=4.585
c130 22 0 1.86602e-19 $X=3.25 $Y=2.765
c131 21 0 6.79641e-20 $X=3.53 $Y=2.765
c132 15 0 6.36774e-20 $X=3.175 $Y=4.585
r133 56 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.85
+ $X2=0.69 $Y2=1.85
r134 55 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.11 $Y=1.85
+ $X2=3.255 $Y2=1.85
r135 55 56 2.19056 $w=1.7e-07 $l=2.275e-06 $layer=MET1_cond $X=3.11 $Y=1.85
+ $X2=0.835 $Y2=1.85
r136 52 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.255 $Y=1.85
+ $X2=3.255 $Y2=1.85
r137 52 54 4.94595 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=3.255 $Y=1.81
+ $X2=3.345 $Y2=1.81
r138 47 54 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=1.935
+ $X2=3.345 $Y2=1.81
r139 47 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.345 $Y=1.935
+ $X2=3.345 $Y2=2.765
r140 43 45 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=4.815
+ $X2=0.69 $Y2=5.835
r141 41 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=1.85
r142 41 43 193.439 $w=1.68e-07 $l=2.965e-06 $layer=LI1_cond $X=0.69 $Y=1.85
+ $X2=0.69 $Y2=4.815
r143 39 41 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.69 $Y=1.165
+ $X2=0.69 $Y2=1.85
r144 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.08
+ $X2=0.69 $Y2=1.165
r145 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.08
+ $X2=0.345 $Y2=1.08
r146 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.995
+ $X2=0.345 $Y2=1.08
r147 33 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.26 $Y=0.995
+ $X2=0.26 $Y2=0.825
r148 29 31 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=3.605 $Y=2.9
+ $X2=3.605 $Y2=4.585
r149 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.605 $Y=1.715
+ $X2=3.605 $Y2=1.075
r150 24 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=2.765 $X2=3.345 $Y2=2.765
r151 22 24 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=2.765
+ $X2=3.345 $Y2=2.765
r152 21 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.53 $Y=2.765
+ $X2=3.605 $Y2=2.9
r153 21 24 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=2.765
+ $X2=3.345 $Y2=2.765
r154 20 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.85 $X2=3.345 $Y2=1.85
r155 18 20 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.25 $Y=1.85
+ $X2=3.345 $Y2=1.85
r156 17 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.53 $Y=1.85
+ $X2=3.605 $Y2=1.715
r157 17 20 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.53 $Y=1.85
+ $X2=3.345 $Y2=1.85
r158 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=2.9
+ $X2=3.25 $Y2=2.765
r159 13 15 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=3.175 $Y=2.9
+ $X2=3.175 $Y2=4.585
r160 9 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.175 $Y=1.715
+ $X2=3.25 $Y2=1.85
r161 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.175 $Y=1.715
+ $X2=3.175 $Y2=1.075
r162 3 45 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=5.835
r163 3 43 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=4.085 $X2=0.69 $Y2=4.815
r164 1 35 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%A_428_89# 1 3 9 11 13 14 15 18 20 24 26
+ 29 32 35 37 38 40 41 43 49 52 55 60 61 64 68
c188 35 0 1.98654e-19 $X=2.335 $Y=1.76
c189 18 0 1.12321e-19 $X=2.815 $Y=4.585
r190 66 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=3.185
+ $X2=5.845 $Y2=3.185
r191 62 64 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.57 $Y=2.25
+ $X2=5.845 $Y2=2.25
r192 60 68 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=3.1
+ $X2=5.845 $Y2=3.185
r193 59 64 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.335
+ $X2=5.845 $Y2=2.25
r194 59 60 47.1364 $w=1.78e-07 $l=7.65e-07 $layer=LI1_cond $X=5.845 $Y=2.335
+ $X2=5.845 $Y2=3.1
r195 55 57 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=5.57 $Y=3.455
+ $X2=5.57 $Y2=5.835
r196 53 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=3.27
+ $X2=5.57 $Y2=3.185
r197 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.57 $Y=3.27
+ $X2=5.57 $Y2=3.455
r198 52 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=2.165
+ $X2=5.57 $Y2=2.25
r199 51 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.935
+ $X2=5.57 $Y2=1.85
r200 51 52 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.57 $Y=1.935
+ $X2=5.57 $Y2=2.165
r201 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.765
+ $X2=5.57 $Y2=1.85
r202 47 49 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.57 $Y=1.765
+ $X2=5.57 $Y2=0.825
r203 43 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=1.85
+ $X2=5.57 $Y2=1.85
r204 43 45 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.485 $Y=1.85
+ $X2=4.505 $Y2=1.85
r205 40 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=1.85 $X2=4.505 $Y2=1.85
r206 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.85
+ $X2=4.505 $Y2=2.015
r207 40 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.85
+ $X2=4.505 $Y2=1.685
r208 33 35 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.215 $Y=1.76
+ $X2=2.335 $Y2=1.76
r209 32 41 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.565 $Y=1.075
+ $X2=4.565 $Y2=1.685
r210 29 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.445 $Y=2.225
+ $X2=4.445 $Y2=2.015
r211 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=2.3
+ $X2=3.965 $Y2=2.3
r212 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.37 $Y=2.3
+ $X2=4.445 $Y2=2.225
r213 26 27 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.37 $Y=2.3
+ $X2=4.04 $Y2=2.3
r214 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.965 $Y=2.375
+ $X2=3.965 $Y2=2.3
r215 22 24 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=3.965 $Y=2.375
+ $X2=3.965 $Y2=4.585
r216 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.89 $Y=2.3
+ $X2=2.815 $Y2=2.3
r217 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.89 $Y=2.3
+ $X2=3.965 $Y2=2.3
r218 20 21 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.89 $Y=2.3 $X2=2.89
+ $Y2=2.3
r219 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.815 $Y=2.375
+ $X2=2.815 $Y2=2.3
r220 16 18 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=2.815 $Y=2.375
+ $X2=2.815 $Y2=4.585
r221 14 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.74 $Y=2.3
+ $X2=2.815 $Y2=2.3
r222 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.74 $Y=2.3
+ $X2=2.41 $Y2=2.3
r223 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.335 $Y=2.225
+ $X2=2.41 $Y2=2.3
r224 12 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.335 $Y=1.835
+ $X2=2.335 $Y2=1.76
r225 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.335 $Y=1.835
+ $X2=2.335 $Y2=2.225
r226 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.215 $Y=1.685
+ $X2=2.215 $Y2=1.76
r227 9 11 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.215 $Y=1.685
+ $X2=2.215 $Y2=1.075
r228 3 57 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5.43
+ $Y=3.085 $X2=5.57 $Y2=5.835
r229 3 55 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5.43
+ $Y=3.085 $X2=5.57 $Y2=3.455
r230 1 49 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.43
+ $Y=0.575 $X2=5.57 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%A_970_89# 1 3 11 15 23 27 30 34 35 38 39
+ 40 42 48 50 51 53 56 62 65 66 67 72
c166 39 0 8.77106e-20 $X=7.66 $Y=2.855
c167 34 0 2.20654e-19 $X=7.57 $Y=2.19
r168 67 69 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.13 $Y=2.19
+ $X2=4.985 $Y2=2.19
r169 66 72 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.425 $Y=2.19
+ $X2=7.57 $Y2=2.19
r170 66 67 2.20982 $w=1.7e-07 $l=2.295e-06 $layer=MET1_cond $X=7.425 $Y=2.19
+ $X2=5.13 $Y2=2.19
r171 62 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.57 $Y=2.19
+ $X2=7.57 $Y2=2.19
r172 60 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=2.19
+ $X2=6.52 $Y2=2.19
r173 60 62 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=6.605 $Y=2.19
+ $X2=7.57 $Y2=2.19
r174 56 58 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.52 $Y=4.815
+ $X2=6.52 $Y2=5.835
r175 54 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.275
+ $X2=6.52 $Y2=2.19
r176 54 56 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=6.52 $Y=2.275
+ $X2=6.52 $Y2=4.815
r177 53 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.105
+ $X2=6.52 $Y2=2.19
r178 52 53 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.52 $Y=1.165
+ $X2=6.52 $Y2=2.105
r179 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.435 $Y=1.08
+ $X2=6.52 $Y2=1.165
r180 50 51 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.435 $Y=1.08
+ $X2=6.175 $Y2=1.08
r181 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.09 $Y=0.995
+ $X2=6.175 $Y2=1.08
r182 46 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.09 $Y=0.995
+ $X2=6.09 $Y2=0.825
r183 42 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.985 $Y=2.19
+ $X2=4.985 $Y2=2.19
r184 39 40 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=2.855
+ $X2=7.66 $Y2=3.005
r185 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=1.65 $X2=7.66
+ $Y2=1.8
r186 36 39 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.635 $Y=2.355
+ $X2=7.635 $Y2=2.855
r187 35 38 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.635 $Y=2.025
+ $X2=7.635 $Y2=1.8
r188 34 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=2.19 $X2=7.57 $Y2=2.19
r189 34 36 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=2.19
+ $X2=7.572 $Y2=2.355
r190 34 35 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.572 $Y=2.19
+ $X2=7.572 $Y2=2.025
r191 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=2.19 $X2=4.985 $Y2=2.19
r192 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=2.19
+ $X2=4.985 $Y2=2.355
r193 30 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=2.19
+ $X2=4.985 $Y2=2.025
r194 27 40 1066.55 $w=1.5e-07 $l=2.08e-06 $layer=POLY_cond $X=7.685 $Y=5.085
+ $X2=7.685 $Y2=3.005
r195 23 37 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=7.685 $Y=0.945
+ $X2=7.685 $Y2=1.65
r196 15 32 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=4.925 $Y=4.585
+ $X2=4.925 $Y2=2.355
r197 11 31 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.925 $Y=1.075
+ $X2=4.925 $Y2=2.025
r198 3 58 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=4.085 $X2=6.52 $Y2=5.835
r199 3 56 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=4.085 $X2=6.52 $Y2=4.815
r200 1 48 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=5.965
+ $Y=0.575 $X2=6.09 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%A_808_115# 1 3 11 15 20 25 26 27 28 29
+ 32 36 41 45 46 51
c128 46 0 1.5821e-19 $X=3.83 $Y=1.85
c129 26 0 1.67294e-19 $X=4.095 $Y=1.43
c130 25 0 1.57671e-19 $X=3.685 $Y=1.85
r131 46 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.83 $Y=1.85
+ $X2=3.685 $Y2=1.85
r132 45 51 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.955 $Y=1.85
+ $X2=6.1 $Y2=1.85
r133 45 46 2.04612 $w=1.7e-07 $l=2.125e-06 $layer=MET1_cond $X=5.955 $Y=1.85
+ $X2=3.83 $Y2=1.85
r134 41 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.1 $Y=1.85 $X2=6.1
+ $Y2=1.85
r135 36 38 69.1466 $w=3.38e-07 $l=2.04e-06 $layer=LI1_cond $X=4.265 $Y=3.795
+ $X2=4.265 $Y2=5.835
r136 34 36 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=4.265 $Y=3.27
+ $X2=4.265 $Y2=3.795
r137 30 32 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=4.265 $Y=1.345
+ $X2=4.265 $Y2=0.825
r138 28 34 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=3.185
+ $X2=4.265 $Y2=3.27
r139 28 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=3.185
+ $X2=3.77 $Y2=3.185
r140 26 30 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.095 $Y=1.43
+ $X2=4.265 $Y2=1.345
r141 26 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.095 $Y=1.43
+ $X2=3.77 $Y2=1.43
r142 25 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.685 $Y=1.85
+ $X2=3.685 $Y2=1.85
r143 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=3.1
+ $X2=3.77 $Y2=3.185
r144 23 25 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.685 $Y=3.1
+ $X2=3.685 $Y2=1.85
r145 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=1.515
+ $X2=3.77 $Y2=1.43
r146 22 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.685 $Y=1.515
+ $X2=3.685 $Y2=1.85
r147 18 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.1
+ $Y=1.85 $X2=6.1 $Y2=1.85
r148 18 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.1 $Y=1.85
+ $X2=6.305 $Y2=1.85
r149 13 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=2.015
+ $X2=6.305 $Y2=1.85
r150 13 15 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=6.305 $Y=2.015
+ $X2=6.305 $Y2=5.085
r151 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.685
+ $X2=6.305 $Y2=1.85
r152 9 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.305 $Y=1.685
+ $X2=6.305 $Y2=0.945
r153 3 38 171.429 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=3 $X=4.04
+ $Y=3.085 $X2=4.265 $Y2=5.835
r154 3 36 171.429 $w=1.7e-07 $l=8.1477e-07 $layer=licon1_PDIFF $count=3 $X=4.04
+ $Y=3.085 $X2=4.265 $Y2=3.795
r155 1 32 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=4.04
+ $Y=0.575 $X2=4.265 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c83 44 0 8.77106e-20 $X=7.475 $Y=2.96
c84 35 0 9.99996e-20 $X=7.97 $Y=2.765
c85 33 0 1.20654e-19 $X=7.97 $Y=1.85
r86 42 44 0.00294811 $w=2.12e-07 $l=5e-09 $layer=MET1_cond $X=7.47 $Y=2.96
+ $X2=7.475 $Y2=2.96
r87 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.055 $Y=2.68
+ $X2=8.055 $Y2=2.395
r88 37 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.055 $Y=1.935
+ $X2=8.055 $Y2=2.395
r89 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=2.765
+ $X2=8.055 $Y2=2.68
r90 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=2.765
+ $X2=7.555 $Y2=2.765
r91 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=1.85
+ $X2=8.055 $Y2=1.935
r92 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=1.85
+ $X2=7.555 $Y2=1.85
r93 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.47 $Y=4.475
+ $X2=7.47 $Y2=5.835
r94 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.47 $Y=2.96
+ $X2=7.47 $Y2=2.96
r95 27 29 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=7.47 $Y=2.96
+ $X2=7.47 $Y2=4.475
r96 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=2.85
+ $X2=7.555 $Y2=2.765
r97 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.47 $Y=2.85
+ $X2=7.47 $Y2=2.96
r98 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.47 $Y=1.765
+ $X2=7.555 $Y2=1.85
r99 21 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=7.47 $Y=1.765
+ $X2=7.47 $Y2=0.825
r100 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=2.395 $X2=8.055 $Y2=2.395
r101 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.395
+ $X2=8.055 $Y2=2.56
r102 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.395
+ $X2=8.055 $Y2=2.23
r103 15 20 1294.73 $w=1.5e-07 $l=2.525e-06 $layer=POLY_cond $X=8.115 $Y=5.085
+ $X2=8.115 $Y2=2.56
r104 11 19 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=8.115 $Y=0.945
+ $X2=8.115 $Y2=2.23
r105 3 31 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=4.085 $X2=7.47 $Y2=5.835
r106 3 29 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=4.085 $X2=7.47 $Y2=4.475
r107 1 23 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.575 $X2=7.47 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__DFFS_L%Q 1 3 11 15 20 23 27 30
r22 27 28 6.40639 $w=2.19e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=3.287
+ $X2=8.445 $Y2=3.287
r23 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.325 $Y=3.33
+ $X2=8.325 $Y2=3.33
r24 26 27 0.278539 $w=2.19e-07 $l=5e-09 $layer=LI1_cond $X=8.325 $Y=3.287
+ $X2=8.33 $Y2=3.287
r25 21 23 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=1.515
+ $X2=8.445 $Y2=1.515
r26 20 28 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.445 $Y=3.16
+ $X2=8.445 $Y2=3.287
r27 19 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=1.6
+ $X2=8.445 $Y2=1.515
r28 19 20 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=8.445 $Y=1.6
+ $X2=8.445 $Y2=3.16
r29 15 17 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=8.33 $Y=4.475
+ $X2=8.33 $Y2=5.835
r30 13 27 2.22295 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.33 $Y=3.415
+ $X2=8.33 $Y2=3.287
r31 13 15 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=8.33 $Y=3.415
+ $X2=8.33 $Y2=4.475
r32 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=1.43 $X2=8.33
+ $Y2=1.515
r33 9 11 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.33 $Y=1.43
+ $X2=8.33 $Y2=0.825
r34 3 17 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=4.085 $X2=8.33 $Y2=5.835
r35 3 15 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=4.085 $X2=8.33 $Y2=4.475
r36 1 11 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.575 $X2=8.33 $Y2=0.825
.ends

