* File: sky130_osu_sc_15T_hs__oai21_l.pxi.spice
* Created: Fri Nov 12 14:32:14 2021
* 
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%GND N_GND_M1004_d N_GND_M1004_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_15T_HS__OAI21_L%GND
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%VDD N_VDD_M1002_d N_VDD_M1005_b N_VDD_c_43_p
+ N_VDD_c_49_p N_VDD_c_55_p VDD N_VDD_c_44_p
+ PM_SKY130_OSU_SC_15T_HS__OAI21_L%VDD
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%A0 N_A0_c_68_n N_A0_M1004_g N_A0_M1005_g
+ N_A0_c_72_n N_A0_c_73_n N_A0_c_74_n N_A0_c_75_n A0
+ PM_SKY130_OSU_SC_15T_HS__OAI21_L%A0
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%A1 N_A1_M1002_g N_A1_M1000_g N_A1_c_110_n
+ N_A1_c_111_n N_A1_c_112_n A1 PM_SKY130_OSU_SC_15T_HS__OAI21_L%A1
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%B0 N_B0_M1003_g N_B0_M1001_g N_B0_c_164_n
+ N_B0_c_165_n N_B0_c_166_n N_B0_c_167_n N_B0_c_168_n N_B0_c_169_n B0
+ PM_SKY130_OSU_SC_15T_HS__OAI21_L%B0
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%Y N_Y_M1001_d N_Y_M1005_s N_Y_M1003_d
+ N_Y_c_224_n N_Y_c_227_n N_Y_c_240_n N_Y_c_218_n N_Y_c_231_n N_Y_c_219_n
+ N_Y_c_234_n Y N_Y_c_222_n N_Y_c_223_n PM_SKY130_OSU_SC_15T_HS__OAI21_L%Y
x_PM_SKY130_OSU_SC_15T_HS__OAI21_L%A_27_115# N_A_27_115#_M1004_s
+ N_A_27_115#_M1000_d N_A_27_115#_c_280_n N_A_27_115#_c_283_n
+ N_A_27_115#_c_286_n N_A_27_115#_c_287_n
+ PM_SKY130_OSU_SC_15T_HS__OAI21_L%A_27_115#
cc_1 N_GND_M1004_b N_A0_c_68_n 0.0239294f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.34
cc_2 N_GND_c_2_p N_A0_c_68_n 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=1.34
cc_3 N_GND_c_3_p N_A0_c_68_n 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=1.34
cc_4 N_GND_c_4_p N_A0_c_68_n 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=1.34
cc_5 N_GND_M1004_b N_A0_c_72_n 0.0341998f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.465
cc_6 N_GND_M1004_b N_A0_c_73_n 0.0342885f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.5
cc_7 N_GND_M1004_b N_A0_c_74_n 0.0620905f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.335
cc_8 N_GND_M1004_b N_A0_c_75_n 0.0028102f $X=-0.045 $Y=0 $X2=0.415 $Y2=2.5
cc_9 N_GND_M1004_b N_A1_M1002_g 0.0270518f $X=-0.045 $Y=0 $X2=0.835 $Y2=3.825
cc_10 N_GND_M1004_b N_A1_M1000_g 0.0502927f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.895
cc_11 N_GND_c_3_p N_A1_M1000_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905 $Y2=0.895
cc_12 N_GND_c_4_p N_A1_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=0.895
cc_13 N_GND_M1004_b N_A1_c_110_n 0.0317916f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.96
cc_14 N_GND_M1004_b N_A1_c_111_n 0.00507239f $X=-0.045 $Y=0 $X2=0.845 $Y2=1.96
cc_15 N_GND_M1004_b N_A1_c_112_n 8.57225e-19 $X=-0.045 $Y=0 $X2=0.895 $Y2=2.7
cc_16 N_GND_M1004_b A1 0.00292188f $X=-0.045 $Y=0 $X2=0.895 $Y2=2.7
cc_17 N_GND_M1004_b N_B0_M1003_g 0.0488857f $X=-0.045 $Y=0 $X2=1.325 $Y2=4.195
cc_18 N_GND_M1004_b N_B0_M1001_g 0.0301537f $X=-0.045 $Y=0 $X2=1.335 $Y2=0.895
cc_19 N_GND_c_4_p N_B0_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=1.335 $Y2=0.895
cc_20 N_GND_M1004_b N_B0_c_164_n 0.0152666f $X=-0.045 $Y=0 $X2=1.395 $Y2=1.49
cc_21 N_GND_M1004_b N_B0_c_165_n 0.0155448f $X=-0.045 $Y=0 $X2=1.395 $Y2=1.62
cc_22 N_GND_M1004_b N_B0_c_166_n 0.0108952f $X=-0.045 $Y=0 $X2=1.39 $Y2=1.785
cc_23 N_GND_M1004_b N_B0_c_167_n 0.00586489f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.33
cc_24 N_GND_M1004_b N_B0_c_168_n 0.00505195f $X=-0.045 $Y=0 $X2=1.285 $Y2=1.62
cc_25 N_GND_M1004_b N_B0_c_169_n 0.00240282f $X=-0.045 $Y=0 $X2=1.395 $Y2=1.62
cc_26 N_GND_M1004_b B0 0.0119375f $X=-0.045 $Y=0 $X2=1.2 $Y2=2.33
cc_27 N_GND_M1004_b N_Y_c_218_n 0.0317947f $X=-0.045 $Y=0 $X2=1.54 $Y2=1.96
cc_28 N_GND_M1004_b N_Y_c_219_n 0.012848f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.86
cc_29 N_GND_c_4_p N_Y_c_219_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.55 $Y2=0.86
cc_30 N_GND_M1004_b Y 0.0139051f $X=-0.045 $Y=0 $X2=1.54 $Y2=1.96
cc_31 N_GND_M1004_b N_Y_c_222_n 0.019044f $X=-0.045 $Y=0 $X2=1.54 $Y2=1.845
cc_32 N_GND_M1004_b N_Y_c_223_n 0.0105874f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.22
cc_33 N_GND_M1004_b N_A_27_115#_c_280_n 0.0015601f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.865
cc_34 N_GND_c_2_p N_A_27_115#_c_280_n 0.00735421f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.865
cc_35 N_GND_c_4_p N_A_27_115#_c_280_n 0.00476028f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.865
cc_36 N_GND_M1004_d N_A_27_115#_c_283_n 0.00176461f $X=0.55 $Y=0.575 $X2=1.035
+ $Y2=1.16
cc_37 N_GND_M1004_b N_A_27_115#_c_283_n 0.0125622f $X=-0.045 $Y=0 $X2=1.035
+ $Y2=1.16
cc_38 N_GND_c_3_p N_A_27_115#_c_283_n 0.0135055f $X=0.69 $Y=0.74 $X2=1.035
+ $Y2=1.16
cc_39 N_GND_M1004_b N_A_27_115#_c_286_n 0.00619673f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.16
cc_40 N_GND_M1004_b N_A_27_115#_c_287_n 0.00888269f $X=-0.045 $Y=0 $X2=1.12
+ $Y2=0.865
cc_41 N_GND_c_4_p N_A_27_115#_c_287_n 0.00475544f $X=1.02 $Y=0.19 $X2=1.12
+ $Y2=0.865
cc_42 N_VDD_M1005_b N_A0_M1005_g 0.0241999f $X=-0.045 $Y=2.645 $X2=0.475
+ $Y2=3.825
cc_43 N_VDD_c_43_p N_A0_M1005_g 0.00496961f $X=0.965 $Y=5.397 $X2=0.475
+ $Y2=3.825
cc_44 N_VDD_c_44_p N_A0_M1005_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.475 $Y2=3.825
cc_45 N_VDD_M1005_b N_A0_c_73_n 0.00574563f $X=-0.045 $Y=2.645 $X2=0.415 $Y2=2.5
cc_46 N_VDD_M1005_b N_A0_c_75_n 0.00549657f $X=-0.045 $Y=2.645 $X2=0.415 $Y2=2.5
cc_47 N_VDD_M1005_b N_A1_M1002_g 0.0189209f $X=-0.045 $Y=2.645 $X2=0.835
+ $Y2=3.825
cc_48 N_VDD_c_43_p N_A1_M1002_g 0.00496961f $X=0.965 $Y=5.397 $X2=0.835
+ $Y2=3.825
cc_49 N_VDD_c_49_p N_A1_M1002_g 0.00383116f $X=1.05 $Y=4.225 $X2=0.835 $Y2=3.825
cc_50 N_VDD_c_44_p N_A1_M1002_g 0.00429146f $X=1.02 $Y=5.36 $X2=0.835 $Y2=3.825
cc_51 N_VDD_M1005_b N_A1_c_112_n 0.00163533f $X=-0.045 $Y=2.645 $X2=0.895
+ $Y2=2.7
cc_52 N_VDD_M1005_b A1 0.00594612f $X=-0.045 $Y=2.645 $X2=0.895 $Y2=2.7
cc_53 N_VDD_M1005_b N_B0_M1003_g 0.069243f $X=-0.045 $Y=2.645 $X2=1.325
+ $Y2=4.195
cc_54 N_VDD_c_49_p N_B0_M1003_g 0.010481f $X=1.05 $Y=4.225 $X2=1.325 $Y2=4.195
cc_55 N_VDD_c_55_p N_B0_M1003_g 0.00496961f $X=1.02 $Y=5.36 $X2=1.325 $Y2=4.195
cc_56 N_VDD_c_44_p N_B0_M1003_g 0.00429146f $X=1.02 $Y=5.36 $X2=1.325 $Y2=4.195
cc_57 N_VDD_M1005_b N_Y_c_224_n 0.00199838f $X=-0.045 $Y=2.645 $X2=0.26
+ $Y2=3.885
cc_58 N_VDD_c_43_p N_Y_c_224_n 0.00452684f $X=0.965 $Y=5.397 $X2=0.26 $Y2=3.885
cc_59 N_VDD_c_44_p N_Y_c_224_n 0.00435496f $X=1.02 $Y=5.36 $X2=0.26 $Y2=3.885
cc_60 N_VDD_M1002_d N_Y_c_227_n 0.00888984f $X=0.91 $Y=2.825 $X2=1.455 $Y2=3.41
cc_61 N_VDD_M1005_b N_Y_c_227_n 0.00886322f $X=-0.045 $Y=2.645 $X2=1.455
+ $Y2=3.41
cc_62 N_VDD_c_49_p N_Y_c_227_n 0.00639099f $X=1.05 $Y=4.225 $X2=1.455 $Y2=3.41
cc_63 N_VDD_M1005_b N_Y_c_218_n 0.032421f $X=-0.045 $Y=2.645 $X2=1.54 $Y2=1.96
cc_64 N_VDD_M1005_b N_Y_c_231_n 0.00509863f $X=-0.045 $Y=2.645 $X2=1.54
+ $Y2=4.225
cc_65 N_VDD_c_55_p N_Y_c_231_n 0.00477009f $X=1.02 $Y=5.36 $X2=1.54 $Y2=4.225
cc_66 N_VDD_c_44_p N_Y_c_231_n 0.00435496f $X=1.02 $Y=5.36 $X2=1.54 $Y2=4.225
cc_67 N_VDD_M1005_b N_Y_c_234_n 0.00720662f $X=-0.045 $Y=2.645 $X2=1.54 $Y2=3.41
cc_68 N_A0_c_73_n N_A1_M1002_g 0.159152f $X=0.415 $Y=2.5 $X2=0.835 $Y2=3.825
cc_69 N_A0_c_74_n N_A1_M1002_g 0.00894734f $X=0.415 $Y=2.335 $X2=0.835 $Y2=3.825
cc_70 N_A0_c_75_n N_A1_M1002_g 0.00413298f $X=0.415 $Y=2.5 $X2=0.835 $Y2=3.825
cc_71 A0 N_A1_M1002_g 0.00376364f $X=0.415 $Y=3.07 $X2=0.835 $Y2=3.825
cc_72 N_A0_c_68_n N_A1_M1000_g 0.0359415f $X=0.475 $Y=1.34 $X2=0.905 $Y2=0.895
cc_73 N_A0_c_74_n N_A1_M1000_g 0.00745632f $X=0.415 $Y=2.335 $X2=0.905 $Y2=0.895
cc_74 N_A0_c_74_n N_A1_c_110_n 0.014675f $X=0.415 $Y=2.335 $X2=0.845 $Y2=1.96
cc_75 N_A0_c_73_n N_A1_c_111_n 8.44103e-19 $X=0.415 $Y=2.5 $X2=0.845 $Y2=1.96
cc_76 N_A0_c_74_n N_A1_c_111_n 0.00346793f $X=0.415 $Y=2.335 $X2=0.845 $Y2=1.96
cc_77 N_A0_c_75_n N_A1_c_111_n 0.0189532f $X=0.415 $Y=2.5 $X2=0.845 $Y2=1.96
cc_78 N_A0_M1005_g N_A1_c_112_n 8.44103e-19 $X=0.475 $Y=3.825 $X2=0.895 $Y2=2.7
cc_79 N_A0_c_73_n A1 0.00357623f $X=0.415 $Y=2.5 $X2=0.895 $Y2=2.7
cc_80 N_A0_c_75_n A1 0.00685942f $X=0.415 $Y=2.5 $X2=0.895 $Y2=2.7
cc_81 N_A0_c_75_n N_Y_M1005_s 0.00842425f $X=0.415 $Y=2.5 $X2=0.135 $Y2=2.825
cc_82 A0 N_Y_M1005_s 0.0119025f $X=0.415 $Y=3.07 $X2=0.135 $Y2=2.825
cc_83 N_A0_M1005_g N_Y_c_227_n 0.0157489f $X=0.475 $Y=3.825 $X2=1.455 $Y2=3.41
cc_84 N_A0_c_75_n N_Y_c_227_n 0.0069936f $X=0.415 $Y=2.5 $X2=1.455 $Y2=3.41
cc_85 A0 N_Y_c_227_n 0.0116431f $X=0.415 $Y=3.07 $X2=1.455 $Y2=3.41
cc_86 N_A0_c_73_n N_Y_c_240_n 0.00152768f $X=0.415 $Y=2.5 $X2=0.345 $Y2=3.41
cc_87 N_A0_c_75_n N_Y_c_240_n 9.01113e-19 $X=0.415 $Y=2.5 $X2=0.345 $Y2=3.41
cc_88 A0 N_Y_c_240_n 0.00385855f $X=0.415 $Y=3.07 $X2=0.345 $Y2=3.41
cc_89 A0 A_110_565# 0.0100173f $X=0.415 $Y=3.07 $X2=0.55 $Y2=2.825
cc_90 N_A0_c_68_n N_A_27_115#_c_283_n 0.0200828f $X=0.475 $Y=1.34 $X2=1.035
+ $Y2=1.16
cc_91 N_A0_c_72_n N_A_27_115#_c_283_n 0.00245797f $X=0.475 $Y=1.465 $X2=1.035
+ $Y2=1.16
cc_92 N_A0_c_72_n N_A_27_115#_c_286_n 0.00338493f $X=0.475 $Y=1.465 $X2=0.345
+ $Y2=1.16
cc_93 N_A1_M1002_g N_B0_M1003_g 0.0838551f $X=0.835 $Y=3.825 $X2=1.325 $Y2=4.195
cc_94 N_A1_c_110_n N_B0_M1003_g 0.014032f $X=0.845 $Y=1.96 $X2=1.325 $Y2=4.195
cc_95 N_A1_c_111_n N_B0_M1003_g 0.00248808f $X=0.845 $Y=1.96 $X2=1.325 $Y2=4.195
cc_96 N_A1_c_112_n N_B0_M1003_g 0.00113925f $X=0.895 $Y=2.7 $X2=1.325 $Y2=4.195
cc_97 A1 N_B0_M1003_g 0.00395308f $X=0.895 $Y=2.7 $X2=1.325 $Y2=4.195
cc_98 N_A1_M1000_g N_B0_M1001_g 0.0379553f $X=0.905 $Y=0.895 $X2=1.335 $Y2=0.895
cc_99 N_A1_M1000_g N_B0_c_166_n 0.00505587f $X=0.905 $Y=0.895 $X2=1.39 $Y2=1.785
cc_100 N_A1_M1002_g N_B0_c_167_n 9.28322e-19 $X=0.835 $Y=3.825 $X2=1.2 $Y2=2.33
cc_101 N_A1_M1000_g N_B0_c_167_n 0.00209141f $X=0.905 $Y=0.895 $X2=1.2 $Y2=2.33
cc_102 N_A1_c_110_n N_B0_c_167_n 0.00180004f $X=0.845 $Y=1.96 $X2=1.2 $Y2=2.33
cc_103 N_A1_c_111_n N_B0_c_167_n 0.0395776f $X=0.845 $Y=1.96 $X2=1.2 $Y2=2.33
cc_104 A1 N_B0_c_167_n 2.28089e-19 $X=0.895 $Y=2.7 $X2=1.2 $Y2=2.33
cc_105 N_A1_M1000_g N_B0_c_168_n 0.00444244f $X=0.905 $Y=0.895 $X2=1.285
+ $Y2=1.62
cc_106 N_A1_c_110_n B0 0.00173697f $X=0.845 $Y=1.96 $X2=1.2 $Y2=2.33
cc_107 N_A1_c_111_n B0 0.00816163f $X=0.845 $Y=1.96 $X2=1.2 $Y2=2.33
cc_108 N_A1_c_112_n B0 2.4196e-19 $X=0.895 $Y=2.7 $X2=1.2 $Y2=2.33
cc_109 A1 B0 0.0191116f $X=0.895 $Y=2.7 $X2=1.2 $Y2=2.33
cc_110 N_A1_M1002_g N_Y_c_227_n 0.0165071f $X=0.835 $Y=3.825 $X2=1.455 $Y2=3.41
cc_111 N_A1_c_112_n N_Y_c_227_n 0.00294448f $X=0.895 $Y=2.7 $X2=1.455 $Y2=3.41
cc_112 A1 N_Y_c_227_n 0.0102328f $X=0.895 $Y=2.7 $X2=1.455 $Y2=3.41
cc_113 N_A1_c_111_n N_Y_c_218_n 0.00577978f $X=0.845 $Y=1.96 $X2=1.54 $Y2=1.96
cc_114 N_A1_c_112_n N_Y_c_218_n 0.00365175f $X=0.895 $Y=2.7 $X2=1.54 $Y2=1.96
cc_115 A1 N_Y_c_218_n 0.00695805f $X=0.895 $Y=2.7 $X2=1.54 $Y2=1.96
cc_116 N_A1_M1000_g N_Y_c_222_n 7.34237e-19 $X=0.905 $Y=0.895 $X2=1.54 $Y2=1.845
cc_117 N_A1_M1000_g N_Y_c_223_n 4.01461e-19 $X=0.905 $Y=0.895 $X2=1.55 $Y2=1.22
cc_118 N_A1_M1000_g N_A_27_115#_c_283_n 0.0170892f $X=0.905 $Y=0.895 $X2=1.035
+ $Y2=1.16
cc_119 N_A1_c_110_n N_A_27_115#_c_283_n 0.00300229f $X=0.845 $Y=1.96 $X2=1.035
+ $Y2=1.16
cc_120 N_A1_c_111_n N_A_27_115#_c_283_n 0.00544104f $X=0.845 $Y=1.96 $X2=1.035
+ $Y2=1.16
cc_121 N_B0_M1003_g N_Y_c_227_n 0.0210988f $X=1.325 $Y=4.195 $X2=1.455 $Y2=3.41
cc_122 N_B0_M1003_g N_Y_c_218_n 0.0418701f $X=1.325 $Y=4.195 $X2=1.54 $Y2=1.96
cc_123 N_B0_c_166_n N_Y_c_218_n 0.00154865f $X=1.39 $Y=1.785 $X2=1.54 $Y2=1.96
cc_124 N_B0_c_167_n N_Y_c_218_n 0.0348659f $X=1.2 $Y=2.33 $X2=1.54 $Y2=1.96
cc_125 N_B0_c_169_n N_Y_c_218_n 0.00728781f $X=1.395 $Y=1.62 $X2=1.54 $Y2=1.96
cc_126 B0 N_Y_c_218_n 0.00659213f $X=1.2 $Y=2.33 $X2=1.54 $Y2=1.96
cc_127 N_B0_M1003_g N_Y_c_231_n 0.0128297f $X=1.325 $Y=4.195 $X2=1.54 $Y2=4.225
cc_128 N_B0_M1001_g N_Y_c_219_n 0.00727144f $X=1.335 $Y=0.895 $X2=1.55 $Y2=0.86
cc_129 N_B0_c_164_n N_Y_c_219_n 0.00145376f $X=1.395 $Y=1.49 $X2=1.55 $Y2=0.86
cc_130 N_B0_c_169_n N_Y_c_219_n 0.00486612f $X=1.395 $Y=1.62 $X2=1.55 $Y2=0.86
cc_131 N_B0_M1003_g Y 0.00488821f $X=1.325 $Y=4.195 $X2=1.54 $Y2=1.96
cc_132 N_B0_c_166_n Y 0.00140404f $X=1.39 $Y=1.785 $X2=1.54 $Y2=1.96
cc_133 N_B0_c_167_n Y 0.00656407f $X=1.2 $Y=2.33 $X2=1.54 $Y2=1.96
cc_134 N_B0_c_169_n Y 0.00199558f $X=1.395 $Y=1.62 $X2=1.54 $Y2=1.96
cc_135 N_B0_M1003_g N_Y_c_222_n 0.00137073f $X=1.325 $Y=4.195 $X2=1.54 $Y2=1.845
cc_136 N_B0_M1001_g N_Y_c_222_n 4.4405e-19 $X=1.335 $Y=0.895 $X2=1.54 $Y2=1.845
cc_137 N_B0_c_164_n N_Y_c_222_n 0.0045285f $X=1.395 $Y=1.49 $X2=1.54 $Y2=1.845
cc_138 N_B0_c_165_n N_Y_c_222_n 0.00122529f $X=1.395 $Y=1.62 $X2=1.54 $Y2=1.845
cc_139 N_B0_c_166_n N_Y_c_222_n 0.00223575f $X=1.39 $Y=1.785 $X2=1.54 $Y2=1.845
cc_140 N_B0_c_167_n N_Y_c_222_n 0.00553065f $X=1.2 $Y=2.33 $X2=1.54 $Y2=1.845
cc_141 N_B0_c_169_n N_Y_c_222_n 0.0118918f $X=1.395 $Y=1.62 $X2=1.54 $Y2=1.845
cc_142 N_B0_M1001_g N_Y_c_223_n 0.00586282f $X=1.335 $Y=0.895 $X2=1.55 $Y2=1.22
cc_143 N_B0_c_164_n N_Y_c_223_n 0.00116649f $X=1.395 $Y=1.49 $X2=1.55 $Y2=1.22
cc_144 N_B0_c_169_n N_Y_c_223_n 0.00157776f $X=1.395 $Y=1.62 $X2=1.55 $Y2=1.22
cc_145 N_B0_M1001_g N_A_27_115#_c_283_n 8.81328e-19 $X=1.335 $Y=0.895 $X2=1.035
+ $Y2=1.16
cc_146 N_B0_c_168_n N_A_27_115#_c_283_n 0.00579405f $X=1.285 $Y=1.62 $X2=1.035
+ $Y2=1.16
cc_147 N_Y_c_227_n A_110_565# 0.00573878f $X=1.455 $Y=3.41 $X2=0.55 $Y2=2.825
cc_148 N_Y_c_219_n N_A_27_115#_c_283_n 0.0026548f $X=1.55 $Y=0.86 $X2=1.035
+ $Y2=1.16
cc_149 N_Y_c_223_n N_A_27_115#_c_283_n 0.00369865f $X=1.55 $Y=1.22 $X2=1.035
+ $Y2=1.16
