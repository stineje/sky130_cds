* File: sky130_osu_sc_15T_ls__and2_l.spice
* Created: Fri Nov 12 14:54:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_15T_ls__and2_l.pex.spice"
.subckt sky130_osu_sc_15T_ls__and2_l  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1003_b NSHORT L=0.15 W=0.52
+ AD=0.091 AS=0.0546 PD=0.87 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75000.5
+ SB=75000.7 A=0.078 P=1.34 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1001_d N_GND_M1003_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.091 PD=1.57 PS=0.87 NRD=0 NRS=16.152 M=1 R=3.46667
+ SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1002 N_A_27_115#_M1002_d N_A_M1002_g N_VDD_M1002_s N_VDD_M1002_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_B_M1005_g N_A_27_115#_M1002_d N_VDD_M1002_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_A_27_115#_M1004_g N_VDD_M1005_d N_VDD_M1002_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=5.64925 P=9.73
pX7_noxref noxref_8 A A PROBETYPE=1
pX8_noxref noxref_9 B B PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_15T_ls__and2_l.pxi.spice"
*
.ends
*
*
