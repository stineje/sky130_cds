* File: sky130_osu_sc_12T_ls__addh_1.spice
* Created: Fri Nov 12 15:33:21 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__addh_1.pex.spice"
.subckt sky130_osu_sc_12T_ls__addh_1  GND VDD CON B A S CO
* 
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_CON_M1006_g N_S_M1006_s N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0884 AS=0.1378 PD=0.86 PS=1.57 NRD=13.836 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1007 A_208_115# N_B_M1007_g N_GND_M1006_d N_GND_M1006_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.0884 PD=0.73 PS=0.86 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.7
+ SB=75000.5 A=0.078 P=1.34 MULT=1
MM1008 N_A_208_521#_M1008_d N_A_M1008_g A_208_115# N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.0546 PD=1.57 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_A_208_521#_M1001_g N_CO_M1001_s N_GND_M1006_b NSHORT
+ L=0.15 W=0.52 AD=0.0884 AS=0.1378 PD=0.86 PS=1.57 NRD=13.836 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75001.5 A=0.078 P=1.34 MULT=1
MM1010 N_CON_M1010_d N_A_208_521#_M1010_g N_GND_M1001_d N_GND_M1006_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.0884 PD=0.8 PS=0.86 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.7 SB=75001 A=0.078 P=1.34 MULT=1
MM1003 N_CON_M1010_d N_B_M1003_g N_CON_M1010_d N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.1
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1005 N_CON_M1010_d N_A_M1005_g N_CON_M1010_d N_GND_M1006_b NSHORT L=0.15
+ W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.5
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1004 N_VDD_M1004_d N_CON_M1004_g N_S_M1004_s N_VDD_M1004_b PHIGHVT L=0.15
+ W=1.26 AD=0.2142 AS=0.3339 PD=1.6 PS=3.05 NRD=9.3772 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1011 N_A_208_521#_M1011_d N_B_M1011_g N_VDD_M1004_d N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.2142 PD=1.54 PS=1.6 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.7 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 N_VDD_M1002_d N_A_M1002_g N_A_208_521#_M1011_d N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.2142 AS=0.1764 PD=1.6 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1009 N_CO_M1009_d N_A_208_521#_M1009_g N_VDD_M1002_d N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.2142 PD=3.05 PS=1.6 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75001.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_VDD_M1000_d N_A_208_521#_M1000_g N_CON_M1000_s N_VDD_M1004_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001 A=0.189 P=2.82 MULT=1
MM1012 A_668_521# N_B_M1012_g N_VDD_M1000_d N_VDD_M1004_b PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_CON_M1013_d N_A_M1013_g A_668_521# N_VDD_M1004_b PHIGHVT L=0.15 W=1.26
+ AD=0.3528 AS=0.1323 PD=3.08 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref N_GND_M1006_b N_VDD_M1004_b NWDIODE A=8.7138 P=12.58
pX15_noxref noxref_11 S S PROBETYPE=1
pX16_noxref noxref_12 CO CO PROBETYPE=1
pX17_noxref noxref_13 B B PROBETYPE=1
pX18_noxref noxref_14 CON CON PROBETYPE=1
pX19_noxref noxref_15 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_ls__addh_1.pxi.spice"
*
.ends
*
*
