* File: sky130_osu_sc_18T_hs__nand2_1.spice
* Created: Thu Oct 29 17:09:00 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_hs__nand2_1.pex.spice"
.subckt sky130_osu_sc_18T_hs__nand2_1  GND VDD A B Y
* 
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A_M1003_g N_Y_M1003_s N_GND_M1003_b NLOWVT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1003_b NLOWVT L=0.15 W=1
+ AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VDD_M1002_s N_VDD_M1002_b PSHORT L=0.15 W=3
+ AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2 SB=75000.6
+ A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_B_M1000_g N_Y_M1002_d N_VDD_M1002_b PSHORT L=0.15 W=3
+ AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75000.6 SB=75000.2
+ A=0.45 P=6.3 MULT=1
DX4_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=5.605 P=10.55
pX5_noxref noxref_7 A A PROBETYPE=1
pX6_noxref noxref_8 Y Y PROBETYPE=1
pX7_noxref noxref_9 B B PROBETYPE=1
c_157 A_110_115# 0 4.69618e-20 $X=0.55 $Y=0.575
*
.include "sky130_osu_sc_18T_hs__nand2_1.pxi.spice"
*
.ends
*
*
