* File: sky130_osu_sc_18T_hs__or2_4.spice
* Created: Fri Nov 12 13:52:39 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_hs__or2_4.pex.spice"
.subckt sky130_osu_sc_18T_hs__or2_4  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1005 N_A_27_617#_M1005_d N_B_M1005_g N_GND_M1005_s N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_A_27_617#_M1005_d N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1003_d N_A_27_617#_M1003_g N_GND_M1001_d N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1003_d N_A_27_617#_M1008_g N_GND_M1008_s N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1009 N_Y_M1009_d N_A_27_617#_M1009_g N_GND_M1008_s N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_Y_M1009_d N_A_27_617#_M1011_g N_GND_M1011_s N_GND_M1005_b NLOWVT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 A_110_617# N_B_M1004_g N_A_27_617#_M1004_s N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=5.5751 NRS=0 M=1 R=20 SA=75000.2
+ SB=75002.3 A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g A_110_617# N_VDD_M1004_b PSHORT L=0.15 W=3
+ AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=5.5751 M=1 R=20 SA=75000.6
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1002 N_Y_M1002_d N_A_27_617#_M1002_g N_VDD_M1000_d N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001 SB=75001.5
+ A=0.45 P=6.3 MULT=1
MM1006 N_Y_M1002_d N_A_27_617#_M1006_g N_VDD_M1006_s N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.5 SB=75001
+ A=0.45 P=6.3 MULT=1
MM1007 N_Y_M1007_d N_A_27_617#_M1007_g N_VDD_M1006_s N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.9 SB=75000.6
+ A=0.45 P=6.3 MULT=1
MM1010 N_Y_M1007_d N_A_27_617#_M1010_g N_VDD_M1010_s N_VDD_M1004_b PSHORT L=0.15
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75002.3
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX12_noxref N_GND_M1005_b N_VDD_M1004_b NWDIODE A=12.293 P=14.07
pX13_noxref noxref_8 B B PROBETYPE=1
pX14_noxref noxref_9 A A PROBETYPE=1
pX15_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_hs__or2_4.pxi.spice"
*
.ends
*
*
