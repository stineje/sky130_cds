* File: sky130_osu_sc_12T_ms__nor2_l.pex.spice
* Created: Fri Nov 12 15:25:37 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_L%GND 1 2 21 25 27 35 41 44
r26 41 44 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r27 33 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.74
r28 27 33 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.305
r29 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.74
r30 21 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r31 21 23 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r32 21 28 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r33 21 27 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r34 21 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r35 2 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.74
r36 1 25 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_L%VDD 1 13 15 21 27 30
r17 27 30 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=4.287
+ $X2=1.02 $Y2=4.287
r18 24 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=4.25
+ $X2=1.02 $Y2=4.25
r19 19 24 4.25596 $w=1.7e-07 $l=2.13185e-07 $layer=LI1_cond $X=1.05 $Y=4.135
+ $X2=1.197 $Y2=4.287
r20 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.05 $Y=4.135
+ $X2=1.05 $Y2=3.275
r21 15 24 3.30228 $w=3.05e-07 $l=2.32e-07 $layer=LI1_cond $X=0.965 $Y=4.287
+ $X2=1.197 $Y2=4.287
r22 15 17 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.965 $Y=4.287
+ $X2=0.34 $Y2=4.287
r23 13 24 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=4.135 $X2=1.02 $Y2=4.22
r24 13 17 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=4.135 $X2=0.34 $Y2=4.22
r25 1 21 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=3.025 $X2=1.05 $Y2=3.275
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_L%B 3 7 10 13 19 22
r47 19 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.65 $Y=2.85
+ $X2=0.65 $Y2=2.85
r48 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.65 $Y=2.065
+ $X2=0.65 $Y2=2.85
r49 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=1.98
+ $X2=0.65 $Y2=2.065
r50 13 15 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.565 $Y=1.98
+ $X2=0.415 $Y2=1.98
r51 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.98 $X2=0.415 $Y2=1.98
r52 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.98
+ $X2=0.415 $Y2=2.145
r53 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.98
+ $X2=0.415 $Y2=1.815
r54 7 12 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=0.475 $Y=3.445
+ $X2=0.475 $Y2=2.145
r55 3 11 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.475 $Y=0.755
+ $X2=0.475 $Y2=1.815
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_L%A 3 7 10 14 20
c31 20 0 1.46366e-19 $X=0.99 $Y=2.48
r32 14 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.99 $Y=2.48
+ $X2=0.99 $Y2=2.48
r33 14 17 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=2.48
+ $X2=0.99 $Y2=2.645
r34 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.645 $X2=0.99 $Y2=2.645
r35 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.645
+ $X2=0.942 $Y2=2.81
r36 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.942 $Y=2.645
+ $X2=0.942 $Y2=2.48
r37 7 11 884.521 $w=1.5e-07 $l=1.725e-06 $layer=POLY_cond $X=0.905 $Y=0.755
+ $X2=0.905 $Y2=2.48
r38 3 12 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.835 $Y=3.445
+ $X2=0.835 $Y2=2.81
.ends

.subckt PM_SKY130_OSU_SC_12T_MS__NOR2_L%Y 1 3 10 16 24 27 29 33 34
c39 10 0 1.46366e-19 $X=0.26 $Y=2.48
r40 33 34 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.69 $Y=1.37
+ $X2=0.545 $Y2=1.37
r41 29 30 0.0784968 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=0.26 $Y=2.48
+ $X2=0.26 $Y2=2.365
r42 27 34 0.181017 $w=1.75e-07 $l=2e-07 $layer=MET1_cond $X=0.345 $Y=1.367
+ $X2=0.545 $Y2=1.367
r43 24 30 0.615458 $w=1.75e-07 $l=6.8e-07 $layer=MET1_cond $X=0.257 $Y=1.685
+ $X2=0.257 $Y2=2.365
r44 21 27 0.0698411 $w=1.75e-07 $l=1.24451e-07 $layer=MET1_cond $X=0.257
+ $Y=1.455 $X2=0.345 $Y2=1.367
r45 21 24 0.20817 $w=1.75e-07 $l=2.3e-07 $layer=MET1_cond $X=0.257 $Y=1.455
+ $X2=0.257 $Y2=1.685
r46 19 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.37
+ $X2=0.69 $Y2=1.37
r47 16 19 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.69 $Y=0.74
+ $X2=0.69 $Y2=1.37
r48 10 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.48
+ $X2=0.26 $Y2=2.48
r49 10 13 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.26 $Y=2.48
+ $X2=0.26 $Y2=3.275
r50 3 13 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=3.025 $X2=0.26 $Y2=3.275
r51 1 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.74
.ends

