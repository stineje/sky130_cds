* File: sky130_osu_sc_12T_hs__or2_1.spice
* Created: Fri Nov 12 15:12:34 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_hs__or2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_1  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_A_27_521#_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_A_27_521#_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A_27_521#_M1002_g N_GND_M1001_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_B_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_M1004_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_521#_M1005_g N_VDD_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9449 P=7.95
pX7_noxref noxref_8 B B PROBETYPE=1
pX8_noxref noxref_9 A A PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_1.pxi.spice"
*
.ends
*
*
