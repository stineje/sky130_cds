* File: sky130_osu_sc_18T_hs__dffr_1.pex.spice
* Created: Thu Oct 29 17:07:28 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%GND 1 2 3 4 5 6 7 8 9 84 88 90 97 99 106
+ 115 117 127 129 139 141 148 150 157 159 166 185 187
c221 139 0 1.67294e-19 $X=6.09 $Y=0.825
c222 115 0 3.07193e-19 $X=2.59 $Y=0.825
c223 84 0 1.27355e-19 $X=-0.05 $Y=0
r224 185 187 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=0.152
+ $X2=9.175 $Y2=0.152
r225 179 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.152
+ $X2=8.85 $Y2=0.152
r226 164 180 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.152
r227 164 166 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.85 $Y=0.305
+ $X2=8.85 $Y2=0.825
r228 159 180 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.152
+ $X2=8.85 $Y2=0.152
r229 155 157 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.9 $Y=0.305
+ $X2=7.9 $Y2=0.825
r230 151 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.152
+ $X2=7.04 $Y2=0.152
r231 146 175 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.152
r232 146 148 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.04 $Y=0.305
+ $X2=7.04 $Y2=0.825
r233 142 174 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.152
+ $X2=6.09 $Y2=0.152
r234 141 175 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.152
+ $X2=7.04 $Y2=0.152
r235 137 174 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.152
r236 137 139 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=0.305
+ $X2=6.09 $Y2=0.825
r237 129 174 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.152
+ $X2=6.09 $Y2=0.152
r238 125 127 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.34 $Y=0.305
+ $X2=4.34 $Y2=0.825
r239 118 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.152
+ $X2=2.59 $Y2=0.152
r240 113 170 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.152
r241 113 115 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.59 $Y=0.305
+ $X2=2.59 $Y2=0.825
r242 109 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.152
+ $X2=2.07 $Y2=0.152
r243 108 170 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.152
+ $X2=2.59 $Y2=0.152
r244 104 169 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.152
r245 104 106 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.07 $Y=0.305
+ $X2=2.07 $Y2=0.825
r246 100 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.152
+ $X2=1.21 $Y2=0.152
r247 99 169 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.152
+ $X2=2.07 $Y2=0.152
r248 95 168 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.152
r249 95 97 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.21 $Y=0.305
+ $X2=1.21 $Y2=0.825
r250 90 168 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.152
+ $X2=1.21 $Y2=0.152
r251 86 88 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r252 84 86 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r253 84 91 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r254 84 179 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=9.175 $Y=0.152
+ $X2=8.935 $Y2=0.152
r255 84 187 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175 $Y=0.17
+ $X2=9.175 $Y2=0.17
r256 84 185 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335 $Y=0.17
+ $X2=0.335 $Y2=0.17
r257 84 155 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.9 $Y2=0.305
r258 84 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.815 $Y2=0.152
r259 84 160 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.152
+ $X2=7.985 $Y2=0.152
r260 84 125 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.34 $Y2=0.305
r261 84 117 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.255 $Y2=0.152
r262 84 130 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.152
+ $X2=4.425 $Y2=0.152
r263 84 159 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=8.765 $Y2=0.152
r264 84 160 19.2704 $w=3.03e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.152
+ $X2=7.985 $Y2=0.152
r265 84 150 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.815 $Y2=0.152
r266 84 151 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=7.135 $Y=0.152
+ $X2=7.125 $Y2=0.152
r267 84 141 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.955 $Y2=0.152
r268 84 142 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.455 $Y=0.152
+ $X2=6.175 $Y2=0.152
r269 84 129 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=5.775 $Y=0.152
+ $X2=6.005 $Y2=0.152
r270 84 130 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=0.152
+ $X2=4.425 $Y2=0.152
r271 84 117 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=0.152
+ $X2=4.255 $Y2=0.152
r272 84 118 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0.152
+ $X2=2.675 $Y2=0.152
r273 84 108 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.505 $Y2=0.152
r274 84 109 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=2.375 $Y=0.152
+ $X2=2.155 $Y2=0.152
r275 84 99 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.985 $Y2=0.152
r276 84 100 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=1.695 $Y=0.152
+ $X2=1.295 $Y2=0.152
r277 84 90 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=1.125 $Y2=0.152
r278 84 91 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.152
+ $X2=0.345 $Y2=0.152
r279 9 166 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.575 $X2=8.85 $Y2=0.825
r280 8 157 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.575 $X2=7.9 $Y2=0.825
r281 7 148 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.575 $X2=7.04 $Y2=0.825
r282 6 139 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.95
+ $Y=0.575 $X2=6.09 $Y2=0.825
r283 5 127 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.575 $X2=4.34 $Y2=0.825
r284 4 115 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=2.465
+ $Y=0.575 $X2=2.59 $Y2=0.825
r285 3 106 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.575 $X2=2.07 $Y2=0.825
r286 2 97 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.575 $X2=1.21 $Y2=0.825
r287 1 88 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%VDD 1 2 3 4 5 6 7 64 68 72 80 90 94 102
+ 106 114 118 126 130 136 150 155 159
r117 155 159 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.175
+ $Y=6.49 $X2=9.175 $Y2=6.49
r118 150 155 4.11698 $w=3.05e-07 $l=8.84e-06 $layer=MET1_cond $X=0.335 $Y=6.507
+ $X2=9.175 $Y2=6.507
r119 150 153 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.335
+ $Y=6.49 $X2=0.335 $Y2=6.49
r120 147 159 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=8.935 $Y=6.507
+ $X2=9.175 $Y2=6.507
r121 147 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=6.507
+ $X2=8.85 $Y2=6.507
r122 136 139 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=8.85 $Y=4.475
+ $X2=8.85 $Y2=5.835
r123 134 148 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.85 $Y=6.355
+ $X2=8.85 $Y2=6.507
r124 134 139 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.85 $Y=6.355
+ $X2=8.85 $Y2=5.835
r125 131 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=6.507
+ $X2=7.83 $Y2=6.507
r126 131 133 21.9153 $w=3.03e-07 $l=5.8e-07 $layer=LI1_cond $X=7.915 $Y=6.507
+ $X2=8.495 $Y2=6.507
r127 130 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=6.507
+ $X2=8.85 $Y2=6.507
r128 130 133 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=8.765 $Y=6.507
+ $X2=8.495 $Y2=6.507
r129 126 129 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.83 $Y=4.475
+ $X2=7.83 $Y2=5.835
r130 124 146 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.83 $Y=6.355
+ $X2=7.83 $Y2=6.507
r131 124 129 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.83 $Y=6.355
+ $X2=7.83 $Y2=5.835
r132 121 123 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.455 $Y=6.507
+ $X2=7.135 $Y2=6.507
r133 119 144 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.09 $Y2=6.507
r134 119 121 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6.175 $Y=6.507
+ $X2=6.455 $Y2=6.507
r135 118 146 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=6.507
+ $X2=7.83 $Y2=6.507
r136 118 123 23.0489 $w=3.03e-07 $l=6.1e-07 $layer=LI1_cond $X=7.745 $Y=6.507
+ $X2=7.135 $Y2=6.507
r137 114 117 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.09 $Y=3.455
+ $X2=6.09 $Y2=5.835
r138 112 144 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=6.507
r139 112 117 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.09 $Y=6.355
+ $X2=6.09 $Y2=5.835
r140 109 111 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=6.507
+ $X2=5.775 $Y2=6.507
r141 107 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=6.507
+ $X2=4.34 $Y2=6.507
r142 107 109 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.425 $Y=6.507
+ $X2=5.095 $Y2=6.507
r143 106 144 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=6.09 $Y2=6.507
r144 106 111 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=6.005 $Y=6.507
+ $X2=5.775 $Y2=6.507
r145 102 105 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.34 $Y=3.795
+ $X2=4.34 $Y2=5.835
r146 100 143 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.34 $Y=6.355
+ $X2=4.34 $Y2=6.507
r147 100 105 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.34 $Y=6.355
+ $X2=4.34 $Y2=5.835
r148 97 99 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=6.507
+ $X2=3.735 $Y2=6.507
r149 95 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=6.507
+ $X2=2.59 $Y2=6.507
r150 95 97 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.675 $Y=6.507
+ $X2=3.055 $Y2=6.507
r151 94 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=6.507
+ $X2=4.34 $Y2=6.507
r152 94 99 19.6482 $w=3.03e-07 $l=5.2e-07 $layer=LI1_cond $X=4.255 $Y=6.507
+ $X2=3.735 $Y2=6.507
r153 90 93 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.59 $Y=3.795
+ $X2=2.59 $Y2=5.835
r154 88 141 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.59 $Y=6.355
+ $X2=2.59 $Y2=6.507
r155 88 93 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.59 $Y=6.355
+ $X2=2.59 $Y2=5.835
r156 85 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=6.507
+ $X2=2 $Y2=6.507
r157 85 87 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=2.085 $Y=6.507
+ $X2=2.375 $Y2=6.507
r158 84 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=6.507
+ $X2=2.59 $Y2=6.507
r159 84 87 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=6.507
+ $X2=2.375 $Y2=6.507
r160 80 83 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2 $Y=4.475 $X2=2
+ $Y2=5.835
r161 78 140 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2 $Y=6.355 $X2=2
+ $Y2=6.507
r162 78 83 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2 $Y=6.355 $X2=2
+ $Y2=5.835
r163 75 77 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.015 $Y=6.507
+ $X2=1.695 $Y2=6.507
r164 73 153 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=0.172 $Y2=6.507
r165 73 75 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.345 $Y=6.507
+ $X2=1.015 $Y2=6.507
r166 72 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=6.507
+ $X2=2 $Y2=6.507
r167 72 77 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=1.915 $Y=6.507
+ $X2=1.695 $Y2=6.507
r168 68 71 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r169 66 153 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.172 $Y2=6.507
r170 66 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=6.355
+ $X2=0.26 $Y2=5.835
r171 64 153 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.13 $Y=6.355 $X2=0.335 $Y2=6.44
r172 64 159 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.97 $Y=6.355 $X2=9.175 $Y2=6.44
r173 64 146 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=7.61 $Y=6.355 $X2=7.815 $Y2=6.44
r174 64 143 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.21 $Y=6.355 $X2=4.415 $Y2=6.44
r175 64 133 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=8.29 $Y=6.355 $X2=8.495 $Y2=6.44
r176 64 123 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.93 $Y=6.355 $X2=7.135 $Y2=6.44
r177 64 121 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.25 $Y=6.355 $X2=6.455 $Y2=6.44
r178 64 111 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.57 $Y=6.355 $X2=5.775 $Y2=6.44
r179 64 109 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.89 $Y=6.355 $X2=5.095 $Y2=6.44
r180 64 99 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.53 $Y=6.355 $X2=3.735 $Y2=6.44
r181 64 97 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.85 $Y=6.355 $X2=3.055 $Y2=6.44
r182 64 87 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.17 $Y=6.355 $X2=2.375 $Y2=6.44
r183 64 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.49 $Y=6.355 $X2=1.695 $Y2=6.44
r184 64 75 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.81 $Y=6.355 $X2=1.015 $Y2=6.44
r185 7 139 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=3.085 $X2=8.85 $Y2=5.835
r186 7 136 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=3.085 $X2=8.85 $Y2=4.475
r187 6 129 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=4.085 $X2=7.83 $Y2=5.835
r188 6 126 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=4.085 $X2=7.83 $Y2=4.475
r189 5 117 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=5.95
+ $Y=3.085 $X2=6.09 $Y2=5.835
r190 5 114 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=5.95
+ $Y=3.085 $X2=6.09 $Y2=3.455
r191 4 105 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=4.2
+ $Y=3.085 $X2=4.34 $Y2=5.835
r192 4 102 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=4.2
+ $Y=3.085 $X2=4.34 $Y2=3.795
r193 3 93 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3
+ $X=2.465 $Y=3.085 $X2=2.59 $Y2=5.835
r194 3 90 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3
+ $X=2.465 $Y=3.085 $X2=2.59 $Y2=3.795
r195 2 83 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=4.085 $X2=2 $Y2=5.835
r196 2 80 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=4.085 $X2=2 $Y2=4.475
r197 1 71 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r198 1 68 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%RN 3 5 7 9 16 17
c38 17 0 7.48684e-20 $X=0.325 $Y=3.33
c39 3 0 1.0751e-19 $X=0.475 $Y=1.075
r40 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.32 $Y=3.33
+ $X2=0.32 $Y2=3.33
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=2.305 $X2=0.53 $Y2=2.305
r42 10 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.32 $Y=2.47 $X2=0.32
+ $Y2=3.33
r43 9 12 8.98947 $w=2.85e-07 $l=2.1e-07 $layer=LI1_cond $X=0.32 $Y=2.305
+ $X2=0.53 $Y2=2.305
r44 9 10 3.76007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.305
+ $X2=0.32 $Y2=2.47
r45 5 13 38.945 $w=2.68e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.53 $Y2=2.305
r46 5 7 1084.5 $w=1.5e-07 $l=2.115e-06 $layer=POLY_cond $X=0.475 $Y=2.47
+ $X2=0.475 $Y2=4.585
r47 1 13 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.53 $Y2=2.305
r48 1 3 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.475 $Y=2.135
+ $X2=0.475 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_110_115# 1 2 7 9 12 16 18 20 23 27 32
+ 33 34 40 42 43 46 49 50 56 63
c173 46 0 9.11346e-20 $X=1.23 $Y=1.48
c174 43 0 1.63751e-20 $X=1.375 $Y=1.48
c175 40 0 7.48684e-20 $X=0.87 $Y=2.74
c176 16 0 1.88625e-19 $X=7.615 $Y=5.085
r177 60 63 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.685 $Y=1.59
+ $X2=7.81 $Y2=1.59
r178 58 60 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.615 $Y=1.59
+ $X2=7.685 $Y2=1.59
r179 54 56 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.23 $Y=1.59
+ $X2=1.425 $Y2=1.59
r180 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.59 $X2=1.23 $Y2=1.59
r181 50 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.81
+ $Y=1.59 $X2=7.81 $Y2=1.59
r182 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.81 $Y=1.48
+ $X2=7.81 $Y2=1.48
r183 46 53 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.23 $Y=1.48
+ $X2=1.23 $Y2=1.59
r184 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.48
+ $X2=1.23 $Y2=1.48
r185 43 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.375 $Y=1.48
+ $X2=1.23 $Y2=1.48
r186 42 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.665 $Y=1.48
+ $X2=7.81 $Y2=1.48
r187 42 43 6.05653 $w=1.7e-07 $l=6.29e-06 $layer=MET1_cond $X=7.665 $Y=1.48
+ $X2=1.375 $Y2=1.48
r188 38 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=2.74
+ $X2=0.87 $Y2=2.74
r189 35 37 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.87 $Y2=1.59
r190 34 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=1.59
+ $X2=0.87 $Y2=1.59
r191 33 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=1.23 $Y2=1.59
r192 33 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.145 $Y=1.59
+ $X2=0.955 $Y2=1.59
r193 32 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.655
+ $X2=0.87 $Y2=2.74
r194 31 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=1.59
r195 31 32 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.87 $Y=1.675
+ $X2=0.87 $Y2=2.655
r196 27 29 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.69 $Y=3.455
+ $X2=0.69 $Y2=5.835
r197 25 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=2.74
r198 25 27 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.69 $Y=2.825
+ $X2=0.69 $Y2=3.455
r199 21 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=1.59
r200 21 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=0.825
r201 18 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.685 $Y=1.425
+ $X2=7.685 $Y2=1.59
r202 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.685 $Y=1.425
+ $X2=7.685 $Y2=0.945
r203 14 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.755
+ $X2=7.615 $Y2=1.59
r204 14 16 1707.51 $w=1.5e-07 $l=3.33e-06 $layer=POLY_cond $X=7.615 $Y=1.755
+ $X2=7.615 $Y2=5.085
r205 10 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.755
+ $X2=1.425 $Y2=1.59
r206 10 12 1707.51 $w=1.5e-07 $l=3.33e-06 $layer=POLY_cond $X=1.425 $Y=1.755
+ $X2=1.425 $Y2=5.085
r207 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.425
+ $X2=1.425 $Y2=1.59
r208 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.425
+ $X2=1.425 $Y2=0.945
r209 2 29 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r210 2 27 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=3.455
r211 1 23 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_342_518# 1 2 9 13 16 18 19 20 21 22 24
+ 27 31 37 39 42
c86 42 0 1.71621e-19 $X=3.457 $Y=1.415
c87 19 0 1.29912e-19 $X=3.28 $Y=1.765
r88 41 42 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.457 $Y=1.245
+ $X2=3.457 $Y2=1.415
r89 37 45 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.755
+ $X2=1.892 $Y2=2.92
r90 37 44 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.892 $Y=2.755
+ $X2=1.892 $Y2=2.59
r91 36 39 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.94 $Y=2.755
+ $X2=2.11 $Y2=2.755
r92 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.755 $X2=1.94 $Y2=2.755
r93 31 33 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=3.465 $Y=3.455
+ $X2=3.465 $Y2=5.835
r94 29 31 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=3.465 $Y=3.27
+ $X2=3.465 $Y2=3.455
r95 27 41 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=3.465 $Y=0.825
+ $X2=3.465 $Y2=1.245
r96 24 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=1.68
+ $X2=3.365 $Y2=1.415
r97 21 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.295 $Y=3.185
+ $X2=3.465 $Y2=3.27
r98 21 22 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.295 $Y=3.185
+ $X2=2.195 $Y2=3.185
r99 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=1.765
+ $X2=3.365 $Y2=1.68
r100 19 20 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.28 $Y=1.765
+ $X2=2.195 $Y2=1.765
r101 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=3.1
+ $X2=2.195 $Y2=3.185
r102 17 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=2.92
+ $X2=2.11 $Y2=2.755
r103 17 18 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.11 $Y=2.92
+ $X2=2.11 $Y2=3.1
r104 16 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=2.59
+ $X2=2.11 $Y2=2.755
r105 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=1.85
+ $X2=2.195 $Y2=1.765
r106 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.11 $Y=1.85
+ $X2=2.11 $Y2=2.59
r107 13 44 843.5 $w=1.5e-07 $l=1.645e-06 $layer=POLY_cond $X=1.855 $Y=0.945
+ $X2=1.855 $Y2=2.59
r108 9 45 1110.14 $w=1.5e-07 $l=2.165e-06 $layer=POLY_cond $X=1.785 $Y=5.085
+ $X2=1.785 $Y2=2.92
r109 2 33 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=3.24
+ $Y=3.085 $X2=3.465 $Y2=5.835
r110 2 31 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=3.24
+ $Y=3.085 $X2=3.465 $Y2=3.455
r111 1 27 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=3.24
+ $Y=0.575 $X2=3.465 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%D 3 7 10 12 16
c41 16 0 1.12321e-19 $X=2.865 $Y=2.22
c42 10 0 1.41836e-19 $X=2.865 $Y=2.22
r43 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=2.22
+ $X2=2.865 $Y2=2.385
r44 16 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=2.22
+ $X2=2.865 $Y2=2.055
r45 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=2.22 $X2=2.865 $Y2=2.22
r46 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.865 $Y=2.22
+ $X2=2.865 $Y2=2.22
r47 7 18 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=2.805 $Y=4.585
+ $X2=2.805 $Y2=2.385
r48 3 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.805 $Y=1.075
+ $X2=2.805 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%CK 3 7 10 13 17 18 20 23 24 25 26 30 31
+ 35 36 38 39 40 41 42 43 46 50 52 54 59 63 66 70
c219 63 0 1.29912e-19 $X=3.705 $Y=1.685
c220 59 0 1.41836e-19 $X=3.225 $Y=2.765
c221 39 0 6.79641e-20 $X=5.06 $Y=2.59
c222 30 0 1.98654e-19 $X=3.705 $Y=1.85
c223 26 0 1.86602e-19 $X=3.62 $Y=2.59
r224 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=2.765 $X2=6.45 $Y2=2.765
r225 70 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=2.765
+ $X2=5.455 $Y2=2.93
r226 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=2.765 $X2=5.455 $Y2=2.765
r227 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.765
+ $X2=3.225 $Y2=2.93
r228 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=2.765 $X2=3.225 $Y2=2.765
r229 54 74 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.45 $Y=2.59
+ $X2=6.45 $Y2=2.765
r230 52 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.45 $Y=2.59
+ $X2=6.45 $Y2=2.59
r231 50 69 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.455 $Y=2.59
+ $X2=5.455 $Y2=2.765
r232 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.455 $Y=2.59
+ $X2=5.455 $Y2=2.59
r233 46 58 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.225 $Y=2.59
+ $X2=3.225 $Y2=2.765
r234 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.225 $Y=2.59
+ $X2=3.225 $Y2=2.59
r235 43 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.6 $Y=2.59
+ $X2=5.455 $Y2=2.59
r236 42 52 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.305 $Y=2.59
+ $X2=6.45 $Y2=2.59
r237 42 43 0.678832 $w=1.7e-07 $l=7.05e-07 $layer=MET1_cond $X=6.305 $Y=2.59
+ $X2=5.6 $Y2=2.59
r238 41 45 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.37 $Y=2.59
+ $X2=3.225 $Y2=2.59
r239 40 49 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.31 $Y=2.59
+ $X2=5.455 $Y2=2.59
r240 40 41 1.86799 $w=1.7e-07 $l=1.94e-06 $layer=MET1_cond $X=5.31 $Y=2.59
+ $X2=3.37 $Y2=2.59
r241 38 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.59
+ $X2=5.455 $Y2=2.59
r242 38 39 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.37 $Y=2.59
+ $X2=5.06 $Y2=2.59
r243 36 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.85
+ $X2=4.975 $Y2=1.685
r244 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.85 $X2=4.975 $Y2=1.85
r245 33 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=2.505
+ $X2=5.06 $Y2=2.59
r246 33 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.975 $Y=2.505
+ $X2=4.975 $Y2=1.85
r247 31 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.85
+ $X2=3.705 $Y2=1.685
r248 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.85 $X2=3.705 $Y2=1.85
r249 28 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.705 $Y=2.505
+ $X2=3.705 $Y2=1.85
r250 27 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.59
+ $X2=3.225 $Y2=2.59
r251 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.59
+ $X2=3.705 $Y2=2.505
r252 26 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.62 $Y=2.59
+ $X2=3.31 $Y2=2.59
r253 24 25 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.332 $Y=1.685
+ $X2=6.332 $Y2=1.835
r254 23 75 38.571 $w=3.25e-07 $l=1.87029e-07 $layer=POLY_cond $X=6.36 $Y=2.6
+ $X2=6.407 $Y2=2.765
r255 23 25 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.36 $Y=2.6
+ $X2=6.36 $Y2=1.835
r256 18 75 38.571 $w=3.25e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.305 $Y=2.93
+ $X2=6.407 $Y2=2.765
r257 18 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=6.305 $Y=2.93
+ $X2=6.305 $Y2=4.585
r258 17 24 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.305 $Y=1.075
+ $X2=6.305 $Y2=1.685
r259 13 72 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.515 $Y=4.585
+ $X2=5.515 $Y2=2.93
r260 10 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.915 $Y=1.075
+ $X2=4.915 $Y2=1.685
r261 7 63 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.765 $Y=1.075
+ $X2=3.765 $Y2=1.685
r262 3 61 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.165 $Y=4.585
+ $X2=3.165 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_217_817# 1 2 9 13 17 21 23 24 25 26 29
+ 33 34 37 41 42 48 49 56
c140 41 0 1.35571e-19 $X=4.06 $Y=1.85
c141 37 0 1.5821e-19 $X=4.295 $Y=2.765
c142 26 0 6.79641e-20 $X=4.48 $Y=2.765
c143 24 0 1.86602e-19 $X=4.2 $Y=2.765
c144 21 0 6.36774e-20 $X=4.555 $Y=4.585
c145 13 0 6.36774e-20 $X=4.125 $Y=4.585
r146 49 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.85 $X2=4.295 $Y2=1.85
r147 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.205 $Y=1.85
+ $X2=4.205 $Y2=1.85
r148 45 56 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=1.64 $Y=1.85
+ $X2=1.64 $Y2=0.825
r149 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.64 $Y=1.85
+ $X2=1.64 $Y2=1.85
r150 42 44 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.785 $Y=1.85
+ $X2=1.64 $Y2=1.85
r151 41 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.85
+ $X2=4.205 $Y2=1.85
r152 41 42 2.19056 $w=1.7e-07 $l=2.275e-06 $layer=MET1_cond $X=4.06 $Y=1.85
+ $X2=1.785 $Y2=1.85
r153 40 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=1.935
+ $X2=1.64 $Y2=1.85
r154 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=2.765 $X2=4.295 $Y2=2.765
r155 35 49 2.3025 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.295 $Y=1.935
+ $X2=4.205 $Y2=1.81
r156 35 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.295 $Y=1.935
+ $X2=4.295 $Y2=2.765
r157 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=2.02
+ $X2=1.64 $Y2=1.935
r158 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.555 $Y=2.02
+ $X2=1.295 $Y2=2.02
r159 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.21 $Y=4.475
+ $X2=1.21 $Y2=5.835
r160 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.295 $Y2=2.02
r161 27 29 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=1.21 $Y=2.105
+ $X2=1.21 $Y2=4.475
r162 26 38 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=2.765
+ $X2=4.295 $Y2=2.765
r163 25 53 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=4.48 $Y=1.85
+ $X2=4.295 $Y2=1.85
r164 24 38 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=2.765
+ $X2=4.295 $Y2=2.765
r165 23 53 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=4.2 $Y=1.85
+ $X2=4.295 $Y2=1.85
r166 19 26 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.48 $Y2=2.765
r167 19 21 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.555 $Y=2.9
+ $X2=4.555 $Y2=4.585
r168 15 25 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.48 $Y2=1.85
r169 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.555 $Y=1.715
+ $X2=4.555 $Y2=1.075
r170 11 24 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=2.9
+ $X2=4.2 $Y2=2.765
r171 11 13 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=4.125 $Y=2.9
+ $X2=4.125 $Y2=4.585
r172 7 23 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.125 $Y=1.715
+ $X2=4.2 $Y2=1.85
r173 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.125 $Y=1.715
+ $X2=4.125 $Y2=1.075
r174 2 31 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=4.085 $X2=1.21 $Y2=5.835
r175 2 29 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=4.085 $X2=1.21 $Y2=4.475
r176 1 56 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.575 $X2=1.64 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_618_89# 1 2 7 9 11 12 13 16 18 22 24
+ 27 30 33 35 36 37 40 44 47 50 55 56 59 63 66
c187 33 0 1.98654e-19 $X=3.285 $Y=1.76
c188 16 0 1.12321e-19 $X=3.765 $Y=4.585
r189 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=3.185
+ $X2=6.795 $Y2=3.185
r190 57 59 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.52 $Y=2.19
+ $X2=6.795 $Y2=2.19
r191 55 63 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=3.1
+ $X2=6.795 $Y2=3.185
r192 54 59 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.275
+ $X2=6.795 $Y2=2.19
r193 54 55 50.8333 $w=1.78e-07 $l=8.25e-07 $layer=LI1_cond $X=6.795 $Y=2.275
+ $X2=6.795 $Y2=3.1
r194 50 52 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.52 $Y=3.455
+ $X2=6.52 $Y2=5.835
r195 48 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=3.27
+ $X2=6.52 $Y2=3.185
r196 48 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.52 $Y=3.27
+ $X2=6.52 $Y2=3.455
r197 47 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.105
+ $X2=6.52 $Y2=2.19
r198 46 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.935
+ $X2=6.52 $Y2=1.85
r199 46 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=1.935
+ $X2=6.52 $Y2=2.105
r200 42 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=1.765
+ $X2=6.52 $Y2=1.85
r201 42 44 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.52 $Y=1.765
+ $X2=6.52 $Y2=0.825
r202 40 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.85
+ $X2=5.455 $Y2=2.015
r203 40 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.85
+ $X2=5.455 $Y2=1.685
r204 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.85 $X2=5.455 $Y2=1.85
r205 37 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=1.85
+ $X2=6.52 $Y2=1.85
r206 37 39 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.435 $Y=1.85
+ $X2=5.455 $Y2=1.85
r207 31 33 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.165 $Y=1.76
+ $X2=3.285 $Y2=1.76
r208 30 66 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.515 $Y=1.075
+ $X2=5.515 $Y2=1.685
r209 27 67 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.395 $Y=2.225
+ $X2=5.395 $Y2=2.015
r210 25 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.99 $Y=2.3
+ $X2=4.915 $Y2=2.3
r211 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.32 $Y=2.3
+ $X2=5.395 $Y2=2.225
r212 24 25 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.32 $Y=2.3
+ $X2=4.99 $Y2=2.3
r213 20 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.915 $Y=2.375
+ $X2=4.915 $Y2=2.3
r214 20 22 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=4.915 $Y=2.375
+ $X2=4.915 $Y2=4.585
r215 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=2.3
+ $X2=3.765 $Y2=2.3
r216 18 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=2.3
+ $X2=4.915 $Y2=2.3
r217 18 19 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.84 $Y=2.3 $X2=3.84
+ $Y2=2.3
r218 14 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=2.375
+ $X2=3.765 $Y2=2.3
r219 14 16 1133.21 $w=1.5e-07 $l=2.21e-06 $layer=POLY_cond $X=3.765 $Y=2.375
+ $X2=3.765 $Y2=4.585
r220 12 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=2.3
+ $X2=3.765 $Y2=2.3
r221 12 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.69 $Y=2.3
+ $X2=3.36 $Y2=2.3
r222 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.285 $Y=2.225
+ $X2=3.36 $Y2=2.3
r223 10 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.835
+ $X2=3.285 $Y2=1.76
r224 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.285 $Y=1.835
+ $X2=3.285 $Y2=2.225
r225 7 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.685
+ $X2=3.165 $Y2=1.76
r226 7 9 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.165 $Y=1.685
+ $X2=3.165 $Y2=1.075
r227 2 52 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=5.835
r228 2 50 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.38
+ $Y=3.085 $X2=6.52 $Y2=3.455
r229 1 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.575 $X2=6.52 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_1160_89# 1 2 9 13 21 24 25 26 27 28 31
+ 35 36 39 42 44 45 46 49 52 53 57 62 63
c160 62 0 2.20654e-19 $X=8.52 $Y=2.19
c161 27 0 8.77106e-20 $X=8.61 $Y=2.855
r162 62 64 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=2.19
+ $X2=8.522 $Y2=2.355
r163 62 63 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.522 $Y=2.19
+ $X2=8.522 $Y2=2.025
r164 57 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=2.19
+ $X2=5.935 $Y2=2.355
r165 57 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=2.19
+ $X2=5.935 $Y2=2.025
r166 53 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.52
+ $Y=2.19 $X2=8.52 $Y2=2.19
r167 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.52 $Y=2.19
+ $X2=8.52 $Y2=2.19
r168 49 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.935
+ $Y=2.19 $X2=5.935 $Y2=2.19
r169 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.935 $Y=2.19
+ $X2=5.935 $Y2=2.19
r170 46 48 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=2.19
+ $X2=5.935 $Y2=2.19
r171 45 52 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.375 $Y=2.19
+ $X2=8.52 $Y2=2.19
r172 45 46 2.20982 $w=1.7e-07 $l=2.295e-06 $layer=MET1_cond $X=8.375 $Y=2.19
+ $X2=6.08 $Y2=2.19
r173 43 53 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.555 $Y=2.19
+ $X2=8.52 $Y2=2.19
r174 43 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=2.19
+ $X2=7.47 $Y2=2.19
r175 41 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=2.275
+ $X2=7.47 $Y2=2.19
r176 41 42 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.47 $Y=2.275
+ $X2=7.47 $Y2=3.695
r177 37 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=2.105
+ $X2=7.47 $Y2=2.19
r178 37 39 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=7.47 $Y=2.105
+ $X2=7.47 $Y2=0.825
r179 35 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=3.78
+ $X2=7.47 $Y2=3.695
r180 35 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.385 $Y=3.78
+ $X2=7.125 $Y2=3.78
r181 31 33 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.04 $Y=4.475
+ $X2=7.04 $Y2=5.835
r182 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=3.865
+ $X2=7.125 $Y2=3.78
r183 29 31 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.04 $Y=3.865
+ $X2=7.04 $Y2=4.475
r184 27 28 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=2.855
+ $X2=8.61 $Y2=3.005
r185 27 64 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=8.585 $Y=2.855
+ $X2=8.585 $Y2=2.355
r186 26 63 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.585 $Y=1.8
+ $X2=8.585 $Y2=2.025
r187 25 26 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.61 $Y=1.65 $X2=8.61
+ $Y2=1.8
r188 24 28 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=8.635 $Y=4.585
+ $X2=8.635 $Y2=3.005
r189 21 25 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.635 $Y=1.075
+ $X2=8.635 $Y2=1.65
r190 13 59 1143.47 $w=1.5e-07 $l=2.23e-06 $layer=POLY_cond $X=5.875 $Y=4.585
+ $X2=5.875 $Y2=2.355
r191 9 58 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.875 $Y=1.075
+ $X2=5.875 $Y2=2.025
r192 2 33 240 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=4.085 $X2=7.04 $Y2=5.835
r193 2 31 240 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=2 $X=6.915
+ $Y=4.085 $X2=7.04 $Y2=4.475
r194 1 39 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.575 $X2=7.47 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%A_998_115# 1 2 9 11 13 15 16 17 18 21 25
+ 31 32 35 38 39
c131 35 0 1.57671e-19 $X=4.635 $Y=1.85
c132 32 0 1.5821e-19 $X=4.78 $Y=1.85
c133 15 0 1.67294e-19 $X=5.045 $Y=1.43
r134 39 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.85 $X2=7.13 $Y2=1.85
r135 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=1.85
+ $X2=7.13 $Y2=1.85
r136 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=1.85
+ $X2=4.635 $Y2=1.85
r137 32 34 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.78 $Y=1.85
+ $X2=4.635 $Y2=1.85
r138 31 38 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=1.85
+ $X2=7.13 $Y2=1.85
r139 31 32 2.12316 $w=1.7e-07 $l=2.205e-06 $layer=MET1_cond $X=6.985 $Y=1.85
+ $X2=4.78 $Y2=1.85
r140 30 35 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.635 $Y=3.1
+ $X2=4.635 $Y2=1.85
r141 29 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.635 $Y=1.515
+ $X2=4.635 $Y2=1.85
r142 25 27 69.1466 $w=3.38e-07 $l=2.04e-06 $layer=LI1_cond $X=5.215 $Y=3.795
+ $X2=5.215 $Y2=5.835
r143 23 25 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=5.215 $Y=3.27
+ $X2=5.215 $Y2=3.795
r144 19 21 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=5.215 $Y=1.345
+ $X2=5.215 $Y2=0.825
r145 18 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.72 $Y=3.185
+ $X2=4.635 $Y2=3.1
r146 17 23 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=3.185
+ $X2=5.215 $Y2=3.27
r147 17 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=3.185
+ $X2=4.72 $Y2=3.185
r148 16 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.72 $Y=1.43
+ $X2=4.635 $Y2=1.515
r149 15 19 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.045 $Y=1.43
+ $X2=5.215 $Y2=1.345
r150 15 16 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.045 $Y=1.43
+ $X2=4.72 $Y2=1.43
r151 11 43 38.6212 $w=3.33e-07 $l=2.06325e-07 $layer=POLY_cond $X=7.255 $Y=2.015
+ $X2=7.162 $Y2=1.85
r152 11 13 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=7.255 $Y=2.015
+ $X2=7.255 $Y2=5.085
r153 7 43 39.3449 $w=3.33e-07 $l=2.11447e-07 $layer=POLY_cond $X=7.255 $Y=1.68
+ $X2=7.162 $Y2=1.85
r154 7 9 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=7.255 $Y=1.68
+ $X2=7.255 $Y2=0.945
r155 2 27 171.429 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=3 $X=4.99
+ $Y=3.085 $X2=5.215 $Y2=5.835
r156 2 25 171.429 $w=1.7e-07 $l=8.1477e-07 $layer=licon1_PDIFF $count=3 $X=4.99
+ $Y=3.085 $X2=5.215 $Y2=3.795
r157 1 21 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=4.99
+ $Y=0.575 $X2=5.215 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%QN 1 2 9 13 17 19 20 21 22 26 27 31 32
c80 32 0 8.77106e-20 $X=8.425 $Y=2.96
c81 21 0 9.99996e-20 $X=8.92 $Y=2.765
c82 19 0 1.20654e-19 $X=8.92 $Y=1.85
c83 17 0 1.88625e-19 $X=8.42 $Y=0.825
r84 39 41 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=8.42 $Y=4.475
+ $X2=8.42 $Y2=5.835
r85 31 39 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=8.42 $Y=2.96
+ $X2=8.42 $Y2=4.475
r86 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.42 $Y=2.96
+ $X2=8.42 $Y2=2.96
r87 28 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.42 $Y=2.85
+ $X2=8.42 $Y2=2.96
r88 27 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=2.395
+ $X2=9.005 $Y2=2.56
r89 27 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=2.395
+ $X2=9.005 $Y2=2.23
r90 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=2.395 $X2=9.005 $Y2=2.395
r91 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.005 $Y=2.68
+ $X2=9.005 $Y2=2.395
r92 23 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.005 $Y=1.935
+ $X2=9.005 $Y2=2.395
r93 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.505 $Y=2.765
+ $X2=8.42 $Y2=2.85
r94 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=2.765
+ $X2=9.005 $Y2=2.68
r95 21 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=2.765
+ $X2=8.505 $Y2=2.765
r96 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=1.85
+ $X2=9.005 $Y2=1.935
r97 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.92 $Y=1.85
+ $X2=8.505 $Y2=1.85
r98 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=1.765
+ $X2=8.505 $Y2=1.85
r99 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=8.42 $Y=1.765
+ $X2=8.42 $Y2=0.825
r100 13 36 1038.35 $w=1.5e-07 $l=2.025e-06 $layer=POLY_cond $X=9.065 $Y=4.585
+ $X2=9.065 $Y2=2.56
r101 9 35 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=9.065 $Y=1.075
+ $X2=9.065 $Y2=2.23
r102 2 41 240 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=3.085 $X2=8.42 $Y2=5.835
r103 2 39 240 $w=1.7e-07 $l=1.45115e-06 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=3.085 $X2=8.42 $Y2=4.475
r104 1 17 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.575 $X2=8.42 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__DFFR_1%Q 1 2 9 13 18 21 24 26
r21 26 29 6.68493 $w=2.19e-07 $l=1.2e-07 $layer=LI1_cond $X=9.275 $Y=3.287
+ $X2=9.395 $Y2=3.287
r22 24 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=3.33
+ $X2=9.275 $Y2=3.33
r23 19 21 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.28 $Y=1.515
+ $X2=9.395 $Y2=1.515
r24 18 29 2.22295 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.395 $Y=3.16
+ $X2=9.395 $Y2=3.287
r25 17 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.6
+ $X2=9.395 $Y2=1.515
r26 17 18 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=9.395 $Y=1.6
+ $X2=9.395 $Y2=3.16
r27 13 15 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=9.28 $Y=4.475
+ $X2=9.28 $Y2=5.835
r28 11 26 2.22295 $w=1.7e-07 $l=1.30476e-07 $layer=LI1_cond $X=9.28 $Y=3.415
+ $X2=9.275 $Y2=3.287
r29 11 13 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=9.28 $Y=3.415
+ $X2=9.28 $Y2=4.475
r30 7 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=1.43 $X2=9.28
+ $Y2=1.515
r31 7 9 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.28 $Y=1.43 $X2=9.28
+ $Y2=0.825
r32 2 15 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=3.085 $X2=9.28 $Y2=5.835
r33 2 13 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=3.085 $X2=9.28 $Y2=4.475
r34 1 9 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.575 $X2=9.28 $Y2=0.825
.ends

