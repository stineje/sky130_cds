* File: sky130_osu_sc_18T_ls__or2_8.spice
* Created: Thu Oct 29 17:38:10 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ls__or2_8.pex.spice"
.subckt sky130_osu_sc_18T_ls__or2_8  GND VDD B A Y
* 
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1006 N_A_27_617#_M1006_d N_B_M1006_g N_GND_M1006_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1000 N_GND_M1000_d N_A_M1000_g N_A_27_617#_M1006_d N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A_27_617#_M1001_g N_GND_M1000_d N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1001_d N_A_27_617#_M1007_g N_GND_M1007_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1010_d N_A_27_617#_M1010_g N_GND_M1007_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1010_d N_A_27_617#_M1012_g N_GND_M1012_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1013 N_Y_M1013_d N_A_27_617#_M1013_g N_GND_M1012_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1013_d N_A_27_617#_M1015_g N_GND_M1015_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1016 N_Y_M1016_d N_A_27_617#_M1016_g N_GND_M1015_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1018 N_Y_M1016_d N_A_27_617#_M1018_g N_GND_M1018_s N_GND_M1006_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 A_110_617# N_B_M1005_g N_A_27_617#_M1005_s N_VDD_M1005_b PHIGHVT L=0.15
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=5.5751 NRS=0 M=1 R=20 SA=75000.2
+ SB=75004.1 A=0.45 P=6.3 MULT=1
MM1017 N_VDD_M1017_d N_A_M1017_g A_110_617# N_VDD_M1005_b PHIGHVT L=0.15 W=3
+ AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=5.5751 M=1 R=20 SA=75000.6
+ SB=75003.6 A=0.45 P=6.3 MULT=1
MM1002 N_VDD_M1017_d N_A_27_617#_M1002_g N_Y_M1002_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001
+ SB=75003.2 A=0.45 P=6.3 MULT=1
MM1003 N_VDD_M1003_d N_A_27_617#_M1003_g N_Y_M1002_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.5
+ SB=75002.8 A=0.45 P=6.3 MULT=1
MM1004 N_VDD_M1003_d N_A_27_617#_M1004_g N_Y_M1004_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.9
+ SB=75002.3 A=0.45 P=6.3 MULT=1
MM1008 N_VDD_M1008_d N_A_27_617#_M1008_g N_Y_M1004_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.3
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1009 N_VDD_M1008_d N_A_27_617#_M1009_g N_Y_M1009_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75002.8
+ SB=75001.5 A=0.45 P=6.3 MULT=1
MM1011 N_VDD_M1011_d N_A_27_617#_M1011_g N_Y_M1009_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.2
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1014 N_VDD_M1011_d N_A_27_617#_M1014_g N_Y_M1014_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75003.6
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1019 N_VDD_M1019_d N_A_27_617#_M1019_g N_Y_M1014_s N_VDD_M1005_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75004.1
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX20_noxref N_GND_M1006_b N_VDD_M1005_b NWDIODE A=18.981 P=17.59
pX21_noxref noxref_8 B B PROBETYPE=1
pX22_noxref noxref_9 A A PROBETYPE=1
pX23_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ls__or2_8.pxi.spice"
*
.ends
*
*
