* File: sky130_osu_sc_12T_ls__aoi21_l.pxi.spice
* Created: Fri Nov 12 15:34:40 2021
* 
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%GND N_GND_M1003_s N_GND_M1004_d N_GND_M1003_b
+ N_GND_c_3_p N_GND_c_4_p N_GND_c_21_p GND N_GND_c_5_p
+ PM_SKY130_OSU_SC_12T_LS__AOI21_L%GND
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_47_p
+ N_VDD_c_48_p N_VDD_c_53_p VDD N_VDD_c_49_p
+ PM_SKY130_OSU_SC_12T_LS__AOI21_L%VDD
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%A0 N_A0_c_72_n N_A0_c_73_n N_A0_M1003_g
+ N_A0_M1001_g N_A0_c_77_n N_A0_c_79_n N_A0_c_80_n A0
+ PM_SKY130_OSU_SC_12T_LS__AOI21_L%A0
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%A1 N_A1_M1000_g N_A1_M1005_g N_A1_c_110_n
+ N_A1_c_111_n N_A1_c_112_n A1 PM_SKY130_OSU_SC_12T_LS__AOI21_L%A1
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%B0 N_B0_M1004_g N_B0_c_170_n N_B0_M1002_g
+ N_B0_c_161_n N_B0_c_162_n N_B0_c_163_n N_B0_c_165_n N_B0_c_166_n N_B0_c_167_n
+ B0 PM_SKY130_OSU_SC_12T_LS__AOI21_L%B0
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%A_27_521# N_A_27_521#_M1001_s
+ N_A_27_521#_M1005_d N_A_27_521#_c_212_n N_A_27_521#_c_215_n
+ N_A_27_521#_c_222_n N_A_27_521#_c_217_n
+ PM_SKY130_OSU_SC_12T_LS__AOI21_L%A_27_521#
x_PM_SKY130_OSU_SC_12T_LS__AOI21_L%Y N_Y_M1000_d N_Y_M1002_d N_Y_c_227_n
+ N_Y_c_230_n N_Y_c_231_n Y N_Y_c_236_n N_Y_c_240_n
+ PM_SKY130_OSU_SC_12T_LS__AOI21_L%Y
cc_1 N_GND_M1003_b N_A0_c_72_n 0.0653521f $X=-0.05 $Y=0 $X2=0.295 $Y2=2.15
cc_2 N_GND_M1003_b N_A0_c_73_n 0.0202714f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.21
cc_3 N_GND_c_3_p N_A0_c_73_n 0.00502587f $X=0.26 $Y=0.735 $X2=0.475 $Y2=1.21
cc_4 N_GND_c_4_p N_A0_c_73_n 0.00606f $X=1.455 $Y=0.15 $X2=0.475 $Y2=1.21
cc_5 N_GND_c_5_p N_A0_c_73_n 0.00467791f $X=1.02 $Y=0.185 $X2=0.475 $Y2=1.21
cc_6 N_GND_M1003_b N_A0_c_77_n 0.0299759f $X=-0.05 $Y=0 $X2=0.475 $Y2=1.29
cc_7 N_GND_c_3_p N_A0_c_77_n 0.00531179f $X=0.26 $Y=0.735 $X2=0.475 $Y2=1.29
cc_8 N_GND_M1003_b N_A0_c_79_n 0.0395437f $X=-0.05 $Y=0 $X2=0.475 $Y2=2.285
cc_9 N_GND_M1003_b N_A0_c_80_n 0.0018756f $X=-0.05 $Y=0 $X2=0.385 $Y2=2.11
cc_10 N_GND_M1003_b A0 0.00934615f $X=-0.05 $Y=0 $X2=0.385 $Y2=2.11
cc_11 N_GND_M1003_b N_A1_M1000_g 0.0410177f $X=-0.05 $Y=0 $X2=0.835 $Y2=0.83
cc_12 N_GND_c_4_p N_A1_M1000_g 0.00606f $X=1.455 $Y=0.15 $X2=0.835 $Y2=0.83
cc_13 N_GND_c_5_p N_A1_M1000_g 0.00467791f $X=1.02 $Y=0.185 $X2=0.835 $Y2=0.83
cc_14 N_GND_M1003_b N_A1_M1005_g 0.0278255f $X=-0.05 $Y=0 $X2=0.905 $Y2=3.235
cc_15 N_GND_M1003_b N_A1_c_110_n 0.0355292f $X=-0.05 $Y=0 $X2=0.815 $Y2=1.775
cc_16 N_GND_M1003_b N_A1_c_111_n 0.00802017f $X=-0.05 $Y=0 $X2=0.725 $Y2=2.48
cc_17 N_GND_M1003_b N_A1_c_112_n 0.00478352f $X=-0.05 $Y=0 $X2=0.815 $Y2=1.775
cc_18 N_GND_M1003_b A1 0.00144495f $X=-0.05 $Y=0 $X2=0.725 $Y2=2.48
cc_19 N_GND_M1003_b N_B0_M1004_g 0.0307266f $X=-0.05 $Y=0 $X2=1.325 $Y2=0.75
cc_20 N_GND_c_4_p N_B0_M1004_g 0.00606f $X=1.455 $Y=0.15 $X2=1.325 $Y2=0.75
cc_21 N_GND_c_21_p N_B0_M1004_g 0.00502587f $X=1.54 $Y=0.735 $X2=1.325 $Y2=0.75
cc_22 N_GND_c_5_p N_B0_M1004_g 0.0046779f $X=1.02 $Y=0.185 $X2=1.325 $Y2=0.75
cc_23 N_GND_M1003_b N_B0_c_161_n 0.0564218f $X=-0.05 $Y=0 $X2=1.47 $Y2=2.37
cc_24 N_GND_M1003_b N_B0_c_162_n 0.0109551f $X=-0.05 $Y=0 $X2=1.47 $Y2=2.445
cc_25 N_GND_M1003_b N_B0_c_163_n 0.0497584f $X=-0.05 $Y=0 $X2=1.47 $Y2=1.38
cc_26 N_GND_c_21_p N_B0_c_163_n 0.00293502f $X=1.54 $Y=0.735 $X2=1.47 $Y2=1.38
cc_27 N_GND_M1003_b N_B0_c_165_n 0.0141127f $X=-0.05 $Y=0 $X2=1.165 $Y2=2.11
cc_28 N_GND_M1003_b N_B0_c_166_n 0.00388118f $X=-0.05 $Y=0 $X2=1.25 $Y2=1.38
cc_29 N_GND_M1003_b N_B0_c_167_n 0.011995f $X=-0.05 $Y=0 $X2=1.53 $Y2=1.38
cc_30 N_GND_c_21_p N_B0_c_167_n 0.00383173f $X=1.54 $Y=0.735 $X2=1.53 $Y2=1.38
cc_31 N_GND_M1003_b B0 0.0175171f $X=-0.05 $Y=0 $X2=1.165 $Y2=2.11
cc_32 N_GND_M1003_b N_Y_c_227_n 0.00322987f $X=-0.05 $Y=0 $X2=1.05 $Y2=0.735
cc_33 N_GND_c_4_p N_Y_c_227_n 0.00721589f $X=1.455 $Y=0.15 $X2=1.05 $Y2=0.735
cc_34 N_GND_c_5_p N_Y_c_227_n 0.0047087f $X=1.02 $Y=0.185 $X2=1.05 $Y2=0.735
cc_35 N_GND_M1003_b N_Y_c_230_n 0.0224787f $X=-0.05 $Y=0 $X2=1.55 $Y2=1.74
cc_36 N_GND_M1004_d N_Y_c_231_n 0.00291716f $X=1.4 $Y=0.57 $X2=1.465 $Y2=1.002
cc_37 N_GND_M1003_b N_Y_c_231_n 0.00762392f $X=-0.05 $Y=0 $X2=1.465 $Y2=1.002
cc_38 N_GND_c_4_p N_Y_c_231_n 0.00464239f $X=1.455 $Y=0.15 $X2=1.465 $Y2=1.002
cc_39 N_GND_c_21_p N_Y_c_231_n 0.00771134f $X=1.54 $Y=0.735 $X2=1.465 $Y2=1.002
cc_40 N_GND_M1003_b Y 0.00901344f $X=-0.05 $Y=0 $X2=1.55 $Y2=1.59
cc_41 N_GND_M1003_b N_Y_c_236_n 0.00559119f $X=-0.05 $Y=0 $X2=1.165 $Y2=1
cc_42 N_GND_c_3_p N_Y_c_236_n 8.83982e-19 $X=0.26 $Y=0.735 $X2=1.165 $Y2=1
cc_43 N_GND_c_4_p N_Y_c_236_n 0.00199024f $X=1.455 $Y=0.15 $X2=1.165 $Y2=1
cc_44 N_GND_c_21_p N_Y_c_236_n 3.97553e-19 $X=1.54 $Y=0.735 $X2=1.165 $Y2=1
cc_45 N_GND_M1003_b N_Y_c_240_n 0.0114144f $X=-0.05 $Y=0 $X2=1.55 $Y2=1.74
cc_46 N_VDD_M1001_b N_A0_M1001_g 0.0287852f $X=-0.05 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_47 N_VDD_c_47_p N_A0_M1001_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475
+ $Y2=3.235
cc_48 N_VDD_c_48_p N_A0_M1001_g 0.00339848f $X=0.69 $Y=3.63 $X2=0.475 $Y2=3.235
cc_49 N_VDD_c_49_p N_A0_M1001_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.235
cc_50 N_VDD_M1001_b N_A0_c_80_n 0.0024763f $X=-0.05 $Y=2.425 $X2=0.385 $Y2=2.11
cc_51 N_VDD_M1001_b N_A1_M1005_g 0.0189812f $X=-0.05 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_52 N_VDD_c_48_p N_A1_M1005_g 0.00339848f $X=0.69 $Y=3.63 $X2=0.905 $Y2=3.235
cc_53 N_VDD_c_53_p N_A1_M1005_g 0.00606474f $X=1.02 $Y=4.22 $X2=0.905 $Y2=3.235
cc_54 N_VDD_c_49_p N_A1_M1005_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.905 $Y2=3.235
cc_55 N_VDD_M1001_b N_A1_c_111_n 0.00500056f $X=-0.05 $Y=2.425 $X2=0.725
+ $Y2=2.48
cc_56 N_VDD_M1001_b A1 0.00652734f $X=-0.05 $Y=2.425 $X2=0.725 $Y2=2.48
cc_57 N_VDD_M1001_b N_B0_c_170_n 0.0192717f $X=-0.05 $Y=2.425 $X2=1.335 $Y2=2.52
cc_58 N_VDD_c_53_p N_B0_c_170_n 0.00606474f $X=1.02 $Y=4.22 $X2=1.335 $Y2=2.52
cc_59 N_VDD_c_49_p N_B0_c_170_n 0.00468827f $X=1.02 $Y=4.25 $X2=1.335 $Y2=2.52
cc_60 N_VDD_M1001_b N_B0_c_162_n 0.0127892f $X=-0.05 $Y=2.425 $X2=1.47 $Y2=2.445
cc_61 N_VDD_M1001_b N_A_27_521#_c_212_n 0.00156053f $X=-0.05 $Y=2.425 $X2=0.26
+ $Y2=3.63
cc_62 N_VDD_c_47_p N_A_27_521#_c_212_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=3.63
cc_63 N_VDD_c_49_p N_A_27_521#_c_212_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26
+ $Y2=3.63
cc_64 N_VDD_M1001_d N_A_27_521#_c_215_n 0.00460359f $X=0.55 $Y=2.605 $X2=1.035
+ $Y2=3.145
cc_65 N_VDD_c_48_p N_A_27_521#_c_215_n 0.0135055f $X=0.69 $Y=3.63 $X2=1.035
+ $Y2=3.145
cc_66 N_VDD_M1001_b N_A_27_521#_c_217_n 0.00155118f $X=-0.05 $Y=2.425 $X2=1.12
+ $Y2=3.635
cc_67 N_VDD_c_53_p N_A_27_521#_c_217_n 0.00734006f $X=1.02 $Y=4.22 $X2=1.12
+ $Y2=3.635
cc_68 N_VDD_c_49_p N_A_27_521#_c_217_n 0.00475776f $X=1.02 $Y=4.25 $X2=1.12
+ $Y2=3.635
cc_69 N_VDD_M1001_b N_Y_c_230_n 0.00833139f $X=-0.05 $Y=2.425 $X2=1.55 $Y2=1.74
cc_70 N_VDD_c_53_p N_Y_c_230_n 0.00757793f $X=1.02 $Y=4.22 $X2=1.55 $Y2=1.74
cc_71 N_VDD_c_49_p N_Y_c_230_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.55 $Y2=1.74
cc_72 N_A0_c_72_n N_A1_M1000_g 0.00899556f $X=0.295 $Y=2.15 $X2=0.835 $Y2=0.83
cc_73 N_A0_c_73_n N_A1_M1000_g 0.0577959f $X=0.475 $Y=1.21 $X2=0.835 $Y2=0.83
cc_74 N_A0_c_72_n N_A1_M1005_g 0.00400739f $X=0.295 $Y=2.15 $X2=0.905 $Y2=3.235
cc_75 N_A0_c_79_n N_A1_M1005_g 0.063953f $X=0.475 $Y=2.285 $X2=0.905 $Y2=3.235
cc_76 N_A0_c_72_n N_A1_c_110_n 0.0125472f $X=0.295 $Y=2.15 $X2=0.815 $Y2=1.775
cc_77 N_A0_c_72_n N_A1_c_111_n 0.00200886f $X=0.295 $Y=2.15 $X2=0.725 $Y2=2.48
cc_78 N_A0_c_79_n N_A1_c_111_n 0.00432627f $X=0.475 $Y=2.285 $X2=0.725 $Y2=2.48
cc_79 N_A0_c_80_n N_A1_c_111_n 0.0279489f $X=0.385 $Y=2.11 $X2=0.725 $Y2=2.48
cc_80 A0 N_A1_c_111_n 0.00329388f $X=0.385 $Y=2.11 $X2=0.725 $Y2=2.48
cc_81 N_A0_c_72_n N_A1_c_112_n 0.00661569f $X=0.295 $Y=2.15 $X2=0.815 $Y2=1.775
cc_82 N_A0_c_79_n A1 0.00417236f $X=0.475 $Y=2.285 $X2=0.725 $Y2=2.48
cc_83 N_A0_c_80_n A1 0.00265232f $X=0.385 $Y=2.11 $X2=0.725 $Y2=2.48
cc_84 A0 A1 0.00563601f $X=0.385 $Y=2.11 $X2=0.725 $Y2=2.48
cc_85 A0 B0 0.0169035f $X=0.385 $Y=2.11 $X2=1.165 $Y2=2.11
cc_86 N_A0_M1001_g N_A_27_521#_c_215_n 0.0196156f $X=0.475 $Y=3.235 $X2=1.035
+ $Y2=3.145
cc_87 N_A0_c_80_n N_A_27_521#_c_215_n 0.00272894f $X=0.385 $Y=2.11 $X2=1.035
+ $Y2=3.145
cc_88 N_A0_c_79_n N_A_27_521#_c_222_n 0.00266419f $X=0.475 $Y=2.285 $X2=0.345
+ $Y2=3.145
cc_89 N_A0_c_80_n N_A_27_521#_c_222_n 0.00150818f $X=0.385 $Y=2.11 $X2=0.345
+ $Y2=3.145
cc_90 N_A0_c_73_n N_Y_c_236_n 0.00104705f $X=0.475 $Y=1.21 $X2=1.165 $Y2=1
cc_91 N_A1_M1000_g N_B0_M1004_g 0.0273492f $X=0.835 $Y=0.83 $X2=1.325 $Y2=0.75
cc_92 N_A1_c_110_n N_B0_c_161_n 0.0174043f $X=0.815 $Y=1.775 $X2=1.47 $Y2=2.37
cc_93 N_A1_M1005_g N_B0_c_162_n 0.0533932f $X=0.905 $Y=3.235 $X2=1.47 $Y2=2.445
cc_94 A1 N_B0_c_162_n 0.00107545f $X=0.725 $Y=2.48 $X2=1.47 $Y2=2.445
cc_95 N_A1_M1000_g N_B0_c_163_n 0.0039494f $X=0.835 $Y=0.83 $X2=1.47 $Y2=1.38
cc_96 N_A1_M1000_g N_B0_c_165_n 0.00326852f $X=0.835 $Y=0.83 $X2=1.165 $Y2=2.11
cc_97 N_A1_c_110_n N_B0_c_165_n 0.00506769f $X=0.815 $Y=1.775 $X2=1.165 $Y2=2.11
cc_98 N_A1_c_111_n N_B0_c_165_n 0.0109205f $X=0.725 $Y=2.48 $X2=1.165 $Y2=2.11
cc_99 N_A1_c_112_n N_B0_c_165_n 0.0226306f $X=0.815 $Y=1.775 $X2=1.165 $Y2=2.11
cc_100 N_A1_M1000_g N_B0_c_166_n 0.00477017f $X=0.835 $Y=0.83 $X2=1.25 $Y2=1.38
cc_101 N_A1_M1005_g B0 0.00588076f $X=0.905 $Y=3.235 $X2=1.165 $Y2=2.11
cc_102 N_A1_c_111_n B0 0.00258971f $X=0.725 $Y=2.48 $X2=1.165 $Y2=2.11
cc_103 A1 B0 0.00582284f $X=0.725 $Y=2.48 $X2=1.165 $Y2=2.11
cc_104 N_A1_M1005_g N_A_27_521#_c_215_n 0.0157671f $X=0.905 $Y=3.235 $X2=1.035
+ $Y2=3.145
cc_105 N_A1_c_111_n N_A_27_521#_c_215_n 0.00325705f $X=0.725 $Y=2.48 $X2=1.035
+ $Y2=3.145
cc_106 A1 N_A_27_521#_c_215_n 0.0109287f $X=0.725 $Y=2.48 $X2=1.035 $Y2=3.145
cc_107 N_A1_M1000_g N_Y_c_227_n 0.00218184f $X=0.835 $Y=0.83 $X2=1.05 $Y2=0.735
cc_108 N_A1_c_110_n N_Y_c_227_n 3.5348e-19 $X=0.815 $Y=1.775 $X2=1.05 $Y2=0.735
cc_109 N_A1_M1005_g N_Y_c_230_n 0.00114141f $X=0.905 $Y=3.235 $X2=1.55 $Y2=1.74
cc_110 N_A1_c_111_n N_Y_c_230_n 0.00648983f $X=0.725 $Y=2.48 $X2=1.55 $Y2=1.74
cc_111 A1 N_Y_c_230_n 0.00498789f $X=0.725 $Y=2.48 $X2=1.55 $Y2=1.74
cc_112 N_A1_M1000_g Y 3.27704e-19 $X=0.835 $Y=0.83 $X2=1.55 $Y2=1.59
cc_113 N_A1_M1000_g N_Y_c_236_n 0.00542417f $X=0.835 $Y=0.83 $X2=1.165 $Y2=1
cc_114 N_A1_c_110_n N_Y_c_236_n 0.00171207f $X=0.815 $Y=1.775 $X2=1.165 $Y2=1
cc_115 N_B0_M1004_g N_Y_c_227_n 0.00643266f $X=1.325 $Y=0.75 $X2=1.05 $Y2=0.735
cc_116 N_B0_c_166_n N_Y_c_227_n 0.00325506f $X=1.25 $Y=1.38 $X2=1.05 $Y2=0.735
cc_117 N_B0_c_170_n N_Y_c_230_n 0.0129182f $X=1.335 $Y=2.52 $X2=1.55 $Y2=1.74
cc_118 N_B0_c_161_n N_Y_c_230_n 0.0233833f $X=1.47 $Y=2.37 $X2=1.55 $Y2=1.74
cc_119 N_B0_c_162_n N_Y_c_230_n 0.00827561f $X=1.47 $Y=2.445 $X2=1.55 $Y2=1.74
cc_120 N_B0_c_163_n N_Y_c_230_n 0.00170788f $X=1.47 $Y=1.38 $X2=1.55 $Y2=1.74
cc_121 N_B0_c_165_n N_Y_c_230_n 0.027719f $X=1.165 $Y=2.11 $X2=1.55 $Y2=1.74
cc_122 N_B0_c_167_n N_Y_c_230_n 0.0101032f $X=1.53 $Y=1.38 $X2=1.55 $Y2=1.74
cc_123 B0 N_Y_c_230_n 0.00715529f $X=1.165 $Y=2.11 $X2=1.55 $Y2=1.74
cc_124 N_B0_M1004_g N_Y_c_231_n 0.00766738f $X=1.325 $Y=0.75 $X2=1.465 $Y2=1.002
cc_125 N_B0_c_163_n N_Y_c_231_n 0.00146003f $X=1.47 $Y=1.38 $X2=1.465 $Y2=1.002
cc_126 N_B0_c_166_n N_Y_c_231_n 0.00438276f $X=1.25 $Y=1.38 $X2=1.465 $Y2=1.002
cc_127 N_B0_c_167_n N_Y_c_231_n 0.00722649f $X=1.53 $Y=1.38 $X2=1.465 $Y2=1.002
cc_128 N_B0_M1004_g Y 0.00266245f $X=1.325 $Y=0.75 $X2=1.55 $Y2=1.59
cc_129 N_B0_c_161_n Y 0.00138242f $X=1.47 $Y=2.37 $X2=1.55 $Y2=1.59
cc_130 N_B0_c_163_n Y 0.01116f $X=1.47 $Y=1.38 $X2=1.55 $Y2=1.59
cc_131 N_B0_c_165_n Y 0.00642461f $X=1.165 $Y=2.11 $X2=1.55 $Y2=1.59
cc_132 N_B0_c_167_n Y 0.0195669f $X=1.53 $Y=1.38 $X2=1.55 $Y2=1.59
cc_133 N_B0_M1004_g N_Y_c_236_n 6.32765e-19 $X=1.325 $Y=0.75 $X2=1.165 $Y2=1
cc_134 N_B0_c_166_n N_Y_c_236_n 0.00324068f $X=1.25 $Y=1.38 $X2=1.165 $Y2=1
cc_135 N_B0_c_161_n N_Y_c_240_n 0.00516977f $X=1.47 $Y=2.37 $X2=1.55 $Y2=1.74
cc_136 N_B0_c_163_n N_Y_c_240_n 8.18646e-19 $X=1.47 $Y=1.38 $X2=1.55 $Y2=1.74
cc_137 N_B0_c_165_n N_Y_c_240_n 0.00655582f $X=1.165 $Y=2.11 $X2=1.55 $Y2=1.74
cc_138 N_B0_c_167_n N_Y_c_240_n 0.00438887f $X=1.53 $Y=1.38 $X2=1.55 $Y2=1.74
