* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_osu_sc_18T_ms__nor2_l
** N=9 EP=0 IP=0 FDC=8
M0 Y B gnd gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=400 $Y=575 $D=9
M1 gnd A Y gnd nshort L=0.15 W=0.74 m=1 r=4.93333 a=0.111 p=1.78 mult=1 $X=830 $Y=575 $D=9
M2 6 B Y vdd pshort L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=400 $Y=4085 $D=79
M3 vdd A 6 vdd pshort L=0.15 W=2 m=1 r=13.3333 a=0.3 p=4.3 mult=1 $X=760 $Y=4085 $D=79
X4 gnd vdd Dpar a=5.605 p=10.55 m=1 $[nwdiode] $X=-45 $Y=2905 $D=185
X5 7 B Probe probetype=1 $[B] $X=648 $Y=2958 $D=289
X6 8 Y Probe probetype=1 $[Y] $X=683 $Y=1963 $D=289
X7 9 A Probe probetype=1 $[A] $X=988 $Y=3328 $D=289
.ENDS
***************************************
