magic
tech sky130A
magscale 1 2
timestamp 1606864601
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 374 1341
<< nmos >>
rect 80 115 110 315
rect 152 115 182 315
rect 250 115 280 263
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
rect 252 617 282 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 115 152 315
rect 182 267 235 315
rect 182 131 193 267
rect 227 263 235 267
rect 227 131 250 263
rect 182 115 250 131
rect 280 199 333 263
rect 280 131 291 199
rect 325 131 333 199
rect 280 115 333 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 166 1217
rect 110 861 121 1201
rect 155 861 166 1201
rect 110 617 166 861
rect 196 1201 252 1217
rect 196 793 207 1201
rect 241 793 252 1201
rect 196 617 252 793
rect 282 1201 335 1217
rect 282 725 293 1201
rect 327 725 335 1201
rect 282 617 335 725
<< ndiffc >>
rect 35 131 69 267
rect 193 131 227 267
rect 291 131 325 199
<< pdiffc >>
rect 35 793 69 1201
rect 121 861 155 1201
rect 207 793 241 1201
rect 293 725 327 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 252 1217 282 1243
rect 80 580 110 617
rect 44 570 110 580
rect 44 536 60 570
rect 94 536 110 570
rect 44 526 110 536
rect 44 370 74 526
rect 166 484 196 617
rect 252 579 282 617
rect 252 549 309 579
rect 134 468 196 484
rect 134 434 146 468
rect 180 434 196 468
rect 134 418 196 434
rect 44 338 110 370
rect 80 315 110 338
rect 152 315 182 418
rect 279 405 309 549
rect 279 389 333 405
rect 279 371 289 389
rect 250 355 289 371
rect 323 355 333 389
rect 250 339 333 355
rect 250 263 280 339
rect 80 89 110 115
rect 152 89 182 115
rect 250 89 280 115
<< polycont >>
rect 60 536 94 570
rect 146 434 180 468
rect 289 355 323 389
<< locali >>
rect 0 1311 374 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 374 1311
rect 35 1201 69 1217
rect 121 1201 155 1271
rect 121 845 155 861
rect 207 1201 241 1217
rect 69 793 207 811
rect 35 777 241 793
rect 293 1201 327 1217
rect 60 570 94 649
rect 60 520 94 536
rect 128 484 162 575
rect 128 468 180 484
rect 128 434 146 468
rect 128 418 180 434
rect 216 389 250 501
rect 293 461 327 725
rect 216 355 289 389
rect 323 355 339 389
rect 35 267 69 283
rect 35 61 69 131
rect 193 267 227 279
rect 193 115 227 131
rect 291 199 325 215
rect 291 61 325 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 60 649 94 683
rect 128 575 162 609
rect 216 501 250 535
rect 293 427 327 461
rect 193 279 227 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 374 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 374 1311
rect 0 1271 374 1277
rect 48 683 106 689
rect 48 649 60 683
rect 94 649 128 683
rect 48 643 106 649
rect 116 609 174 615
rect 116 575 128 609
rect 162 575 196 609
rect 116 569 174 575
rect 204 535 262 541
rect 182 501 216 535
rect 250 501 262 535
rect 204 495 262 501
rect 281 461 339 467
rect 281 427 293 461
rect 327 427 339 461
rect 281 421 339 427
rect 181 313 239 319
rect 293 313 327 421
rect 181 279 193 313
rect 227 279 327 313
rect 181 273 239 279
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 77 666 77 666 1 A0
port 1 n
rlabel metal1 233 518 233 518 1 B0
port 2 n
rlabel metal1 310 414 310 414 1 Y
port 3 n
rlabel metal1 145 592 145 592 1 A1
port 4 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
