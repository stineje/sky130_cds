* File: sky130_osu_sc_15T_ls__dlat_l.pxi.spice
* Created: Fri Nov 12 14:56:50 2021
* 
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%GND N_GND_M1001_s N_GND_M1004_d N_GND_M1007_s
+ N_GND_M1008_d N_GND_M1001_b N_GND_c_4_p N_GND_c_5_p N_GND_c_25_p N_GND_c_39_p
+ N_GND_c_9_p N_GND_c_10_p N_GND_c_76_p GND N_GND_c_6_p
+ PM_SKY130_OSU_SC_15T_LS__DLAT_L%GND
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%VDD N_VDD_M1009_s N_VDD_M1012_d N_VDD_M1014_s
+ N_VDD_M1005_d N_VDD_M1009_b N_VDD_c_116_p N_VDD_c_117_p N_VDD_c_132_p
+ N_VDD_c_133_p N_VDD_c_120_p N_VDD_c_121_p N_VDD_c_155_p N_VDD_c_163_p VDD
+ N_VDD_c_118_p PM_SKY130_OSU_SC_15T_LS__DLAT_L%VDD
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%D N_D_M1015_d N_D_M1003_d N_D_c_175_n
+ N_D_c_176_n N_D_M1001_g N_D_M1009_g N_D_c_182_n N_D_M1007_g N_D_M1014_g
+ N_D_c_187_n N_D_c_188_n N_D_c_190_n N_D_c_191_n N_D_c_219_p N_D_c_293_p
+ N_D_c_225_p N_D_c_290_p N_D_c_192_n N_D_c_213_n N_D_c_195_n N_D_c_197_n
+ N_D_c_198_n N_D_c_200_n D N_D_c_202_n PM_SKY130_OSU_SC_15T_LS__DLAT_L%D
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%CK N_CK_M1015_g N_CK_M1010_g N_CK_M1006_g
+ N_CK_c_294_n N_CK_M1002_g N_CK_c_295_n N_CK_c_296_n N_CK_c_297_n N_CK_c_300_n
+ N_CK_c_301_n N_CK_c_306_n N_CK_c_307_n N_CK_c_308_n N_CK_c_309_n N_CK_c_310_n
+ N_CK_c_311_n N_CK_c_312_n N_CK_c_313_n CK PM_SKY130_OSU_SC_15T_LS__DLAT_L%CK
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%A_157_393# N_A_157_393#_M1006_d
+ N_A_157_393#_M1002_d N_A_157_393#_M1003_g N_A_157_393#_c_428_n
+ N_A_157_393#_c_429_n N_A_157_393#_c_430_n N_A_157_393#_M1013_g
+ N_A_157_393#_c_431_n N_A_157_393#_c_432_n N_A_157_393#_c_435_n
+ N_A_157_393#_c_437_n N_A_157_393#_c_441_n N_A_157_393#_c_448_n
+ N_A_157_393#_c_442_n N_A_157_393#_c_443_n N_A_157_393#_c_444_n
+ N_A_157_393#_c_453_n PM_SKY130_OSU_SC_15T_LS__DLAT_L%A_157_393#
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%A_349_89# N_A_349_89#_M1007_d
+ N_A_349_89#_M1014_d N_A_349_89#_M1004_g N_A_349_89#_M1012_g
+ N_A_349_89#_M1008_g N_A_349_89#_M1005_g N_A_349_89#_c_555_n
+ N_A_349_89#_c_556_n N_A_349_89#_c_557_n N_A_349_89#_c_558_n
+ N_A_349_89#_c_559_n N_A_349_89#_c_560_n N_A_349_89#_c_561_n
+ N_A_349_89#_c_562_n N_A_349_89#_c_565_n N_A_349_89#_c_566_n
+ N_A_349_89#_c_567_n N_A_349_89#_c_568_n N_A_349_89#_c_569_n
+ N_A_349_89#_c_570_n PM_SKY130_OSU_SC_15T_LS__DLAT_L%A_349_89#
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%QN N_QN_M1008_s N_QN_M1005_s N_QN_M1011_g
+ N_QN_M1000_g N_QN_c_684_n N_QN_c_685_n N_QN_c_688_n N_QN_c_689_n N_QN_c_691_n
+ N_QN_c_692_n N_QN_c_693_n N_QN_c_694_n QN PM_SKY130_OSU_SC_15T_LS__DLAT_L%QN
x_PM_SKY130_OSU_SC_15T_LS__DLAT_L%Q N_Q_M1011_d N_Q_M1000_d N_Q_c_757_n
+ N_Q_c_762_n N_Q_c_763_n N_Q_c_759_n N_Q_c_761_n Q
+ PM_SKY130_OSU_SC_15T_LS__DLAT_L%Q
cc_1 N_GND_M1001_b N_D_c_175_n 0.0193486f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.88
cc_2 N_GND_M1001_b N_D_c_176_n 0.0111643f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.96
cc_3 N_GND_M1001_b N_D_M1001_g 0.0422121f $X=-0.045 $Y=0 $X2=0.5 $Y2=0.945
cc_4 N_GND_c_4_p N_D_M1001_g 0.00502587f $X=0.285 $Y=0.74 $X2=0.5 $Y2=0.945
cc_5 N_GND_c_5_p N_D_M1001_g 0.00606474f $X=1.95 $Y=0.152 $X2=0.5 $Y2=0.945
cc_6 N_GND_c_6_p N_D_M1001_g 0.00468827f $X=4.42 $Y=0.19 $X2=0.5 $Y2=0.945
cc_7 N_GND_M1001_b N_D_M1009_g 0.035797f $X=-0.045 $Y=0 $X2=0.5 $Y2=3.825
cc_8 N_GND_M1001_b N_D_c_182_n 0.0221119f $X=-0.045 $Y=0 $X2=3.2 $Y2=1.425
cc_9 N_GND_c_9_p N_D_c_182_n 0.00866533f $X=2.985 $Y=0.825 $X2=3.2 $Y2=1.425
cc_10 N_GND_c_10_p N_D_c_182_n 0.00606474f $X=4.28 $Y=0.152 $X2=3.2 $Y2=1.425
cc_11 N_GND_c_6_p N_D_c_182_n 0.00468827f $X=4.42 $Y=0.19 $X2=3.2 $Y2=1.425
cc_12 N_GND_M1001_b N_D_M1014_g 0.0594514f $X=-0.045 $Y=0 $X2=3.2 $Y2=3.825
cc_13 N_GND_M1001_b N_D_c_187_n 0.0173576f $X=-0.045 $Y=0 $X2=0.44 $Y2=2.155
cc_14 N_GND_M1001_b N_D_c_188_n 0.0482669f $X=-0.045 $Y=0 $X2=3.2 $Y2=1.59
cc_15 N_GND_c_9_p N_D_c_188_n 0.00386381f $X=2.985 $Y=0.825 $X2=3.2 $Y2=1.59
cc_16 N_GND_M1001_b N_D_c_190_n 0.00268454f $X=-0.045 $Y=0 $X2=0.58 $Y2=1.59
cc_17 N_GND_M1001_b N_D_c_191_n 0.00380459f $X=-0.045 $Y=0 $X2=0.58 $Y2=2.84
cc_18 N_GND_M1001_b N_D_c_192_n 0.00313975f $X=-0.045 $Y=0 $X2=1.16 $Y2=0.825
cc_19 N_GND_c_5_p N_D_c_192_n 0.0149461f $X=1.95 $Y=0.152 $X2=1.16 $Y2=0.825
cc_20 N_GND_c_6_p N_D_c_192_n 0.00958198f $X=4.42 $Y=0.19 $X2=1.16 $Y2=0.825
cc_21 N_GND_M1001_b N_D_c_195_n 0.00161958f $X=-0.045 $Y=0 $X2=2.995 $Y2=1.59
cc_22 N_GND_c_9_p N_D_c_195_n 0.00509685f $X=2.985 $Y=0.825 $X2=2.995 $Y2=1.59
cc_23 N_GND_M1001_b N_D_c_197_n 0.00166426f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.96
cc_24 N_GND_M1001_b N_D_c_198_n 0.0405753f $X=-0.045 $Y=0 $X2=2.85 $Y2=1.59
cc_25 N_GND_c_25_p N_D_c_198_n 0.00414959f $X=2.035 $Y=0.825 $X2=2.85 $Y2=1.59
cc_26 N_GND_M1001_b N_D_c_200_n 0.00214607f $X=-0.045 $Y=0 $X2=0.725 $Y2=1.59
cc_27 N_GND_M1001_b D 0.0122313f $X=-0.045 $Y=0 $X2=0.44 $Y2=1.96
cc_28 N_GND_M1001_b N_D_c_202_n 9.64388e-19 $X=-0.045 $Y=0 $X2=2.995 $Y2=1.59
cc_29 N_GND_c_9_p N_D_c_202_n 0.00387325f $X=2.985 $Y=0.825 $X2=2.995 $Y2=1.59
cc_30 N_GND_M1001_b N_CK_c_294_n 0.0311248f $X=-0.045 $Y=0 $X2=2.25 $Y2=2.67
cc_31 N_GND_M1001_b N_CK_c_295_n 0.0438842f $X=-0.045 $Y=0 $X2=2.305 $Y2=2.34
cc_32 N_GND_M1001_b N_CK_c_296_n 0.0250297f $X=-0.045 $Y=0 $X2=0.92 $Y2=1.59
cc_33 N_GND_M1001_b N_CK_c_297_n 0.0175305f $X=-0.045 $Y=0 $X2=0.92 $Y2=1.425
cc_34 N_GND_c_5_p N_CK_c_297_n 0.00606474f $X=1.95 $Y=0.152 $X2=0.92 $Y2=1.425
cc_35 N_GND_c_6_p N_CK_c_297_n 0.00468827f $X=4.42 $Y=0.19 $X2=0.92 $Y2=1.425
cc_36 N_GND_M1001_b N_CK_c_300_n 0.0233984f $X=-0.045 $Y=0 $X2=1.4 $Y2=2.505
cc_37 N_GND_M1001_b N_CK_c_301_n 0.0183851f $X=-0.045 $Y=0 $X2=2.277 $Y2=1.425
cc_38 N_GND_c_25_p N_CK_c_301_n 0.00388248f $X=2.035 $Y=0.825 $X2=2.277
+ $Y2=1.425
cc_39 N_GND_c_39_p N_CK_c_301_n 0.00606474f $X=2.9 $Y=0.152 $X2=2.277 $Y2=1.425
cc_40 N_GND_c_9_p N_CK_c_301_n 0.0041071f $X=2.985 $Y=0.825 $X2=2.277 $Y2=1.425
cc_41 N_GND_c_6_p N_CK_c_301_n 0.00468827f $X=4.42 $Y=0.19 $X2=2.277 $Y2=1.425
cc_42 N_GND_M1001_b N_CK_c_306_n 0.01373f $X=-0.045 $Y=0 $X2=2.277 $Y2=1.575
cc_43 N_GND_M1001_b N_CK_c_307_n 0.0077706f $X=-0.045 $Y=0 $X2=0.92 $Y2=1.59
cc_44 N_GND_M1001_b N_CK_c_308_n 0.00513137f $X=-0.045 $Y=0 $X2=1.315 $Y2=2.33
cc_45 N_GND_M1001_b N_CK_c_309_n 9.63154e-19 $X=-0.045 $Y=0 $X2=1.005 $Y2=2.33
cc_46 N_GND_M1001_b N_CK_c_310_n 7.61111e-19 $X=-0.045 $Y=0 $X2=2.395 $Y2=2.33
cc_47 N_GND_M1001_b N_CK_c_311_n 0.00265612f $X=-0.045 $Y=0 $X2=1.4 $Y2=2.33
cc_48 N_GND_M1001_b N_CK_c_312_n 0.0181831f $X=-0.045 $Y=0 $X2=2.25 $Y2=2.33
cc_49 N_GND_M1001_b N_CK_c_313_n 0.0041728f $X=-0.045 $Y=0 $X2=1.545 $Y2=2.33
cc_50 N_GND_M1001_b CK 0.00239232f $X=-0.045 $Y=0 $X2=2.395 $Y2=2.33
cc_51 N_GND_M1001_b N_A_157_393#_M1003_g 0.0292909f $X=-0.045 $Y=0 $X2=0.86
+ $Y2=3.825
cc_52 N_GND_M1001_b N_A_157_393#_c_428_n 0.0294293f $X=-0.045 $Y=0 $X2=1.265
+ $Y2=2.04
cc_53 N_GND_M1001_b N_A_157_393#_c_429_n 0.00679315f $X=-0.045 $Y=0 $X2=0.935
+ $Y2=2.04
cc_54 N_GND_M1001_b N_A_157_393#_c_430_n 0.0138829f $X=-0.045 $Y=0 $X2=1.34
+ $Y2=1.965
cc_55 N_GND_M1001_b N_A_157_393#_c_431_n 0.0265388f $X=-0.045 $Y=0 $X2=1.4
+ $Y2=1.59
cc_56 N_GND_M1001_b N_A_157_393#_c_432_n 0.01755f $X=-0.045 $Y=0 $X2=1.4
+ $Y2=1.425
cc_57 N_GND_c_5_p N_A_157_393#_c_432_n 0.00606474f $X=1.95 $Y=0.152 $X2=1.4
+ $Y2=1.425
cc_58 N_GND_c_6_p N_A_157_393#_c_432_n 0.00468827f $X=4.42 $Y=0.19 $X2=1.4
+ $Y2=1.425
cc_59 N_GND_M1001_b N_A_157_393#_c_435_n 0.0116005f $X=-0.045 $Y=0 $X2=2.38
+ $Y2=1.59
cc_60 N_GND_c_25_p N_A_157_393#_c_435_n 0.00572623f $X=2.035 $Y=0.825 $X2=2.38
+ $Y2=1.59
cc_61 N_GND_M1001_b N_A_157_393#_c_437_n 0.00549177f $X=-0.045 $Y=0 $X2=2.465
+ $Y2=0.825
cc_62 N_GND_c_39_p N_A_157_393#_c_437_n 0.00736239f $X=2.9 $Y=0.152 $X2=2.465
+ $Y2=0.825
cc_63 N_GND_c_9_p N_A_157_393#_c_437_n 0.0247767f $X=2.985 $Y=0.825 $X2=2.465
+ $Y2=0.825
cc_64 N_GND_c_6_p N_A_157_393#_c_437_n 0.00476261f $X=4.42 $Y=0.19 $X2=2.465
+ $Y2=0.825
cc_65 N_GND_M1001_b N_A_157_393#_c_441_n 0.00324634f $X=-0.045 $Y=0 $X2=2.465
+ $Y2=1.845
cc_66 N_GND_M1001_b N_A_157_393#_c_442_n 0.0141454f $X=-0.045 $Y=0 $X2=2.735
+ $Y2=2.84
cc_67 N_GND_M1001_b N_A_157_393#_c_443_n 8.79856e-19 $X=-0.045 $Y=0 $X2=2.465
+ $Y2=1.59
cc_68 N_GND_M1001_b N_A_157_393#_c_444_n 0.0100851f $X=-0.045 $Y=0 $X2=2.735
+ $Y2=1.93
cc_69 N_GND_M1001_b N_A_349_89#_M1004_g 0.0319752f $X=-0.045 $Y=0 $X2=1.82
+ $Y2=0.945
cc_70 N_GND_c_5_p N_A_349_89#_M1004_g 0.00606474f $X=1.95 $Y=0.152 $X2=1.82
+ $Y2=0.945
cc_71 N_GND_c_25_p N_A_349_89#_M1004_g 0.00388248f $X=2.035 $Y=0.825 $X2=1.82
+ $Y2=0.945
cc_72 N_GND_c_6_p N_A_349_89#_M1004_g 0.00468827f $X=4.42 $Y=0.19 $X2=1.82
+ $Y2=0.945
cc_73 N_GND_M1001_b N_A_349_89#_M1012_g 0.0330331f $X=-0.045 $Y=0 $X2=1.82
+ $Y2=3.825
cc_74 N_GND_M1001_b N_A_349_89#_M1008_g 0.0310629f $X=-0.045 $Y=0 $X2=4.15
+ $Y2=0.835
cc_75 N_GND_c_10_p N_A_349_89#_M1008_g 0.00606474f $X=4.28 $Y=0.152 $X2=4.15
+ $Y2=0.835
cc_76 N_GND_c_76_p N_A_349_89#_M1008_g 0.00308284f $X=4.365 $Y=0.74 $X2=4.15
+ $Y2=0.835
cc_77 N_GND_c_6_p N_A_349_89#_M1008_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.15
+ $Y2=0.835
cc_78 N_GND_M1001_b N_A_349_89#_c_555_n 0.0263478f $X=-0.045 $Y=0 $X2=1.88
+ $Y2=1.93
cc_79 N_GND_M1001_b N_A_349_89#_c_556_n 0.0291536f $X=-0.045 $Y=0 $X2=4.035
+ $Y2=1.93
cc_80 N_GND_M1001_b N_A_349_89#_c_557_n 0.0138254f $X=-0.045 $Y=0 $X2=4.037
+ $Y2=1.765
cc_81 N_GND_M1001_b N_A_349_89#_c_558_n 0.0135442f $X=-0.045 $Y=0 $X2=4.125
+ $Y2=1.54
cc_82 N_GND_M1001_b N_A_349_89#_c_559_n 0.0305585f $X=-0.045 $Y=0 $X2=4.125
+ $Y2=2.595
cc_83 N_GND_M1001_b N_A_349_89#_c_560_n 0.00495879f $X=-0.045 $Y=0 $X2=4.125
+ $Y2=2.745
cc_84 N_GND_M1001_b N_A_349_89#_c_561_n 0.0039674f $X=-0.045 $Y=0 $X2=1.88
+ $Y2=1.93
cc_85 N_GND_M1001_b N_A_349_89#_c_562_n 0.0136393f $X=-0.045 $Y=0 $X2=3.415
+ $Y2=0.825
cc_86 N_GND_c_10_p N_A_349_89#_c_562_n 0.00757793f $X=4.28 $Y=0.152 $X2=3.415
+ $Y2=0.825
cc_87 N_GND_c_6_p N_A_349_89#_c_562_n 0.00476261f $X=4.42 $Y=0.19 $X2=3.415
+ $Y2=0.825
cc_88 N_GND_M1001_b N_A_349_89#_c_565_n 0.0162343f $X=-0.045 $Y=0 $X2=3.415
+ $Y2=3.205
cc_89 N_GND_M1001_b N_A_349_89#_c_566_n 0.0123965f $X=-0.045 $Y=0 $X2=4.035
+ $Y2=1.93
cc_90 N_GND_M1001_b N_A_349_89#_c_567_n 0.00241536f $X=-0.045 $Y=0 $X2=3.415
+ $Y2=1.93
cc_91 N_GND_M1001_b N_A_349_89#_c_568_n 0.0515942f $X=-0.045 $Y=0 $X2=3.89
+ $Y2=1.93
cc_92 N_GND_M1001_b N_A_349_89#_c_569_n 0.00189525f $X=-0.045 $Y=0 $X2=2.025
+ $Y2=1.93
cc_93 N_GND_M1001_b N_A_349_89#_c_570_n 0.00128332f $X=-0.045 $Y=0 $X2=4.035
+ $Y2=1.93
cc_94 N_GND_M1001_b N_QN_M1011_g 0.0683285f $X=-0.045 $Y=0 $X2=4.58 $Y2=0.835
cc_95 N_GND_c_76_p N_QN_M1011_g 0.00308284f $X=4.365 $Y=0.74 $X2=4.58 $Y2=0.835
cc_96 N_GND_c_6_p N_QN_M1011_g 0.00468827f $X=4.42 $Y=0.19 $X2=4.58 $Y2=0.835
cc_97 N_GND_M1001_b N_QN_M1000_g 0.0184175f $X=-0.045 $Y=0 $X2=4.58 $Y2=4.195
cc_98 N_GND_M1001_b N_QN_c_684_n 0.0289957f $X=-0.045 $Y=0 $X2=4.52 $Y2=2.135
cc_99 N_GND_M1001_b N_QN_c_685_n 0.0106252f $X=-0.045 $Y=0 $X2=3.935 $Y2=0.74
cc_100 N_GND_c_10_p N_QN_c_685_n 0.00745733f $X=4.28 $Y=0.152 $X2=3.935 $Y2=0.74
cc_101 N_GND_c_6_p N_QN_c_685_n 0.00476261f $X=4.42 $Y=0.19 $X2=3.935 $Y2=0.74
cc_102 N_GND_M1001_b N_QN_c_688_n 0.00102655f $X=-0.045 $Y=0 $X2=3.935 $Y2=2.7
cc_103 N_GND_M1001_b N_QN_c_689_n 0.0139574f $X=-0.045 $Y=0 $X2=4.435 $Y2=1.59
cc_104 N_GND_c_76_p N_QN_c_689_n 0.00556529f $X=4.365 $Y=0.74 $X2=4.435 $Y2=1.59
cc_105 N_GND_M1001_b N_QN_c_691_n 0.00262941f $X=-0.045 $Y=0 $X2=4.02 $Y2=1.59
cc_106 N_GND_M1001_b N_QN_c_692_n 0.0176115f $X=-0.045 $Y=0 $X2=4.435 $Y2=2.505
cc_107 N_GND_M1001_b N_QN_c_693_n 0.00318212f $X=-0.045 $Y=0 $X2=4.02 $Y2=2.505
cc_108 N_GND_M1001_b N_QN_c_694_n 0.0034889f $X=-0.045 $Y=0 $X2=4.52 $Y2=2.135
cc_109 N_GND_M1001_b QN 0.00252171f $X=-0.045 $Y=0 $X2=3.94 $Y2=2.7
cc_110 N_GND_M1001_b N_Q_c_757_n 0.00907452f $X=-0.045 $Y=0 $X2=4.795 $Y2=0.74
cc_111 N_GND_c_6_p N_Q_c_757_n 0.00474541f $X=4.42 $Y=0.19 $X2=4.795 $Y2=0.74
cc_112 N_GND_M1001_b N_Q_c_759_n 0.00819704f $X=-0.045 $Y=0 $X2=4.827 $Y2=1.08
cc_113 N_GND_c_6_p N_Q_c_759_n 0.00148124f $X=4.42 $Y=0.19 $X2=4.827 $Y2=1.08
cc_114 N_GND_M1001_b N_Q_c_761_n 0.0735742f $X=-0.045 $Y=0 $X2=4.827 $Y2=2.9
cc_115 N_VDD_M1009_b N_D_M1009_g 0.0239842f $X=-0.045 $Y=2.645 $X2=0.5 $Y2=3.825
cc_116 N_VDD_c_116_p N_D_M1009_g 0.00751602f $X=0.285 $Y=3.545 $X2=0.5 $Y2=3.825
cc_117 N_VDD_c_117_p N_D_M1009_g 0.00606474f $X=1.95 $Y=5.247 $X2=0.5 $Y2=3.825
cc_118 N_VDD_c_118_p N_D_M1009_g 0.00468827f $X=4.42 $Y=5.21 $X2=0.5 $Y2=3.825
cc_119 N_VDD_M1009_b N_D_M1014_g 0.0260072f $X=-0.045 $Y=2.645 $X2=3.2 $Y2=3.825
cc_120 N_VDD_c_120_p N_D_M1014_g 0.00751602f $X=2.985 $Y=3.545 $X2=3.2 $Y2=3.825
cc_121 N_VDD_c_121_p N_D_M1014_g 0.00606474f $X=4.28 $Y=5.247 $X2=3.2 $Y2=3.825
cc_122 N_VDD_c_118_p N_D_M1014_g 0.00468827f $X=4.42 $Y=5.21 $X2=3.2 $Y2=3.825
cc_123 N_VDD_M1009_b N_D_c_191_n 0.00168314f $X=-0.045 $Y=2.645 $X2=0.58
+ $Y2=2.84
cc_124 N_VDD_M1009_b N_D_c_213_n 0.00313975f $X=-0.045 $Y=2.645 $X2=1.16
+ $Y2=3.205
cc_125 N_VDD_c_117_p N_D_c_213_n 0.0149461f $X=1.95 $Y=5.247 $X2=1.16 $Y2=3.205
cc_126 N_VDD_c_118_p N_D_c_213_n 0.00958198f $X=4.42 $Y=5.21 $X2=1.16 $Y2=3.205
cc_127 N_VDD_M1009_b N_CK_M1010_g 0.020128f $X=-0.045 $Y=2.645 $X2=1.46
+ $Y2=3.825
cc_128 N_VDD_c_117_p N_CK_M1010_g 0.00606474f $X=1.95 $Y=5.247 $X2=1.46
+ $Y2=3.825
cc_129 N_VDD_c_118_p N_CK_M1010_g 0.00468827f $X=4.42 $Y=5.21 $X2=1.46 $Y2=3.825
cc_130 N_VDD_M1009_b N_CK_c_294_n 0.00774555f $X=-0.045 $Y=2.645 $X2=2.25
+ $Y2=2.67
cc_131 N_VDD_M1009_b N_CK_M1002_g 0.0214648f $X=-0.045 $Y=2.645 $X2=2.25
+ $Y2=3.825
cc_132 N_VDD_c_132_p N_CK_M1002_g 0.00362996f $X=2.035 $Y=3.205 $X2=2.25
+ $Y2=3.825
cc_133 N_VDD_c_133_p N_CK_M1002_g 0.00606474f $X=2.9 $Y=5.247 $X2=2.25 $Y2=3.825
cc_134 N_VDD_c_120_p N_CK_M1002_g 0.00607189f $X=2.985 $Y=3.545 $X2=2.25
+ $Y2=3.825
cc_135 N_VDD_c_118_p N_CK_M1002_g 0.00468827f $X=4.42 $Y=5.21 $X2=2.25 $Y2=3.825
cc_136 N_VDD_M1009_b N_CK_c_300_n 0.00487051f $X=-0.045 $Y=2.645 $X2=1.4
+ $Y2=2.505
cc_137 N_VDD_M1009_b N_CK_c_310_n 0.00302835f $X=-0.045 $Y=2.645 $X2=2.395
+ $Y2=2.33
cc_138 N_VDD_M1009_b N_CK_c_311_n 0.0022456f $X=-0.045 $Y=2.645 $X2=1.4 $Y2=2.33
cc_139 N_VDD_c_132_p N_CK_c_312_n 0.00634153f $X=2.035 $Y=3.205 $X2=2.25
+ $Y2=2.33
cc_140 N_VDD_M1009_b N_A_157_393#_M1003_g 0.0214821f $X=-0.045 $Y=2.645 $X2=0.86
+ $Y2=3.825
cc_141 N_VDD_c_117_p N_A_157_393#_M1003_g 0.00606474f $X=1.95 $Y=5.247 $X2=0.86
+ $Y2=3.825
cc_142 N_VDD_c_118_p N_A_157_393#_M1003_g 0.00468827f $X=4.42 $Y=5.21 $X2=0.86
+ $Y2=3.825
cc_143 N_VDD_M1009_b N_A_157_393#_c_448_n 0.00156053f $X=-0.045 $Y=2.645
+ $X2=2.465 $Y2=3.205
cc_144 N_VDD_c_133_p N_A_157_393#_c_448_n 0.00736239f $X=2.9 $Y=5.247 $X2=2.465
+ $Y2=3.205
cc_145 N_VDD_c_120_p N_A_157_393#_c_448_n 0.0657863f $X=2.985 $Y=3.545 $X2=2.465
+ $Y2=3.205
cc_146 N_VDD_c_118_p N_A_157_393#_c_448_n 0.00476261f $X=4.42 $Y=5.21 $X2=2.465
+ $Y2=3.205
cc_147 N_VDD_M1009_b N_A_157_393#_c_442_n 0.00551116f $X=-0.045 $Y=2.645
+ $X2=2.735 $Y2=2.84
cc_148 N_VDD_M1009_b N_A_157_393#_c_453_n 0.013496f $X=-0.045 $Y=2.645 $X2=2.735
+ $Y2=2.925
cc_149 N_VDD_M1009_b N_A_349_89#_M1012_g 0.0197647f $X=-0.045 $Y=2.645 $X2=1.82
+ $Y2=3.825
cc_150 N_VDD_c_117_p N_A_349_89#_M1012_g 0.00606474f $X=1.95 $Y=5.247 $X2=1.82
+ $Y2=3.825
cc_151 N_VDD_c_132_p N_A_349_89#_M1012_g 0.00362996f $X=2.035 $Y=3.205 $X2=1.82
+ $Y2=3.825
cc_152 N_VDD_c_118_p N_A_349_89#_M1012_g 0.00468827f $X=4.42 $Y=5.21 $X2=1.82
+ $Y2=3.825
cc_153 N_VDD_M1009_b N_A_349_89#_M1005_g 0.0614895f $X=-0.045 $Y=2.645 $X2=4.15
+ $Y2=4.195
cc_154 N_VDD_c_121_p N_A_349_89#_M1005_g 0.00606474f $X=4.28 $Y=5.247 $X2=4.15
+ $Y2=4.195
cc_155 N_VDD_c_155_p N_A_349_89#_M1005_g 0.00362996f $X=4.365 $Y=4.225 $X2=4.15
+ $Y2=4.195
cc_156 N_VDD_c_118_p N_A_349_89#_M1005_g 0.00468827f $X=4.42 $Y=5.21 $X2=4.15
+ $Y2=4.195
cc_157 N_VDD_M1009_b N_A_349_89#_c_560_n 0.00913636f $X=-0.045 $Y=2.645
+ $X2=4.125 $Y2=2.745
cc_158 N_VDD_M1009_b N_A_349_89#_c_565_n 0.00558439f $X=-0.045 $Y=2.645
+ $X2=3.415 $Y2=3.205
cc_159 N_VDD_c_121_p N_A_349_89#_c_565_n 0.00757793f $X=4.28 $Y=5.247 $X2=3.415
+ $Y2=3.205
cc_160 N_VDD_c_118_p N_A_349_89#_c_565_n 0.00476261f $X=4.42 $Y=5.21 $X2=3.415
+ $Y2=3.205
cc_161 N_VDD_M1009_b N_QN_M1000_g 0.0693077f $X=-0.045 $Y=2.645 $X2=4.58
+ $Y2=4.195
cc_162 N_VDD_c_155_p N_QN_M1000_g 0.00362996f $X=4.365 $Y=4.225 $X2=4.58
+ $Y2=4.195
cc_163 N_VDD_c_163_p N_QN_M1000_g 0.00606474f $X=4.42 $Y=5.21 $X2=4.58 $Y2=4.195
cc_164 N_VDD_c_118_p N_QN_M1000_g 0.00468827f $X=4.42 $Y=5.21 $X2=4.58 $Y2=4.195
cc_165 N_VDD_M1009_b N_QN_c_688_n 0.0229251f $X=-0.045 $Y=2.645 $X2=3.935
+ $Y2=2.7
cc_166 N_VDD_c_121_p N_QN_c_688_n 0.00745733f $X=4.28 $Y=5.247 $X2=3.935 $Y2=2.7
cc_167 N_VDD_c_118_p N_QN_c_688_n 0.00476261f $X=4.42 $Y=5.21 $X2=3.935 $Y2=2.7
cc_168 N_VDD_M1009_b QN 0.00991454f $X=-0.045 $Y=2.645 $X2=3.94 $Y2=2.7
cc_169 N_VDD_M1009_b N_Q_c_762_n 0.0129218f $X=-0.045 $Y=2.645 $X2=4.795
+ $Y2=3.07
cc_170 N_VDD_M1009_b N_Q_c_763_n 0.0240458f $X=-0.045 $Y=2.645 $X2=4.795
+ $Y2=4.225
cc_171 N_VDD_c_163_p N_Q_c_763_n 0.00757793f $X=4.42 $Y=5.21 $X2=4.795 $Y2=4.225
cc_172 N_VDD_c_118_p N_Q_c_763_n 0.00476261f $X=4.42 $Y=5.21 $X2=4.795 $Y2=4.225
cc_173 N_VDD_M1009_b N_Q_c_761_n 0.0126284f $X=-0.045 $Y=2.645 $X2=4.827 $Y2=2.9
cc_174 N_VDD_M1009_b Q 0.0109219f $X=-0.045 $Y=2.645 $X2=4.795 $Y2=3.07
cc_175 N_D_M1014_g N_CK_c_294_n 0.00448096f $X=3.2 $Y=3.825 $X2=2.25 $Y2=2.67
cc_176 N_D_c_198_n N_CK_c_295_n 0.00128484f $X=2.85 $Y=1.59 $X2=2.305 $Y2=2.34
cc_177 N_D_c_175_n N_CK_c_296_n 0.040252f $X=0.44 $Y=1.88 $X2=0.92 $Y2=1.59
cc_178 N_D_c_219_p N_CK_c_296_n 0.0023548f $X=0.99 $Y=1.17 $X2=0.92 $Y2=1.59
cc_179 N_D_c_198_n N_CK_c_296_n 0.00407483f $X=2.85 $Y=1.59 $X2=0.92 $Y2=1.59
cc_180 N_D_c_200_n N_CK_c_296_n 9.79344e-19 $X=0.725 $Y=1.59 $X2=0.92 $Y2=1.59
cc_181 N_D_M1001_g N_CK_c_297_n 0.040252f $X=0.5 $Y=0.945 $X2=0.92 $Y2=1.425
cc_182 N_D_c_190_n N_CK_c_297_n 0.0052197f $X=0.58 $Y=1.59 $X2=0.92 $Y2=1.425
cc_183 N_D_c_219_p N_CK_c_297_n 0.0149528f $X=0.99 $Y=1.17 $X2=0.92 $Y2=1.425
cc_184 N_D_c_225_p N_CK_c_300_n 0.00150627f $X=0.99 $Y=2.925 $X2=1.4 $Y2=2.505
cc_185 N_D_c_188_n N_CK_c_306_n 0.00662135f $X=3.2 $Y=1.59 $X2=2.277 $Y2=1.575
cc_186 N_D_c_195_n N_CK_c_306_n 3.50905e-19 $X=2.995 $Y=1.59 $X2=2.277 $Y2=1.575
cc_187 N_D_c_198_n N_CK_c_306_n 0.0082638f $X=2.85 $Y=1.59 $X2=2.277 $Y2=1.575
cc_188 N_D_c_175_n N_CK_c_307_n 7.00514e-19 $X=0.44 $Y=1.88 $X2=0.92 $Y2=1.59
cc_189 N_D_c_176_n N_CK_c_307_n 2.73444e-19 $X=0.44 $Y=1.96 $X2=0.92 $Y2=1.59
cc_190 N_D_M1001_g N_CK_c_307_n 4.01349e-19 $X=0.5 $Y=0.945 $X2=0.92 $Y2=1.59
cc_191 N_D_c_190_n N_CK_c_307_n 0.0567541f $X=0.58 $Y=1.59 $X2=0.92 $Y2=1.59
cc_192 N_D_c_219_p N_CK_c_307_n 0.0103829f $X=0.99 $Y=1.17 $X2=0.92 $Y2=1.59
cc_193 N_D_c_198_n N_CK_c_307_n 0.0133835f $X=2.85 $Y=1.59 $X2=0.92 $Y2=1.59
cc_194 N_D_c_200_n N_CK_c_307_n 0.00180575f $X=0.725 $Y=1.59 $X2=0.92 $Y2=1.59
cc_195 D N_CK_c_307_n 0.00563597f $X=0.44 $Y=1.96 $X2=0.92 $Y2=1.59
cc_196 N_D_c_225_p N_CK_c_308_n 0.012157f $X=0.99 $Y=2.925 $X2=1.315 $Y2=2.33
cc_197 N_D_c_198_n N_CK_c_308_n 0.00774794f $X=2.85 $Y=1.59 $X2=1.315 $Y2=2.33
cc_198 N_D_c_191_n N_CK_c_309_n 0.0128995f $X=0.58 $Y=2.84 $X2=1.005 $Y2=2.33
cc_199 N_D_c_225_p N_CK_c_309_n 0.0056307f $X=0.99 $Y=2.925 $X2=1.005 $Y2=2.33
cc_200 N_D_c_191_n N_CK_c_311_n 0.00613815f $X=0.58 $Y=2.84 $X2=1.4 $Y2=2.33
cc_201 N_D_c_225_p N_CK_c_311_n 0.00103871f $X=0.99 $Y=2.925 $X2=1.4 $Y2=2.33
cc_202 N_D_c_198_n N_CK_c_311_n 6.39375e-19 $X=2.85 $Y=1.59 $X2=1.4 $Y2=2.33
cc_203 N_D_c_191_n N_CK_c_313_n 0.00128303f $X=0.58 $Y=2.84 $X2=1.545 $Y2=2.33
cc_204 N_D_c_225_p N_CK_c_313_n 0.00146098f $X=0.99 $Y=2.925 $X2=1.545 $Y2=2.33
cc_205 N_D_c_198_n N_CK_c_313_n 0.0144351f $X=2.85 $Y=1.59 $X2=1.545 $Y2=2.33
cc_206 N_D_c_187_n N_A_157_393#_M1003_g 0.0889164f $X=0.44 $Y=2.155 $X2=0.86
+ $Y2=3.825
cc_207 N_D_c_191_n N_A_157_393#_M1003_g 0.00439102f $X=0.58 $Y=2.84 $X2=0.86
+ $Y2=3.825
cc_208 N_D_c_225_p N_A_157_393#_M1003_g 0.0174985f $X=0.99 $Y=2.925 $X2=0.86
+ $Y2=3.825
cc_209 N_D_c_198_n N_A_157_393#_c_428_n 0.00419102f $X=2.85 $Y=1.59 $X2=1.265
+ $Y2=2.04
cc_210 N_D_c_176_n N_A_157_393#_c_429_n 0.0889164f $X=0.44 $Y=1.96 $X2=0.935
+ $Y2=2.04
cc_211 N_D_c_197_n N_A_157_393#_c_429_n 0.00439102f $X=0.44 $Y=1.96 $X2=0.935
+ $Y2=2.04
cc_212 N_D_c_198_n N_A_157_393#_c_429_n 5.19983e-19 $X=2.85 $Y=1.59 $X2=0.935
+ $Y2=2.04
cc_213 D N_A_157_393#_c_429_n 0.00144527f $X=0.44 $Y=1.96 $X2=0.935 $Y2=2.04
cc_214 N_D_c_175_n N_A_157_393#_c_430_n 0.00201381f $X=0.44 $Y=1.88 $X2=1.34
+ $Y2=1.965
cc_215 N_D_c_219_p N_A_157_393#_c_431_n 0.00182707f $X=0.99 $Y=1.17 $X2=1.4
+ $Y2=1.59
cc_216 N_D_c_198_n N_A_157_393#_c_431_n 0.0113766f $X=2.85 $Y=1.59 $X2=1.4
+ $Y2=1.59
cc_217 N_D_c_219_p N_A_157_393#_c_435_n 0.00435378f $X=0.99 $Y=1.17 $X2=2.38
+ $Y2=1.59
cc_218 N_D_c_198_n N_A_157_393#_c_435_n 0.0492477f $X=2.85 $Y=1.59 $X2=2.38
+ $Y2=1.59
cc_219 N_D_c_182_n N_A_157_393#_c_437_n 0.00724066f $X=3.2 $Y=1.425 $X2=2.465
+ $Y2=0.825
cc_220 N_D_c_188_n N_A_157_393#_c_437_n 0.00153999f $X=3.2 $Y=1.59 $X2=2.465
+ $Y2=0.825
cc_221 N_D_c_202_n N_A_157_393#_c_437_n 0.00126742f $X=2.995 $Y=1.59 $X2=2.465
+ $Y2=0.825
cc_222 N_D_M1014_g N_A_157_393#_c_441_n 0.00201047f $X=3.2 $Y=3.825 $X2=2.465
+ $Y2=1.845
cc_223 N_D_c_188_n N_A_157_393#_c_441_n 0.00153999f $X=3.2 $Y=1.59 $X2=2.465
+ $Y2=1.845
cc_224 N_D_c_202_n N_A_157_393#_c_441_n 0.00126742f $X=2.995 $Y=1.59 $X2=2.465
+ $Y2=1.845
cc_225 N_D_M1014_g N_A_157_393#_c_448_n 0.00932885f $X=3.2 $Y=3.825 $X2=2.465
+ $Y2=3.205
cc_226 N_D_M1014_g N_A_157_393#_c_442_n 0.012583f $X=3.2 $Y=3.825 $X2=2.735
+ $Y2=2.84
cc_227 N_D_c_188_n N_A_157_393#_c_443_n 5.35151e-19 $X=3.2 $Y=1.59 $X2=2.465
+ $Y2=1.59
cc_228 N_D_c_195_n N_A_157_393#_c_443_n 0.00755683f $X=2.995 $Y=1.59 $X2=2.465
+ $Y2=1.59
cc_229 N_D_c_198_n N_A_157_393#_c_443_n 0.0171747f $X=2.85 $Y=1.59 $X2=2.465
+ $Y2=1.59
cc_230 N_D_M1014_g N_A_157_393#_c_444_n 0.0023936f $X=3.2 $Y=3.825 $X2=2.735
+ $Y2=1.93
cc_231 N_D_c_198_n N_A_157_393#_c_444_n 0.00219678f $X=2.85 $Y=1.59 $X2=2.735
+ $Y2=1.93
cc_232 N_D_M1014_g N_A_157_393#_c_453_n 0.00340068f $X=3.2 $Y=3.825 $X2=2.735
+ $Y2=2.925
cc_233 N_D_c_198_n N_A_349_89#_M1004_g 0.00707887f $X=2.85 $Y=1.59 $X2=1.82
+ $Y2=0.945
cc_234 N_D_c_198_n N_A_349_89#_c_555_n 0.00187603f $X=2.85 $Y=1.59 $X2=1.88
+ $Y2=1.93
cc_235 N_D_M1014_g N_A_349_89#_c_556_n 0.0046172f $X=3.2 $Y=3.825 $X2=4.035
+ $Y2=1.93
cc_236 N_D_c_198_n N_A_349_89#_c_561_n 0.00166223f $X=2.85 $Y=1.59 $X2=1.88
+ $Y2=1.93
cc_237 N_D_c_182_n N_A_349_89#_c_562_n 0.0251298f $X=3.2 $Y=1.425 $X2=3.415
+ $Y2=0.825
cc_238 N_D_c_195_n N_A_349_89#_c_562_n 0.0115453f $X=2.995 $Y=1.59 $X2=3.415
+ $Y2=0.825
cc_239 N_D_c_202_n N_A_349_89#_c_562_n 0.00389142f $X=2.995 $Y=1.59 $X2=3.415
+ $Y2=0.825
cc_240 N_D_M1014_g N_A_349_89#_c_565_n 0.025216f $X=3.2 $Y=3.825 $X2=3.415
+ $Y2=3.205
cc_241 N_D_M1014_g N_A_349_89#_c_567_n 0.00245806f $X=3.2 $Y=3.825 $X2=3.415
+ $Y2=1.93
cc_242 N_D_M1014_g N_A_349_89#_c_568_n 0.0167433f $X=3.2 $Y=3.825 $X2=3.89
+ $Y2=1.93
cc_243 N_D_c_188_n N_A_349_89#_c_568_n 0.0041429f $X=3.2 $Y=1.59 $X2=3.89
+ $Y2=1.93
cc_244 N_D_c_195_n N_A_349_89#_c_568_n 0.00508416f $X=2.995 $Y=1.59 $X2=3.89
+ $Y2=1.93
cc_245 N_D_c_198_n N_A_349_89#_c_568_n 0.0735565f $X=2.85 $Y=1.59 $X2=3.89
+ $Y2=1.93
cc_246 N_D_c_202_n N_A_349_89#_c_568_n 0.0291144f $X=2.995 $Y=1.59 $X2=3.89
+ $Y2=1.93
cc_247 N_D_c_198_n N_A_349_89#_c_569_n 0.0289631f $X=2.85 $Y=1.59 $X2=2.025
+ $Y2=1.93
cc_248 N_D_c_225_p A_115_565# 0.00473129f $X=0.99 $Y=2.925 $X2=0.575 $Y2=2.825
cc_249 N_D_c_290_p A_115_565# 0.00144354f $X=0.665 $Y=2.925 $X2=0.575 $Y2=2.825
cc_250 N_D_c_190_n A_115_115# 6.64472e-19 $X=0.58 $Y=1.59 $X2=0.575 $Y2=0.575
cc_251 N_D_c_219_p A_115_115# 0.00317038f $X=0.99 $Y=1.17 $X2=0.575 $Y2=0.575
cc_252 N_D_c_293_p A_115_115# 0.00148865f $X=0.665 $Y=1.17 $X2=0.575 $Y2=0.575
cc_253 N_CK_M1010_g N_A_157_393#_M1003_g 0.0441985f $X=1.46 $Y=3.825 $X2=0.86
+ $Y2=3.825
cc_254 N_CK_c_300_n N_A_157_393#_M1003_g 0.0118393f $X=1.4 $Y=2.505 $X2=0.86
+ $Y2=3.825
cc_255 N_CK_c_307_n N_A_157_393#_M1003_g 0.00391544f $X=0.92 $Y=1.59 $X2=0.86
+ $Y2=3.825
cc_256 N_CK_c_309_n N_A_157_393#_M1003_g 0.0079407f $X=1.005 $Y=2.33 $X2=0.86
+ $Y2=3.825
cc_257 N_CK_c_311_n N_A_157_393#_M1003_g 0.00128351f $X=1.4 $Y=2.33 $X2=0.86
+ $Y2=3.825
cc_258 N_CK_c_313_n N_A_157_393#_M1003_g 4.61617e-19 $X=1.545 $Y=2.33 $X2=0.86
+ $Y2=3.825
cc_259 N_CK_c_300_n N_A_157_393#_c_428_n 0.00904036f $X=1.4 $Y=2.505 $X2=1.265
+ $Y2=2.04
cc_260 N_CK_c_307_n N_A_157_393#_c_428_n 0.00909647f $X=0.92 $Y=1.59 $X2=1.265
+ $Y2=2.04
cc_261 N_CK_c_308_n N_A_157_393#_c_428_n 0.00939103f $X=1.315 $Y=2.33 $X2=1.265
+ $Y2=2.04
cc_262 N_CK_c_311_n N_A_157_393#_c_428_n 0.00102633f $X=1.4 $Y=2.33 $X2=1.265
+ $Y2=2.04
cc_263 N_CK_c_313_n N_A_157_393#_c_428_n 0.00131242f $X=1.545 $Y=2.33 $X2=1.265
+ $Y2=2.04
cc_264 N_CK_c_296_n N_A_157_393#_c_429_n 0.018421f $X=0.92 $Y=1.59 $X2=0.935
+ $Y2=2.04
cc_265 N_CK_c_307_n N_A_157_393#_c_429_n 0.00314767f $X=0.92 $Y=1.59 $X2=0.935
+ $Y2=2.04
cc_266 N_CK_c_307_n N_A_157_393#_c_430_n 0.0045597f $X=0.92 $Y=1.59 $X2=1.34
+ $Y2=1.965
cc_267 N_CK_c_296_n N_A_157_393#_c_431_n 0.0220721f $X=0.92 $Y=1.59 $X2=1.4
+ $Y2=1.59
cc_268 N_CK_c_300_n N_A_157_393#_c_431_n 0.00227671f $X=1.4 $Y=2.505 $X2=1.4
+ $Y2=1.59
cc_269 N_CK_c_307_n N_A_157_393#_c_431_n 0.00131283f $X=0.92 $Y=1.59 $X2=1.4
+ $Y2=1.59
cc_270 N_CK_c_311_n N_A_157_393#_c_431_n 5.27321e-19 $X=1.4 $Y=2.33 $X2=1.4
+ $Y2=1.59
cc_271 N_CK_c_313_n N_A_157_393#_c_431_n 8.78837e-19 $X=1.545 $Y=2.33 $X2=1.4
+ $Y2=1.59
cc_272 N_CK_c_297_n N_A_157_393#_c_432_n 0.0219663f $X=0.92 $Y=1.425 $X2=1.4
+ $Y2=1.425
cc_273 N_CK_c_295_n N_A_157_393#_c_435_n 0.00592387f $X=2.305 $Y=2.34 $X2=2.38
+ $Y2=1.59
cc_274 N_CK_c_296_n N_A_157_393#_c_435_n 8.05876e-19 $X=0.92 $Y=1.59 $X2=2.38
+ $Y2=1.59
cc_275 N_CK_c_300_n N_A_157_393#_c_435_n 5.56676e-19 $X=1.4 $Y=2.505 $X2=2.38
+ $Y2=1.59
cc_276 N_CK_c_306_n N_A_157_393#_c_435_n 0.00762848f $X=2.277 $Y=1.575 $X2=2.38
+ $Y2=1.59
cc_277 N_CK_c_307_n N_A_157_393#_c_435_n 0.00853323f $X=0.92 $Y=1.59 $X2=2.38
+ $Y2=1.59
cc_278 N_CK_c_308_n N_A_157_393#_c_435_n 0.00132148f $X=1.315 $Y=2.33 $X2=2.38
+ $Y2=1.59
cc_279 N_CK_c_310_n N_A_157_393#_c_435_n 8.24249e-19 $X=2.395 $Y=2.33 $X2=2.38
+ $Y2=1.59
cc_280 N_CK_c_311_n N_A_157_393#_c_435_n 0.00261697f $X=1.4 $Y=2.33 $X2=2.38
+ $Y2=1.59
cc_281 N_CK_c_312_n N_A_157_393#_c_435_n 0.00341454f $X=2.25 $Y=2.33 $X2=2.38
+ $Y2=1.59
cc_282 N_CK_c_313_n N_A_157_393#_c_435_n 0.00221563f $X=1.545 $Y=2.33 $X2=2.38
+ $Y2=1.59
cc_283 N_CK_c_301_n N_A_157_393#_c_437_n 0.0109347f $X=2.277 $Y=1.425 $X2=2.465
+ $Y2=0.825
cc_284 N_CK_c_306_n N_A_157_393#_c_437_n 0.0022869f $X=2.277 $Y=1.575 $X2=2.465
+ $Y2=0.825
cc_285 N_CK_c_295_n N_A_157_393#_c_441_n 0.00595506f $X=2.305 $Y=2.34 $X2=2.465
+ $Y2=1.845
cc_286 N_CK_c_294_n N_A_157_393#_c_442_n 0.0033284f $X=2.25 $Y=2.67 $X2=2.735
+ $Y2=2.84
cc_287 N_CK_M1002_g N_A_157_393#_c_442_n 0.00491946f $X=2.25 $Y=3.825 $X2=2.735
+ $Y2=2.84
cc_288 N_CK_c_295_n N_A_157_393#_c_442_n 0.00747875f $X=2.305 $Y=2.34 $X2=2.735
+ $Y2=2.84
cc_289 N_CK_c_310_n N_A_157_393#_c_442_n 0.0288018f $X=2.395 $Y=2.33 $X2=2.735
+ $Y2=2.84
cc_290 CK N_A_157_393#_c_442_n 0.00851352f $X=2.395 $Y=2.33 $X2=2.735 $Y2=2.84
cc_291 N_CK_c_295_n N_A_157_393#_c_443_n 0.00114916f $X=2.305 $Y=2.34 $X2=2.465
+ $Y2=1.59
cc_292 N_CK_c_306_n N_A_157_393#_c_443_n 8.09104e-19 $X=2.277 $Y=1.575 $X2=2.465
+ $Y2=1.59
cc_293 N_CK_c_294_n N_A_157_393#_c_444_n 0.00157237f $X=2.25 $Y=2.67 $X2=2.735
+ $Y2=1.93
cc_294 N_CK_c_295_n N_A_157_393#_c_444_n 0.00436926f $X=2.305 $Y=2.34 $X2=2.735
+ $Y2=1.93
cc_295 N_CK_c_310_n N_A_157_393#_c_444_n 0.00529105f $X=2.395 $Y=2.33 $X2=2.735
+ $Y2=1.93
cc_296 CK N_A_157_393#_c_444_n 8.76467e-19 $X=2.395 $Y=2.33 $X2=2.735 $Y2=1.93
cc_297 N_CK_c_294_n N_A_157_393#_c_453_n 0.00260941f $X=2.25 $Y=2.67 $X2=2.735
+ $Y2=2.925
cc_298 N_CK_c_310_n N_A_157_393#_c_453_n 0.00706443f $X=2.395 $Y=2.33 $X2=2.735
+ $Y2=2.925
cc_299 CK N_A_157_393#_c_453_n 0.00259785f $X=2.395 $Y=2.33 $X2=2.735 $Y2=2.925
cc_300 N_CK_c_295_n N_A_349_89#_M1004_g 0.00697006f $X=2.305 $Y=2.34 $X2=1.82
+ $Y2=0.945
cc_301 N_CK_c_301_n N_A_349_89#_M1004_g 0.0306464f $X=2.277 $Y=1.425 $X2=1.82
+ $Y2=0.945
cc_302 N_CK_c_294_n N_A_349_89#_M1012_g 0.0294691f $X=2.25 $Y=2.67 $X2=1.82
+ $Y2=3.825
cc_303 N_CK_c_295_n N_A_349_89#_M1012_g 0.0175925f $X=2.305 $Y=2.34 $X2=1.82
+ $Y2=3.825
cc_304 N_CK_c_300_n N_A_349_89#_M1012_g 0.156645f $X=1.4 $Y=2.505 $X2=1.82
+ $Y2=3.825
cc_305 N_CK_c_310_n N_A_349_89#_M1012_g 0.0026346f $X=2.395 $Y=2.33 $X2=1.82
+ $Y2=3.825
cc_306 N_CK_c_311_n N_A_349_89#_M1012_g 0.00453616f $X=1.4 $Y=2.33 $X2=1.82
+ $Y2=3.825
cc_307 N_CK_c_312_n N_A_349_89#_M1012_g 0.0112778f $X=2.25 $Y=2.33 $X2=1.82
+ $Y2=3.825
cc_308 N_CK_c_313_n N_A_349_89#_M1012_g 0.00113587f $X=1.545 $Y=2.33 $X2=1.82
+ $Y2=3.825
cc_309 CK N_A_349_89#_M1012_g 3.05655e-19 $X=2.395 $Y=2.33 $X2=1.82 $Y2=3.825
cc_310 N_CK_c_295_n N_A_349_89#_c_555_n 0.0213817f $X=2.305 $Y=2.34 $X2=1.88
+ $Y2=1.93
cc_311 N_CK_c_312_n N_A_349_89#_c_555_n 0.00185875f $X=2.25 $Y=2.33 $X2=1.88
+ $Y2=1.93
cc_312 N_CK_c_295_n N_A_349_89#_c_561_n 8.95026e-19 $X=2.305 $Y=2.34 $X2=1.88
+ $Y2=1.93
cc_313 N_CK_c_312_n N_A_349_89#_c_561_n 0.00488871f $X=2.25 $Y=2.33 $X2=1.88
+ $Y2=1.93
cc_314 N_CK_c_294_n N_A_349_89#_c_568_n 2.34467e-19 $X=2.25 $Y=2.67 $X2=3.89
+ $Y2=1.93
cc_315 N_CK_c_295_n N_A_349_89#_c_568_n 0.0033485f $X=2.305 $Y=2.34 $X2=3.89
+ $Y2=1.93
cc_316 N_CK_c_310_n N_A_349_89#_c_568_n 8.38639e-19 $X=2.395 $Y=2.33 $X2=3.89
+ $Y2=1.93
cc_317 N_CK_c_312_n N_A_349_89#_c_568_n 0.0179446f $X=2.25 $Y=2.33 $X2=3.89
+ $Y2=1.93
cc_318 CK N_A_349_89#_c_568_n 0.0248956f $X=2.395 $Y=2.33 $X2=3.89 $Y2=1.93
cc_319 N_CK_c_295_n N_A_349_89#_c_569_n 8.66236e-19 $X=2.305 $Y=2.34 $X2=2.025
+ $Y2=1.93
cc_320 N_CK_c_312_n N_A_349_89#_c_569_n 0.0247156f $X=2.25 $Y=2.33 $X2=2.025
+ $Y2=1.93
cc_321 N_A_157_393#_c_430_n N_A_349_89#_M1004_g 0.00733314f $X=1.34 $Y=1.965
+ $X2=1.82 $Y2=0.945
cc_322 N_A_157_393#_c_432_n N_A_349_89#_M1004_g 0.081251f $X=1.4 $Y=1.425
+ $X2=1.82 $Y2=0.945
cc_323 N_A_157_393#_c_435_n N_A_349_89#_M1004_g 0.0107575f $X=2.38 $Y=1.59
+ $X2=1.82 $Y2=0.945
cc_324 N_A_157_393#_c_428_n N_A_349_89#_c_555_n 0.00733314f $X=1.265 $Y=2.04
+ $X2=1.88 $Y2=1.93
cc_325 N_A_157_393#_c_435_n N_A_349_89#_c_555_n 0.00290516f $X=2.38 $Y=1.59
+ $X2=1.88 $Y2=1.93
cc_326 N_A_157_393#_c_444_n N_A_349_89#_c_555_n 2.96928e-19 $X=2.735 $Y=1.93
+ $X2=1.88 $Y2=1.93
cc_327 N_A_157_393#_c_430_n N_A_349_89#_c_561_n 0.00352413f $X=1.34 $Y=1.965
+ $X2=1.88 $Y2=1.93
cc_328 N_A_157_393#_c_435_n N_A_349_89#_c_561_n 0.0219931f $X=2.38 $Y=1.59
+ $X2=1.88 $Y2=1.93
cc_329 N_A_157_393#_c_444_n N_A_349_89#_c_561_n 0.00559532f $X=2.735 $Y=1.93
+ $X2=1.88 $Y2=1.93
cc_330 N_A_157_393#_c_442_n N_A_349_89#_c_565_n 0.0285298f $X=2.735 $Y=2.84
+ $X2=3.415 $Y2=3.205
cc_331 N_A_157_393#_c_444_n N_A_349_89#_c_567_n 0.0038132f $X=2.735 $Y=1.93
+ $X2=3.415 $Y2=1.93
cc_332 N_A_157_393#_c_435_n N_A_349_89#_c_568_n 0.00314603f $X=2.38 $Y=1.59
+ $X2=3.89 $Y2=1.93
cc_333 N_A_157_393#_c_441_n N_A_349_89#_c_568_n 6.94255e-19 $X=2.465 $Y=1.845
+ $X2=3.89 $Y2=1.93
cc_334 N_A_157_393#_c_442_n N_A_349_89#_c_568_n 0.00464833f $X=2.735 $Y=2.84
+ $X2=3.89 $Y2=1.93
cc_335 N_A_157_393#_c_444_n N_A_349_89#_c_568_n 0.0225447f $X=2.735 $Y=1.93
+ $X2=3.89 $Y2=1.93
cc_336 N_A_157_393#_c_430_n N_A_349_89#_c_569_n 9.10135e-19 $X=1.34 $Y=1.965
+ $X2=2.025 $Y2=1.93
cc_337 N_A_157_393#_c_435_n N_A_349_89#_c_569_n 0.0010261f $X=2.38 $Y=1.59
+ $X2=2.025 $Y2=1.93
cc_338 N_A_157_393#_c_441_n N_A_349_89#_c_569_n 0.00122156f $X=2.465 $Y=1.845
+ $X2=2.025 $Y2=1.93
cc_339 N_A_349_89#_M1008_g N_QN_M1011_g 0.030339f $X=4.15 $Y=0.835 $X2=4.58
+ $Y2=0.835
cc_340 N_A_349_89#_c_557_n N_QN_M1011_g 0.0153126f $X=4.037 $Y=1.765 $X2=4.58
+ $Y2=0.835
cc_341 N_A_349_89#_c_566_n N_QN_M1011_g 4.79563e-19 $X=4.035 $Y=1.93 $X2=4.58
+ $Y2=0.835
cc_342 N_A_349_89#_c_559_n N_QN_M1000_g 0.0102931f $X=4.125 $Y=2.595 $X2=4.58
+ $Y2=4.195
cc_343 N_A_349_89#_c_560_n N_QN_M1000_g 0.0668032f $X=4.125 $Y=2.745 $X2=4.58
+ $Y2=4.195
cc_344 N_A_349_89#_c_556_n N_QN_c_684_n 0.021196f $X=4.035 $Y=1.93 $X2=4.52
+ $Y2=2.135
cc_345 N_A_349_89#_c_566_n N_QN_c_684_n 3.0115e-19 $X=4.035 $Y=1.93 $X2=4.52
+ $Y2=2.135
cc_346 N_A_349_89#_c_570_n N_QN_c_684_n 4.60229e-19 $X=4.035 $Y=1.93 $X2=4.52
+ $Y2=2.135
cc_347 N_A_349_89#_M1008_g N_QN_c_685_n 0.0144755f $X=4.15 $Y=0.835 $X2=3.935
+ $Y2=0.74
cc_348 N_A_349_89#_c_558_n N_QN_c_685_n 0.00485394f $X=4.125 $Y=1.54 $X2=3.935
+ $Y2=0.74
cc_349 N_A_349_89#_c_562_n N_QN_c_685_n 0.0405988f $X=3.415 $Y=0.825 $X2=3.935
+ $Y2=0.74
cc_350 N_A_349_89#_M1005_g N_QN_c_688_n 0.041548f $X=4.15 $Y=4.195 $X2=3.935
+ $Y2=2.7
cc_351 N_A_349_89#_c_559_n N_QN_c_688_n 0.00567875f $X=4.125 $Y=2.595 $X2=3.935
+ $Y2=2.7
cc_352 N_A_349_89#_c_565_n N_QN_c_688_n 0.0937909f $X=3.415 $Y=3.205 $X2=3.935
+ $Y2=2.7
cc_353 N_A_349_89#_c_557_n N_QN_c_689_n 0.00799433f $X=4.037 $Y=1.765 $X2=4.435
+ $Y2=1.59
cc_354 N_A_349_89#_c_558_n N_QN_c_689_n 0.011031f $X=4.125 $Y=1.54 $X2=4.435
+ $Y2=1.59
cc_355 N_A_349_89#_c_566_n N_QN_c_689_n 0.0110498f $X=4.035 $Y=1.93 $X2=4.435
+ $Y2=1.59
cc_356 N_A_349_89#_c_570_n N_QN_c_689_n 0.00387586f $X=4.035 $Y=1.93 $X2=4.435
+ $Y2=1.59
cc_357 N_A_349_89#_c_556_n N_QN_c_691_n 0.00308111f $X=4.035 $Y=1.93 $X2=4.02
+ $Y2=1.59
cc_358 N_A_349_89#_c_562_n N_QN_c_691_n 0.00869401f $X=3.415 $Y=0.825 $X2=4.02
+ $Y2=1.59
cc_359 N_A_349_89#_c_566_n N_QN_c_691_n 0.0120703f $X=4.035 $Y=1.93 $X2=4.02
+ $Y2=1.59
cc_360 N_A_349_89#_c_568_n N_QN_c_691_n 0.0010572f $X=3.89 $Y=1.93 $X2=4.02
+ $Y2=1.59
cc_361 N_A_349_89#_c_570_n N_QN_c_691_n 0.00336135f $X=4.035 $Y=1.93 $X2=4.02
+ $Y2=1.59
cc_362 N_A_349_89#_c_559_n N_QN_c_692_n 0.016126f $X=4.125 $Y=2.595 $X2=4.435
+ $Y2=2.505
cc_363 N_A_349_89#_c_560_n N_QN_c_692_n 0.00248624f $X=4.125 $Y=2.745 $X2=4.435
+ $Y2=2.505
cc_364 N_A_349_89#_c_566_n N_QN_c_692_n 0.00426371f $X=4.035 $Y=1.93 $X2=4.435
+ $Y2=2.505
cc_365 N_A_349_89#_c_570_n N_QN_c_692_n 0.00253233f $X=4.035 $Y=1.93 $X2=4.435
+ $Y2=2.505
cc_366 N_A_349_89#_c_556_n N_QN_c_693_n 0.00265611f $X=4.035 $Y=1.93 $X2=4.02
+ $Y2=2.505
cc_367 N_A_349_89#_c_565_n N_QN_c_693_n 0.00859877f $X=3.415 $Y=3.205 $X2=4.02
+ $Y2=2.505
cc_368 N_A_349_89#_c_566_n N_QN_c_693_n 0.00471962f $X=4.035 $Y=1.93 $X2=4.02
+ $Y2=2.505
cc_369 N_A_349_89#_c_568_n N_QN_c_693_n 9.40773e-19 $X=3.89 $Y=1.93 $X2=4.02
+ $Y2=2.505
cc_370 N_A_349_89#_c_570_n N_QN_c_693_n 0.00140341f $X=4.035 $Y=1.93 $X2=4.02
+ $Y2=2.505
cc_371 N_A_349_89#_c_556_n N_QN_c_694_n 0.00216137f $X=4.035 $Y=1.93 $X2=4.52
+ $Y2=2.135
cc_372 N_A_349_89#_c_557_n N_QN_c_694_n 0.00323473f $X=4.037 $Y=1.765 $X2=4.52
+ $Y2=2.135
cc_373 N_A_349_89#_c_559_n N_QN_c_694_n 0.00226435f $X=4.125 $Y=2.595 $X2=4.52
+ $Y2=2.135
cc_374 N_A_349_89#_c_566_n N_QN_c_694_n 0.00987106f $X=4.035 $Y=1.93 $X2=4.52
+ $Y2=2.135
cc_375 N_A_349_89#_c_570_n N_QN_c_694_n 0.00377439f $X=4.035 $Y=1.93 $X2=4.52
+ $Y2=2.135
cc_376 N_A_349_89#_M1005_g QN 0.00233644f $X=4.15 $Y=4.195 $X2=3.94 $Y2=2.7
cc_377 N_A_349_89#_c_560_n QN 0.00507218f $X=4.125 $Y=2.745 $X2=3.94 $Y2=2.7
cc_378 N_A_349_89#_c_565_n QN 0.00717604f $X=3.415 $Y=3.205 $X2=3.94 $Y2=2.7
cc_379 N_A_349_89#_c_566_n QN 0.00350993f $X=4.035 $Y=1.93 $X2=3.94 $Y2=2.7
cc_380 N_A_349_89#_c_570_n QN 0.00842298f $X=4.035 $Y=1.93 $X2=3.94 $Y2=2.7
cc_381 N_A_349_89#_M1005_g Q 0.00113884f $X=4.15 $Y=4.195 $X2=4.795 $Y2=3.07
cc_382 N_QN_M1000_g N_Q_c_762_n 0.0347947f $X=4.58 $Y=4.195 $X2=4.795 $Y2=3.07
cc_383 N_QN_M1011_g N_Q_c_761_n 0.0493233f $X=4.58 $Y=0.835 $X2=4.827 $Y2=2.9
cc_384 N_QN_c_689_n N_Q_c_761_n 0.0135849f $X=4.435 $Y=1.59 $X2=4.827 $Y2=2.9
cc_385 N_QN_c_692_n N_Q_c_761_n 0.0135849f $X=4.435 $Y=2.505 $X2=4.827 $Y2=2.9
cc_386 N_QN_c_694_n N_Q_c_761_n 0.052716f $X=4.52 $Y=2.135 $X2=4.827 $Y2=2.9
cc_387 N_QN_M1000_g Q 0.0145734f $X=4.58 $Y=4.195 $X2=4.795 $Y2=3.07
cc_388 N_QN_c_688_n Q 0.00553755f $X=3.935 $Y=2.7 $X2=4.795 $Y2=3.07
cc_389 N_QN_c_692_n Q 0.00245821f $X=4.435 $Y=2.505 $X2=4.795 $Y2=3.07
