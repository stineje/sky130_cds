magic
tech sky130A
magscale 1 2
timestamp 1606864607
<< checkpaint >>
rect -1209 -1243 1481 2575
<< nwell >>
rect -9 581 286 1341
<< nmos >>
rect 80 115 110 315
rect 152 115 182 315
<< pmos >>
rect 80 617 110 1217
rect 166 617 196 1217
<< ndiff >>
rect 27 267 80 315
rect 27 131 35 267
rect 69 131 80 267
rect 27 115 80 131
rect 110 115 152 315
rect 182 267 235 315
rect 182 131 193 267
rect 227 131 235 267
rect 182 115 235 131
<< pdiff >>
rect 27 1201 80 1217
rect 27 793 35 1201
rect 69 793 80 1201
rect 27 617 80 793
rect 110 1201 166 1217
rect 110 657 121 1201
rect 155 657 166 1201
rect 110 617 166 657
rect 196 1201 249 1217
rect 196 725 207 1201
rect 241 725 249 1201
rect 196 617 249 725
<< ndiffc >>
rect 35 131 69 267
rect 193 131 227 267
<< pdiffc >>
rect 35 793 69 1201
rect 121 657 155 1201
rect 207 725 241 1201
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1271 51 1305
rect 85 1271 109 1305
rect 163 1271 187 1305
rect 221 1271 245 1305
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1271 85 1305
rect 187 1271 221 1305
<< poly >>
rect 80 1217 110 1243
rect 166 1217 196 1243
rect 80 570 110 617
rect 37 554 110 570
rect 37 520 47 554
rect 81 520 110 554
rect 37 504 110 520
rect 80 315 110 504
rect 166 477 196 617
rect 152 461 210 477
rect 152 427 166 461
rect 200 427 210 461
rect 152 411 210 427
rect 152 315 182 411
rect 80 89 110 115
rect 152 89 182 115
<< polycont >>
rect 47 520 81 554
rect 166 427 200 461
<< locali >>
rect 0 1311 286 1332
rect 0 1271 51 1311
rect 85 1271 187 1311
rect 221 1271 286 1311
rect 35 1201 69 1271
rect 35 777 69 793
rect 121 1201 155 1217
rect 47 554 81 649
rect 47 504 81 520
rect 207 1201 241 1271
rect 207 709 241 725
rect 121 535 155 657
rect 195 461 229 575
rect 150 427 166 461
rect 200 427 229 461
rect 35 267 69 279
rect 35 115 69 131
rect 193 267 227 283
rect 193 61 227 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 286 61
rect 0 0 286 21
<< viali >>
rect 51 1305 85 1311
rect 51 1277 85 1305
rect 187 1305 221 1311
rect 187 1277 221 1305
rect 47 649 81 683
rect 121 501 155 535
rect 195 575 229 609
rect 35 279 69 313
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1311 286 1332
rect 0 1277 51 1311
rect 85 1277 187 1311
rect 221 1277 286 1311
rect 0 1271 286 1277
rect 35 683 93 689
rect 35 649 47 683
rect 81 649 115 683
rect 35 643 93 649
rect 183 609 241 615
rect 161 575 195 609
rect 229 575 241 609
rect 183 569 241 575
rect 109 535 167 541
rect 109 501 121 535
rect 155 501 167 535
rect 109 495 167 501
rect 23 313 81 319
rect 121 313 155 495
rect 23 279 35 313
rect 69 279 155 313
rect 23 273 81 279
rect 0 55 286 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 286 55
rect 0 0 286 21
<< labels >>
rlabel metal1 136 470 136 470 1 Y
port 1 n
rlabel metal1 64 666 64 666 1 A
port 2 n
rlabel metal1 212 592 212 592 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1284 68 1284 1 vdd
<< end >>
