* File: sky130_osu_sc_18T_ls__dlat_l.spice
* Created: Fri Nov 12 14:16:47 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_18T_ls__dlat_l.pex.spice"
.subckt sky130_osu_sc_18T_ls__dlat_l  GND VDD D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1002 A_115_115# N_D_M1002_g N_GND_M1002_s N_GND_M1002_b NSHORT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=5.988 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1013 N_D_M1013_d N_CK_M1013_g A_115_115# N_GND_M1002_b NSHORT L=0.15 W=1
+ AD=0.225 AS=0.105 PD=1.45 PS=1.21 NRD=10.188 NRS=5.988 M=1 R=6.66667
+ SA=75000.5 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1010 A_307_115# N_A_157_445#_M1010_g N_D_M1013_d N_GND_M1002_b NSHORT L=0.15
+ W=1 AD=0.105 AS=0.225 PD=1.21 PS=1.45 NRD=5.988 NRS=10.188 M=1 R=6.66667
+ SA=75001.1 SB=75001 A=0.15 P=2.3 MULT=1
MM1003 N_GND_M1003_d N_A_349_89#_M1003_g A_307_115# N_GND_M1002_b NSHORT L=0.15
+ W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=5.988 M=1 R=6.66667 SA=75001.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_157_445#_M1005_d N_CK_M1005_g N_GND_M1003_d N_GND_M1002_b NSHORT
+ L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_349_89#_M1006_d N_D_M1006_g N_GND_M1006_s N_GND_M1002_b NSHORT L=0.15
+ W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_GND_M1007_d N_A_349_89#_M1007_g N_QN_M1007_s N_GND_M1002_b NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_Q_M1009_d N_QN_M1009_g N_GND_M1007_d N_GND_M1002_b NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 A_115_617# N_D_M1014_g N_VDD_M1014_s N_VDD_M1014_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.2702 NRS=0 M=1 R=20 SA=75000.2
+ SB=75001.9 A=0.45 P=6.3 MULT=1
MM1011 N_D_M1011_d N_A_157_445#_M1011_g A_115_617# N_VDD_M1014_b PHIGHVT L=0.15
+ W=3 AD=0.675 AS=0.315 PD=3.45 PS=3.21 NRD=5.5751 NRS=3.2702 M=1 R=20
+ SA=75000.5 SB=75001.6 A=0.45 P=6.3 MULT=1
MM1015 A_307_617# N_CK_M1015_g N_D_M1011_d N_VDD_M1014_b PHIGHVT L=0.15 W=3
+ AD=0.315 AS=0.675 PD=3.21 PS=3.45 NRD=3.2702 NRS=5.5751 M=1 R=20 SA=75001.1
+ SB=75001 A=0.45 P=6.3 MULT=1
MM1000 N_VDD_M1000_d N_A_349_89#_M1000_g A_307_617# N_VDD_M1014_b PHIGHVT L=0.15
+ W=3 AD=0.42 AS=0.315 PD=3.28 PS=3.21 NRD=0 NRS=3.2702 M=1 R=20 SA=75001.5
+ SB=75000.6 A=0.45 P=6.3 MULT=1
MM1008 N_A_157_445#_M1008_d N_CK_M1008_g N_VDD_M1000_d N_VDD_M1014_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=20 SA=75001.9
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1001 N_A_349_89#_M1001_d N_D_M1001_g N_VDD_M1001_s N_VDD_M1014_b PHIGHVT
+ L=0.15 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.2 A=0.45 P=6.3 MULT=1
MM1012 N_VDD_M1012_d N_A_349_89#_M1012_g N_QN_M1012_s N_VDD_M1014_b PHIGHVT
+ L=0.15 W=2 AD=0.28 AS=0.53 PD=2.28 PS=4.53 NRD=0 NRS=0 M=1 R=13.3333
+ SA=75000.2 SB=75000.6 A=0.3 P=4.3 MULT=1
MM1004 N_Q_M1004_d N_QN_M1004_g N_VDD_M1012_d N_VDD_M1014_b PHIGHVT L=0.15 W=2
+ AD=0.53 AS=0.28 PD=4.53 PS=2.28 NRD=0 NRS=0 M=1 R=13.3333 SA=75000.6
+ SB=75000.2 A=0.3 P=4.3 MULT=1
DX16_noxref N_GND_M1002_b N_VDD_M1014_b NWDIODE A=19.551 P=17.89
pX17_noxref noxref_13 D D PROBETYPE=1
pX18_noxref noxref_14 CK CK PROBETYPE=1
pX19_noxref noxref_15 QN QN PROBETYPE=1
pX20_noxref noxref_16 Q Q PROBETYPE=1
c_753 A_115_617# 0 1.57671e-19 $X=0.575 $Y=3.085
*
.include "sky130_osu_sc_18T_ls__dlat_l.pxi.spice"
*
.ends
*
*
