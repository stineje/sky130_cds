* File: sky130_osu_sc_18T_ls__aoi22_l.pex.spice
* Created: Thu Oct 29 17:34:25 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%GND 1 2 19 23 27 31 37 39
c44 19 0 6.36774e-20 $X=-0.045 $Y=0
r45 37 39 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.7 $Y2=0.152
r46 31 32 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=0.152
+ $X2=1.91 $Y2=0.152
r47 25 32 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.152
r48 25 27 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.91 $Y=0.305
+ $X2=1.91 $Y2=0.825
r49 21 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.825
r50 19 21 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r51 19 42 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r52 19 31 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.825 $Y2=0.152
r53 19 42 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r54 19 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=0.17 $X2=1.7
+ $Y2=0.17
r55 19 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r56 2 27 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.77
+ $Y=0.575 $X2=1.91 $Y2=0.825
r57 1 23 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%VDD 1 13 17 22 25 30 39
r30 37 39 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r31 30 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.7 $Y=6.49 $X2=1.7
+ $Y2=6.49
r32 25 30 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=1.7 $Y2=6.507
r33 25 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r34 22 34 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r35 22 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r36 21 37 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r37 21 23 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r38 17 20 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.69 $Y=4.475
+ $X2=0.69 $Y2=5.835
r39 15 23 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r40 15 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r41 13 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r42 13 37 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r43 13 34 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r44 1 20 240 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r45 1 17 240 $w=1.7e-07 $l=1.45832e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.475
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%A0 2 3 5 8 12 15 22 24
c35 8 0 6.36774e-20 $X=0.475 $Y=4.585
r36 23 24 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.385 $Y=2.765
+ $X2=0.475 $Y2=2.765
r37 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=2.765 $X2=0.385 $Y2=2.765
r38 19 23 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.295 $Y=2.765
+ $X2=0.385 $Y2=2.765
r39 17 22 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.385 $Y2=2.765
r40 15 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.385 $Y=3.33
+ $X2=0.385 $Y2=3.33
r41 10 12 83.4231 $w=1.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.295 $Y=1.77
+ $X2=0.475 $Y2=1.77
r42 6 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=2.765
r43 6 8 864.011 $w=1.5e-07 $l=1.685e-06 $layer=POLY_cond $X=0.475 $Y=2.9
+ $X2=0.475 $Y2=4.585
r44 3 12 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.475 $Y=1.69 $X2=0.475
+ $Y2=1.77
r45 3 5 197.62 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.475 $Y=1.69
+ $X2=0.475 $Y2=1.075
r46 2 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.295 $Y=2.63
+ $X2=0.295 $Y2=2.765
r47 1 10 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.295 $Y=1.85 $X2=0.295
+ $Y2=1.77
r48 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.295 $Y=1.85
+ $X2=0.295 $Y2=2.63
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%A1 3 5 7 10 15
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=2.255 $X2=0.725 $Y2=2.255
r44 12 15 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.725 $Y=2.96
+ $X2=0.725 $Y2=2.255
r45 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=2.96
+ $X2=0.725 $Y2=2.96
r46 5 16 63.0864 $w=2.95e-07 $l=3.7229e-07 $layer=POLY_cond $X=0.905 $Y=2.57
+ $X2=0.78 $Y2=2.255
r47 5 7 1033.22 $w=1.5e-07 $l=2.015e-06 $layer=POLY_cond $X=0.905 $Y=2.57
+ $X2=0.905 $Y2=4.585
r48 1 16 38.578 $w=2.95e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.835 $Y=2.09
+ $X2=0.78 $Y2=2.255
r49 1 3 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=0.835 $Y=2.09
+ $X2=0.835 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%B0 3 7 9 13 15 17
r44 15 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.165 $Y=2.59
+ $X2=1.165 $Y2=2.59
r45 13 21 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.9
+ $X2=1.265 $Y2=2.065
r46 13 20 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.9
+ $X2=1.265 $Y2=1.735
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.9 $X2=1.255 $Y2=1.9
r48 10 17 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.165 $Y=2.065
+ $X2=1.165 $Y2=2.59
r49 9 12 3.63576 $w=3.02e-07 $l=9e-08 $layer=LI1_cond $X=1.165 $Y=1.9 $X2=1.255
+ $Y2=1.9
r50 9 10 4.10007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=1.9
+ $X2=1.165 $Y2=2.065
r51 7 21 1292.17 $w=1.5e-07 $l=2.52e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.065
r52 3 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=1.735
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%B1 3 7 10 12 15
r26 15 18 26.0127 $w=3.15e-07 $l=1.7e-07 $layer=POLY_cond $X=1.765 $Y=2.205
+ $X2=1.935 $Y2=2.205
r27 14 15 10.7111 $w=3.15e-07 $l=7e-08 $layer=POLY_cond $X=1.695 $Y=2.205
+ $X2=1.765 $Y2=2.205
r28 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=2.225 $X2=1.935 $Y2=2.225
r29 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.935 $Y=2.225
+ $X2=1.935 $Y2=2.225
r30 5 15 20.1192 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.765 $Y=2.39
+ $X2=1.765 $Y2=2.205
r31 5 7 1125.52 $w=1.5e-07 $l=2.195e-06 $layer=POLY_cond $X=1.765 $Y=2.39
+ $X2=1.765 $Y2=4.585
r32 1 14 20.1192 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.695 $Y=2.02
+ $X2=1.695 $Y2=2.205
r33 1 3 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.695 $Y=2.02
+ $X2=1.695 $Y2=1.075
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%A_27_617# 1 2 3 12 16 17 24 25
r23 28 31 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.98 $Y=4.135
+ $X2=1.98 $Y2=5.835
r24 26 31 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.98 $Y=5.915 $X2=1.98
+ $Y2=5.835
r25 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.895 $Y=6
+ $X2=1.98 $Y2=5.915
r26 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=6 $X2=1.205
+ $Y2=6
r27 21 23 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=1.12 $Y=4.135
+ $X2=1.12 $Y2=5.835
r28 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=5.915
+ $X2=1.205 $Y2=6
r29 19 23 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=5.915 $X2=1.12
+ $Y2=5.835
r30 18 21 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=4.055 $X2=1.12
+ $Y2=4.135
r31 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.97
+ $X2=1.12 $Y2=4.055
r32 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.97
+ $X2=0.345 $Y2=3.97
r33 12 14 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.26 $Y=4.135
+ $X2=0.26 $Y2=5.835
r34 10 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=4.055
+ $X2=0.345 $Y2=3.97
r35 10 12 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=4.055 $X2=0.26
+ $Y2=4.135
r36 3 31 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r37 3 28 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=4.135
r38 2 23 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r39 2 21 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=4.135
r40 1 14 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r41 1 12 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__AOI22_L%Y 1 2 9 16 17 21 28 29 33
c40 21 0 5.84789e-20 $X=1.605 $Y=1.7
r41 28 30 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.595 $Y=1.85
+ $X2=1.595 $Y2=1.735
r42 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.595 $Y=1.85
+ $X2=1.595 $Y2=1.85
r43 25 33 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.085 $Y=1.48
+ $X2=1.085 $Y2=0.825
r44 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.085 $Y=1.48
+ $X2=1.085 $Y2=1.48
r45 21 30 0.0337009 $w=1.7e-07 $l=3.5e-08 $layer=MET1_cond $X=1.605 $Y=1.7
+ $X2=1.605 $Y2=1.735
r46 18 21 0.129989 $w=1.7e-07 $l=1.35e-07 $layer=MET1_cond $X=1.605 $Y=1.565
+ $X2=1.605 $Y2=1.7
r47 17 24 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.23 $Y=1.48
+ $X2=1.085 $Y2=1.48
r48 16 18 0.0698411 $w=1.7e-07 $l=1.20208e-07 $layer=MET1_cond $X=1.52 $Y=1.48
+ $X2=1.605 $Y2=1.565
r49 16 17 0.279236 $w=1.7e-07 $l=2.9e-07 $layer=MET1_cond $X=1.52 $Y=1.48
+ $X2=1.23 $Y2=1.48
r50 14 29 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.595 $Y=3.16
+ $X2=1.595 $Y2=1.85
r51 14 15 9.11234 $w=2.13e-07 $l=1.7e-07 $layer=LI1_cond $X=1.572 $Y=3.16
+ $X2=1.572 $Y2=3.33
r52 9 11 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=5.495
r53 9 15 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.55 $Y=4.135
+ $X2=1.55 $Y2=3.33
r54 2 11 240 $w=1.7e-07 $l=2.47901e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.495
r55 2 9 240 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=4.135
r56 1 33 91 $w=1.7e-07 $l=3.2596e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.085 $Y2=0.825
.ends

