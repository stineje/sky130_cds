magic
tech sky130A
magscale 1 2
timestamp 1612373655
<< nwell >>
rect -9 529 374 1119
<< nmoslvt >>
rect 80 115 110 243
rect 166 115 196 243
rect 252 115 282 243
<< pmos >>
rect 80 565 110 965
rect 166 565 196 965
rect 252 565 282 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 166 243
rect 110 131 121 215
rect 155 131 166 215
rect 110 115 166 131
rect 196 215 252 243
rect 196 131 207 215
rect 241 131 252 215
rect 196 115 252 131
rect 282 215 335 243
rect 282 131 293 215
rect 327 131 335 215
rect 282 115 335 131
<< pdiff >>
rect 27 949 80 965
rect 27 673 35 949
rect 69 673 80 949
rect 27 565 80 673
rect 110 565 166 965
rect 196 949 252 965
rect 196 741 207 949
rect 241 741 252 949
rect 196 565 252 741
rect 282 949 335 965
rect 282 605 293 949
rect 327 605 335 949
rect 282 565 335 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
rect 207 131 241 215
rect 293 131 327 215
<< pdiffc >>
rect 35 673 69 949
rect 207 741 241 949
rect 293 605 327 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
rect 163 27 187 61
rect 221 27 245 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
rect 163 1049 187 1083
rect 221 1049 245 1083
<< psubdiffcont >>
rect 51 27 85 61
rect 187 27 221 61
<< nsubdiffcont >>
rect 51 1049 85 1083
rect 187 1049 221 1083
<< poly >>
rect 80 965 110 991
rect 166 965 196 991
rect 252 965 282 991
rect 80 516 110 565
rect 27 500 110 516
rect 27 466 37 500
rect 71 466 110 500
rect 27 450 110 466
rect 166 458 196 565
rect 252 540 282 565
rect 252 510 289 540
rect 80 243 110 450
rect 163 442 217 458
rect 163 408 173 442
rect 207 408 217 442
rect 163 392 217 408
rect 166 243 196 392
rect 259 368 289 510
rect 259 352 313 368
rect 259 332 269 352
rect 252 318 269 332
rect 303 318 313 352
rect 252 302 313 318
rect 252 243 282 302
rect 80 89 110 115
rect 166 89 196 115
rect 252 89 282 115
<< polycont >>
rect 37 466 71 500
rect 173 408 207 442
rect 269 318 303 352
<< locali >>
rect 0 1089 374 1110
rect 0 1049 51 1089
rect 85 1049 187 1089
rect 221 1049 374 1089
rect 35 949 69 965
rect 207 949 241 1049
rect 207 725 241 741
rect 293 949 327 965
rect 69 673 139 691
rect 35 657 139 673
rect 37 500 71 523
rect 37 450 71 466
rect 105 352 139 657
rect 173 442 207 597
rect 293 483 327 605
rect 173 392 207 408
rect 105 318 269 352
rect 303 318 319 352
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 318
rect 121 115 155 131
rect 207 215 241 231
rect 207 61 241 131
rect 293 215 327 227
rect 293 115 327 131
rect 0 21 51 61
rect 85 21 187 61
rect 221 21 374 61
rect 0 0 374 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 187 1083 221 1089
rect 187 1055 221 1083
rect 37 523 71 557
rect 173 597 207 631
rect 293 449 327 483
rect 293 227 327 261
rect 51 27 85 55
rect 51 21 85 27
rect 187 27 221 55
rect 187 21 221 27
<< metal1 >>
rect 0 1089 374 1110
rect 0 1055 51 1089
rect 85 1055 187 1089
rect 221 1055 374 1089
rect 0 1049 374 1055
rect 161 631 219 637
rect 140 597 173 631
rect 207 597 219 631
rect 161 591 219 597
rect 25 557 83 563
rect 25 523 37 557
rect 71 523 105 557
rect 25 517 83 523
rect 281 483 339 489
rect 281 449 293 483
rect 327 449 339 483
rect 281 443 339 449
rect 293 267 327 443
rect 281 261 339 267
rect 281 227 293 261
rect 327 227 339 261
rect 281 221 339 227
rect 0 55 374 61
rect 0 21 51 55
rect 85 21 187 55
rect 221 21 374 55
rect 0 0 374 21
<< labels >>
rlabel metal1 311 392 311 392 1 Y
port 1 n
rlabel viali 190 614 190 614 1 A
port 2 n
rlabel viali 54 540 54 540 1 B
port 3 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
