* File: sky130_osu_sc_18T_ms__tiehi.spice
* Created: Thu Oct 29 17:31:45 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* 
.include "sky130_osu_sc_18T_ms__tiehi.pex.spice"
.subckt sky130_osu_sc_18T_ms__tiehi  GND VDD Y
* 
* Y	Y
* VDD	VDD
* GND	GND
MM1000 N_A_80_89#_M1000_d N_A_80_89#_M1000_g N_GND_M1000_s N_GND_M1000_b NSHORT
+ L=0.15 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A_80_89#_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT L=0.15
+ W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 M=1 R=20 SA=75000.2
+ SB=75000.2 A=0.45 P=6.3 MULT=1
DX2_noxref N_GND_M1000_b N_VDD_M1001_b NWDIODE A=3.952 P=9.68
pX3_noxref noxref_5 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_18T_ms__tiehi.pxi.spice"
*
.ends
*
*
