* File: sky130_osu_sc_15T_ms__and2_1.pex.spice
* Created: Fri Nov 12 14:40:03 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__AND2_1%GND 1 17 19 26 35 38
r36 35 38 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=1.02 $Y2=0.152
r37 24 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r38 17 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r39 17 24 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r40 17 19 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r41 17 19 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r42 1 26 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_1%VDD 1 2 17 21 25 32 40 42 45
r29 42 45 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r30 32 35 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=3.555
+ $X2=1.12 $Y2=4.575
r31 30 40 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r32 30 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.575
r33 28 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.02 $Y=5.36
+ $X2=1.02 $Y2=5.36
r34 26 39 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r35 26 28 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r36 25 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r37 25 28 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r38 21 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.895
+ $X2=0.26 $Y2=4.575
r39 19 39 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r40 19 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.575
r41 17 28 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r42 17 39 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r43 2 35 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r44 2 32 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.555
r45 1 24 400 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r46 1 21 400 $w=1.7e-07 $l=1.13077e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_1%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=3.07
+ $X2=0.275 $Y2=3.07
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.07
+ $X2=0.27 $Y2=3.07
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.505
+ $X2=0.27 $Y2=3.07
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.505 $X2=0.27 $Y2=2.505
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.505
+ $X2=0.475 $Y2=2.505
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=2.505
r38 5 7 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=3.825
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=2.505
r40 1 3 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_1%B 3 7 10 14 22
r41 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.7
+ $X2=0.955 $Y2=2.7
r42 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.7 $X2=0.95
+ $Y2=2.7
r43 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.165
+ $X2=0.95 $Y2=2.7
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.165 $X2=0.95 $Y2=2.165
r45 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2.33
r46 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2
r47 7 12 766.585 $w=1.5e-07 $l=1.495e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.33
r48 3 11 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=2
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_1%A_27_115# 1 3 11 15 16 18 19 24 26 27 32
+ 38 40 41 42
r69 41 42 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.305
+ $X2=0.65 $Y2=3.475
r70 36 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=0.61 $Y2=1.675
r71 36 38 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=1.43 $Y2=1.675
r72 32 34 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=3.555
+ $X2=0.69 $Y2=4.575
r73 32 42 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.555 $X2=0.69
+ $Y2=3.475
r74 28 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.76 $X2=0.61
+ $Y2=1.675
r75 28 41 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=3.305
r76 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.61 $Y2=1.675
r77 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.345 $Y2=1.675
r78 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.345 $Y2=1.675
r79 22 24 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.74
r80 21 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.675 $X2=1.43 $Y2=1.675
r81 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=2.55
+ $X2=1.352 $Y2=2.7
r82 16 21 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.412 $Y2=1.675
r83 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=2.55
r84 15 19 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=3.825
+ $X2=1.335 $Y2=2.7
r85 9 21 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.412 $Y2=1.675
r86 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.945
r87 3 34 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.575
r88 3 32 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.555
r89 1 24 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__AND2_1%Y 1 3 10 16 26 29 32
r35 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r36 24 26 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r37 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r38 23 26 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r39 19 21 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.215
+ $X2=1.55 $Y2=4.575
r40 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r41 16 19 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=3.215
r42 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r43 10 13 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.22
r44 3 21 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.575
r45 3 19 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.215
r46 1 10 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

