* File: sky130_osu_sc_12T_hs__buf_l.pxi.spice
* Created: Fri Nov 12 15:08:45 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__BUF_L%GND N_GND_M1002_d N_GND_M1002_b N_GND_c_2_p
+ N_GND_c_3_p GND N_GND_c_4_p PM_SKY130_OSU_SC_12T_HS__BUF_L%GND
x_PM_SKY130_OSU_SC_12T_HS__BUF_L%VDD N_VDD_M1001_d N_VDD_M1001_b N_VDD_c_28_p
+ N_VDD_c_29_p N_VDD_c_36_p VDD N_VDD_c_30_p PM_SKY130_OSU_SC_12T_HS__BUF_L%VDD
x_PM_SKY130_OSU_SC_12T_HS__BUF_L%A N_A_M1002_g N_A_M1001_g N_A_c_51_n N_A_c_52_n
+ A PM_SKY130_OSU_SC_12T_HS__BUF_L%A
x_PM_SKY130_OSU_SC_12T_HS__BUF_L%A_27_115# N_A_27_115#_M1002_s
+ N_A_27_115#_M1001_s N_A_27_115#_M1000_g N_A_27_115#_c_98_n N_A_27_115#_M1003_g
+ N_A_27_115#_c_88_n N_A_27_115#_c_89_n N_A_27_115#_c_90_n N_A_27_115#_c_91_n
+ N_A_27_115#_c_94_n N_A_27_115#_c_95_n N_A_27_115#_c_96_n N_A_27_115#_c_97_n
+ PM_SKY130_OSU_SC_12T_HS__BUF_L%A_27_115#
x_PM_SKY130_OSU_SC_12T_HS__BUF_L%Y N_Y_M1000_d N_Y_M1003_d N_Y_c_138_n
+ N_Y_c_143_n Y N_Y_c_141_n N_Y_c_142_n PM_SKY130_OSU_SC_12T_HS__BUF_L%Y
cc_1 N_GND_M1002_b N_A_M1002_g 0.0853601f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.785
cc_2 N_GND_c_2_p N_A_M1002_g 0.00606474f $X=0.605 $Y=0.152 $X2=0.475 $Y2=0.785
cc_3 N_GND_c_3_p N_A_M1002_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.475 $Y2=0.785
cc_4 N_GND_c_4_p N_A_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.785
cc_5 N_GND_M1002_b N_A_M1001_g 0.0171588f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.445
cc_6 N_GND_M1002_b N_A_c_51_n 0.0409987f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.37
cc_7 N_GND_M1002_b N_A_c_52_n 0.00399069f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.37
cc_8 N_GND_M1002_b A 0.00826358f $X=-0.045 $Y=0 $X2=0.635 $Y2=2.48
cc_9 N_GND_M1002_b N_A_27_115#_M1000_g 0.0628823f $X=-0.045 $Y=0 $X2=0.905
+ $Y2=0.785
cc_10 N_GND_c_3_p N_A_27_115#_M1000_g 0.00308284f $X=0.69 $Y=0.74 $X2=0.905
+ $Y2=0.785
cc_11 N_GND_c_4_p N_A_27_115#_M1000_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905
+ $Y2=0.785
cc_12 N_GND_M1002_b N_A_27_115#_c_88_n 0.0597491f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.75
cc_13 N_GND_M1002_b N_A_27_115#_c_89_n 0.0562401f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=1.825
cc_14 N_GND_M1002_b N_A_27_115#_c_90_n 0.0168517f $X=-0.045 $Y=0 $X2=1.18
+ $Y2=2.825
cc_15 N_GND_M1002_b N_A_27_115#_c_91_n 0.0375616f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.74
cc_16 N_GND_c_2_p N_A_27_115#_c_91_n 0.00736239f $X=0.605 $Y=0.152 $X2=0.26
+ $Y2=0.74
cc_17 N_GND_c_4_p N_A_27_115#_c_91_n 0.00476261f $X=1.02 $Y=0.19 $X2=0.26
+ $Y2=0.74
cc_18 N_GND_M1002_b N_A_27_115#_c_94_n 0.041318f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=3.275
cc_19 N_GND_M1002_b N_A_27_115#_c_95_n 0.0155884f $X=-0.045 $Y=0 $X2=0.88
+ $Y2=1.825
cc_20 N_GND_M1002_b N_A_27_115#_c_96_n 0.0071553f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=1.825
cc_21 N_GND_M1002_b N_A_27_115#_c_97_n 0.00663593f $X=-0.045 $Y=0 $X2=0.965
+ $Y2=1.825
cc_22 N_GND_M1002_b N_Y_c_138_n 0.0302461f $X=-0.045 $Y=0 $X2=1.12 $Y2=0.74
cc_23 N_GND_c_4_p N_Y_c_138_n 0.00476261f $X=1.02 $Y=0.19 $X2=1.12 $Y2=0.74
cc_24 N_GND_M1002_b Y 0.0167208f $X=-0.045 $Y=0 $X2=1.07 $Y2=2.15
cc_25 N_GND_M1002_b N_Y_c_141_n 0.014537f $X=-0.045 $Y=0 $X2=1.12 $Y2=1.37
cc_26 N_GND_M1002_b N_Y_c_142_n 0.00512926f $X=-0.045 $Y=0 $X2=1.12 $Y2=2.85
cc_27 N_VDD_M1001_b N_A_M1001_g 0.0274536f $X=-0.045 $Y=2.795 $X2=0.475
+ $Y2=3.445
cc_28 N_VDD_c_28_p N_A_M1001_g 0.00606474f $X=0.605 $Y=4.287 $X2=0.475 $Y2=3.445
cc_29 N_VDD_c_29_p N_A_M1001_g 0.00354579f $X=0.69 $Y=3.275 $X2=0.475 $Y2=3.445
cc_30 N_VDD_c_30_p N_A_M1001_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.445
cc_31 N_VDD_c_29_p N_A_c_51_n 0.00204209f $X=0.69 $Y=3.275 $X2=0.635 $Y2=2.37
cc_32 N_VDD_c_29_p N_A_c_52_n 0.00287518f $X=0.69 $Y=3.275 $X2=0.635 $Y2=2.37
cc_33 N_VDD_c_29_p A 0.00514946f $X=0.69 $Y=3.275 $X2=0.635 $Y2=2.48
cc_34 N_VDD_M1001_b N_A_27_115#_c_98_n 0.0222851f $X=-0.045 $Y=2.795 $X2=0.905
+ $Y2=2.9
cc_35 N_VDD_c_29_p N_A_27_115#_c_98_n 0.00354579f $X=0.69 $Y=3.275 $X2=0.905
+ $Y2=2.9
cc_36 N_VDD_c_36_p N_A_27_115#_c_98_n 0.00606474f $X=1.02 $Y=4.22 $X2=0.905
+ $Y2=2.9
cc_37 N_VDD_c_30_p N_A_27_115#_c_98_n 0.00468827f $X=1.02 $Y=4.25 $X2=0.905
+ $Y2=2.9
cc_38 N_VDD_M1001_b N_A_27_115#_c_90_n 0.0187971f $X=-0.045 $Y=2.795 $X2=1.18
+ $Y2=2.825
cc_39 N_VDD_M1001_b N_A_27_115#_c_94_n 0.0129707f $X=-0.045 $Y=2.795 $X2=0.26
+ $Y2=3.275
cc_40 N_VDD_c_28_p N_A_27_115#_c_94_n 0.00736239f $X=0.605 $Y=4.287 $X2=0.26
+ $Y2=3.275
cc_41 N_VDD_c_30_p N_A_27_115#_c_94_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26
+ $Y2=3.275
cc_42 N_VDD_M1001_b N_Y_c_143_n 0.00582211f $X=-0.045 $Y=2.795 $X2=1.12 $Y2=2.85
cc_43 N_VDD_c_36_p N_Y_c_143_n 0.00736239f $X=1.02 $Y=4.22 $X2=1.12 $Y2=2.85
cc_44 N_VDD_c_30_p N_Y_c_143_n 0.00476261f $X=1.02 $Y=4.25 $X2=1.12 $Y2=2.85
cc_45 N_VDD_M1001_b N_Y_c_142_n 0.0107503f $X=-0.045 $Y=2.795 $X2=1.12 $Y2=2.85
cc_46 N_A_M1002_g N_A_27_115#_M1000_g 0.0502049f $X=0.475 $Y=0.785 $X2=0.905
+ $Y2=0.785
cc_47 N_A_M1002_g N_A_27_115#_c_88_n 0.00260138f $X=0.475 $Y=0.785 $X2=1.18
+ $Y2=2.75
cc_48 N_A_M1001_g N_A_27_115#_c_88_n 0.00264714f $X=0.475 $Y=3.445 $X2=1.18
+ $Y2=2.75
cc_49 N_A_c_51_n N_A_27_115#_c_88_n 0.0138474f $X=0.635 $Y=2.37 $X2=1.18
+ $Y2=2.75
cc_50 N_A_c_52_n N_A_27_115#_c_88_n 0.00245678f $X=0.635 $Y=2.37 $X2=1.18
+ $Y2=2.75
cc_51 A N_A_27_115#_c_88_n 6.60003e-19 $X=0.635 $Y=2.48 $X2=1.18 $Y2=2.75
cc_52 N_A_M1001_g N_A_27_115#_c_90_n 0.0204687f $X=0.475 $Y=3.445 $X2=1.18
+ $Y2=2.825
cc_53 N_A_M1002_g N_A_27_115#_c_91_n 0.0290598f $X=0.475 $Y=0.785 $X2=0.26
+ $Y2=0.74
cc_54 N_A_M1002_g N_A_27_115#_c_94_n 0.0390158f $X=0.475 $Y=0.785 $X2=0.26
+ $Y2=3.275
cc_55 N_A_c_52_n N_A_27_115#_c_94_n 0.0210234f $X=0.635 $Y=2.37 $X2=0.26
+ $Y2=3.275
cc_56 A N_A_27_115#_c_94_n 0.0155137f $X=0.635 $Y=2.48 $X2=0.26 $Y2=3.275
cc_57 N_A_M1002_g N_A_27_115#_c_95_n 0.0173663f $X=0.475 $Y=0.785 $X2=0.88
+ $Y2=1.825
cc_58 N_A_c_51_n N_A_27_115#_c_95_n 0.00273049f $X=0.635 $Y=2.37 $X2=0.88
+ $Y2=1.825
cc_59 N_A_c_52_n N_A_27_115#_c_95_n 0.00743028f $X=0.635 $Y=2.37 $X2=0.88
+ $Y2=1.825
cc_60 A N_A_27_115#_c_95_n 0.0090064f $X=0.635 $Y=2.48 $X2=0.88 $Y2=1.825
cc_61 N_A_M1002_g N_A_27_115#_c_97_n 6.59135e-19 $X=0.475 $Y=0.785 $X2=0.965
+ $Y2=1.825
cc_62 N_A_M1001_g N_Y_c_143_n 9.433e-19 $X=0.475 $Y=3.445 $X2=1.12 $Y2=2.85
cc_63 N_A_M1002_g Y 0.00310306f $X=0.475 $Y=0.785 $X2=1.07 $Y2=2.15
cc_64 N_A_M1001_g Y 0.00217977f $X=0.475 $Y=3.445 $X2=1.07 $Y2=2.15
cc_65 N_A_c_51_n Y 0.00257172f $X=0.635 $Y=2.37 $X2=1.07 $Y2=2.15
cc_66 N_A_c_52_n Y 0.00824365f $X=0.635 $Y=2.37 $X2=1.07 $Y2=2.15
cc_67 A Y 0.0185956f $X=0.635 $Y=2.48 $X2=1.07 $Y2=2.15
cc_68 N_A_M1002_g N_Y_c_141_n 0.00102215f $X=0.475 $Y=0.785 $X2=1.12 $Y2=1.37
cc_69 N_A_M1001_g N_Y_c_142_n 0.00126023f $X=0.475 $Y=3.445 $X2=1.12 $Y2=2.85
cc_70 N_A_27_115#_M1000_g N_Y_c_138_n 0.0178582f $X=0.905 $Y=0.785 $X2=1.12
+ $Y2=0.74
cc_71 N_A_27_115#_c_89_n N_Y_c_138_n 0.00477112f $X=1.18 $Y=1.825 $X2=1.12
+ $Y2=0.74
cc_72 N_A_27_115#_c_97_n N_Y_c_138_n 7.50437e-19 $X=0.965 $Y=1.825 $X2=1.12
+ $Y2=0.74
cc_73 N_A_27_115#_c_98_n N_Y_c_143_n 0.00655682f $X=0.905 $Y=2.9 $X2=1.12
+ $Y2=2.85
cc_74 N_A_27_115#_c_90_n N_Y_c_143_n 0.0149803f $X=1.18 $Y=2.825 $X2=1.12
+ $Y2=2.85
cc_75 N_A_27_115#_M1000_g Y 0.00406656f $X=0.905 $Y=0.785 $X2=1.07 $Y2=2.15
cc_76 N_A_27_115#_c_88_n Y 0.0310322f $X=1.18 $Y=2.75 $X2=1.07 $Y2=2.15
cc_77 N_A_27_115#_c_89_n Y 0.0161039f $X=1.18 $Y=1.825 $X2=1.07 $Y2=2.15
cc_78 N_A_27_115#_c_95_n Y 8.73078e-19 $X=0.88 $Y=1.825 $X2=1.07 $Y2=2.15
cc_79 N_A_27_115#_c_97_n Y 0.0121742f $X=0.965 $Y=1.825 $X2=1.07 $Y2=2.15
cc_80 N_A_27_115#_M1000_g N_Y_c_141_n 0.00714414f $X=0.905 $Y=0.785 $X2=1.12
+ $Y2=1.37
cc_81 N_A_27_115#_c_89_n N_Y_c_141_n 0.0014753f $X=1.18 $Y=1.825 $X2=1.12
+ $Y2=1.37
cc_82 N_A_27_115#_c_97_n N_Y_c_141_n 0.00278861f $X=0.965 $Y=1.825 $X2=1.12
+ $Y2=1.37
cc_83 N_A_27_115#_c_98_n N_Y_c_142_n 0.00213138f $X=0.905 $Y=2.9 $X2=1.12
+ $Y2=2.85
cc_84 N_A_27_115#_c_88_n N_Y_c_142_n 0.00226191f $X=1.18 $Y=2.75 $X2=1.12
+ $Y2=2.85
cc_85 N_A_27_115#_c_90_n N_Y_c_142_n 0.00641643f $X=1.18 $Y=2.825 $X2=1.12
+ $Y2=2.85
