* File: sky130_osu_sc_12T_hs__and2_4.pxi.spice
* Created: Fri Nov 12 15:07:01 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__AND2_4%GND N_GND_M1002_d N_GND_M1009_s N_GND_M1011_s
+ N_GND_M1004_b N_GND_c_2_p N_GND_c_8_p N_GND_c_16_p N_GND_c_22_p N_GND_c_30_p
+ N_GND_c_36_p GND N_GND_c_3_p PM_SKY130_OSU_SC_12T_HS__AND2_4%GND
x_PM_SKY130_OSU_SC_12T_HS__AND2_4%VDD N_VDD_M1000_s N_VDD_M1007_d N_VDD_M1005_d
+ N_VDD_M1008_d N_VDD_M1000_b N_VDD_c_77_p N_VDD_c_78_p N_VDD_c_89_p
+ N_VDD_c_96_p N_VDD_c_102_p N_VDD_c_108_p N_VDD_c_113_p VDD N_VDD_c_79_p
+ PM_SKY130_OSU_SC_12T_HS__AND2_4%VDD
x_PM_SKY130_OSU_SC_12T_HS__AND2_4%A N_A_M1004_g N_A_M1000_g N_A_c_132_n
+ N_A_c_133_n A PM_SKY130_OSU_SC_12T_HS__AND2_4%A
x_PM_SKY130_OSU_SC_12T_HS__AND2_4%B N_B_M1002_g N_B_M1007_g N_B_c_166_n
+ N_B_c_167_n B PM_SKY130_OSU_SC_12T_HS__AND2_4%B
x_PM_SKY130_OSU_SC_12T_HS__AND2_4%A_27_115# N_A_27_115#_M1004_s
+ N_A_27_115#_M1000_d N_A_27_115#_M1001_g N_A_27_115#_c_239_n
+ N_A_27_115#_M1003_g N_A_27_115#_c_206_n N_A_27_115#_c_207_n
+ N_A_27_115#_M1009_g N_A_27_115#_c_244_n N_A_27_115#_M1005_g
+ N_A_27_115#_c_212_n N_A_27_115#_c_214_n N_A_27_115#_c_215_n
+ N_A_27_115#_M1010_g N_A_27_115#_c_251_n N_A_27_115#_M1006_g
+ N_A_27_115#_c_220_n N_A_27_115#_c_221_n N_A_27_115#_M1011_g
+ N_A_27_115#_c_256_n N_A_27_115#_M1008_g N_A_27_115#_c_226_n
+ N_A_27_115#_c_227_n N_A_27_115#_c_228_n N_A_27_115#_c_229_n
+ N_A_27_115#_c_230_n N_A_27_115#_c_233_n N_A_27_115#_c_234_n
+ N_A_27_115#_c_263_n N_A_27_115#_c_235_n N_A_27_115#_c_237_n
+ N_A_27_115#_c_238_n N_A_27_115#_c_279_n
+ PM_SKY130_OSU_SC_12T_HS__AND2_4%A_27_115#
x_PM_SKY130_OSU_SC_12T_HS__AND2_4%Y N_Y_M1001_d N_Y_M1010_d N_Y_M1003_s
+ N_Y_M1006_s N_Y_c_337_n N_Y_c_342_n N_Y_c_343_n N_Y_c_347_n N_Y_c_348_n
+ N_Y_c_351_n Y N_Y_c_353_n N_Y_c_357_n N_Y_c_358_n N_Y_c_361_n
+ PM_SKY130_OSU_SC_12T_HS__AND2_4%Y
cc_1 N_GND_M1004_b N_A_M1004_g 0.079001f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_A_M1004_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_A_M1004_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.475 $Y2=0.85
cc_4 N_GND_M1004_b N_A_c_132_n 0.042117f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.285
cc_5 N_GND_M1004_b N_A_c_133_n 0.00270174f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.285
cc_6 N_GND_M1004_b N_B_M1002_g 0.0444472f $X=-0.045 $Y=0 $X2=0.835 $Y2=0.85
cc_7 N_GND_c_2_p N_B_M1002_g 0.00606474f $X=0.965 $Y=0.152 $X2=0.835 $Y2=0.85
cc_8 N_GND_c_8_p N_B_M1002_g 0.00319969f $X=1.05 $Y=0.755 $X2=0.835 $Y2=0.85
cc_9 N_GND_c_3_p N_B_M1002_g 0.00468827f $X=2.38 $Y=0.19 $X2=0.835 $Y2=0.85
cc_10 N_GND_M1004_b N_B_M1007_g 0.0151186f $X=-0.045 $Y=0 $X2=0.905 $Y2=3.235
cc_11 N_GND_M1004_b N_B_c_166_n 0.0333619f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.945
cc_12 N_GND_M1004_b N_B_c_167_n 0.00382966f $X=-0.045 $Y=0 $X2=0.95 $Y2=1.945
cc_13 N_GND_M1004_b B 0.00536919f $X=-0.045 $Y=0 $X2=0.955 $Y2=2.48
cc_14 N_GND_M1004_b N_A_27_115#_M1001_g 0.0199994f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=0.85
cc_15 N_GND_c_8_p N_A_27_115#_M1001_g 0.00610843f $X=1.05 $Y=0.755 $X2=1.335
+ $Y2=0.85
cc_16 N_GND_c_16_p N_A_27_115#_M1001_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=0.85
cc_17 N_GND_c_3_p N_A_27_115#_M1001_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.335
+ $Y2=0.85
cc_18 N_GND_M1004_b N_A_27_115#_c_206_n 0.0470206f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.33
cc_19 N_GND_M1004_b N_A_27_115#_c_207_n 0.00954592f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.405
cc_20 N_GND_M1004_b N_A_27_115#_M1009_g 0.0187696f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=0.85
cc_21 N_GND_c_16_p N_A_27_115#_M1009_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=0.85
cc_22 N_GND_c_22_p N_A_27_115#_M1009_g 0.00311745f $X=1.98 $Y=0.755 $X2=1.765
+ $Y2=0.85
cc_23 N_GND_c_3_p N_A_27_115#_M1009_g 0.00468827f $X=2.38 $Y=0.19 $X2=1.765
+ $Y2=0.85
cc_24 N_GND_M1004_b N_A_27_115#_c_212_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.365
cc_25 N_GND_c_22_p N_A_27_115#_c_212_n 0.00256938f $X=1.98 $Y=0.755 $X2=2.12
+ $Y2=1.365
cc_26 N_GND_M1004_b N_A_27_115#_c_214_n 0.0448266f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.365
cc_27 N_GND_M1004_b N_A_27_115#_c_215_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.405
cc_28 N_GND_M1004_b N_A_27_115#_M1010_g 0.0187674f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=0.85
cc_29 N_GND_c_22_p N_A_27_115#_M1010_g 0.00311745f $X=1.98 $Y=0.755 $X2=2.195
+ $Y2=0.85
cc_30 N_GND_c_30_p N_A_27_115#_M1010_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=0.85
cc_31 N_GND_c_3_p N_A_27_115#_M1010_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.195
+ $Y2=0.85
cc_32 N_GND_M1004_b N_A_27_115#_c_220_n 0.0369419f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.365
cc_33 N_GND_M1004_b N_A_27_115#_c_221_n 0.0268552f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.405
cc_34 N_GND_M1004_b N_A_27_115#_M1011_g 0.0241608f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=0.85
cc_35 N_GND_c_30_p N_A_27_115#_M1011_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=0.85
cc_36 N_GND_c_36_p N_A_27_115#_M1011_g 0.00502587f $X=2.84 $Y=0.755 $X2=2.625
+ $Y2=0.85
cc_37 N_GND_c_3_p N_A_27_115#_M1011_g 0.00468827f $X=2.38 $Y=0.19 $X2=2.625
+ $Y2=0.85
cc_38 N_GND_M1004_b N_A_27_115#_c_226_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.405
cc_39 N_GND_M1004_b N_A_27_115#_c_227_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.405
cc_40 N_GND_M1004_b N_A_27_115#_c_228_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.365
cc_41 N_GND_M1004_b N_A_27_115#_c_229_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.405
cc_42 N_GND_M1004_b N_A_27_115#_c_230_n 0.0128494f $X=-0.045 $Y=0 $X2=0.26
+ $Y2=0.755
cc_43 N_GND_c_2_p N_A_27_115#_c_230_n 0.00736239f $X=0.965 $Y=0.152 $X2=0.26
+ $Y2=0.755
cc_44 N_GND_c_3_p N_A_27_115#_c_230_n 0.00476261f $X=2.38 $Y=0.19 $X2=0.26
+ $Y2=0.755
cc_45 N_GND_M1004_b N_A_27_115#_c_233_n 0.00258316f $X=-0.045 $Y=0 $X2=0.525
+ $Y2=1.455
cc_46 N_GND_M1004_b N_A_27_115#_c_234_n 0.00933193f $X=-0.045 $Y=0 $X2=0.345
+ $Y2=1.455
cc_47 N_GND_M1004_b N_A_27_115#_c_235_n 0.0230268f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.455
cc_48 N_GND_c_8_p N_A_27_115#_c_235_n 0.00704977f $X=1.05 $Y=0.755 $X2=1.43
+ $Y2=1.455
cc_49 N_GND_M1004_b N_A_27_115#_c_237_n 0.00590548f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=1.455
cc_50 N_GND_M1004_b N_A_27_115#_c_238_n 0.00587837f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=3.065
cc_51 N_GND_M1004_b N_Y_c_337_n 0.00154299f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.755
cc_52 N_GND_c_8_p N_Y_c_337_n 0.00806382f $X=1.05 $Y=0.755 $X2=1.55 $Y2=0.755
cc_53 N_GND_c_16_p N_Y_c_337_n 0.00722248f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.755
cc_54 N_GND_c_22_p N_Y_c_337_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=0.755
cc_55 N_GND_c_3_p N_Y_c_337_n 0.0047139f $X=2.38 $Y=0.19 $X2=1.55 $Y2=0.755
cc_56 N_GND_M1004_b N_Y_c_342_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.11
cc_57 N_GND_M1004_b N_Y_c_343_n 0.00154299f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.755
cc_58 N_GND_c_22_p N_Y_c_343_n 8.14297e-19 $X=1.98 $Y=0.755 $X2=2.41 $Y2=0.755
cc_59 N_GND_c_30_p N_Y_c_343_n 0.00718527f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.755
cc_60 N_GND_c_3_p N_Y_c_343_n 0.0047139f $X=2.38 $Y=0.19 $X2=2.41 $Y2=0.755
cc_61 N_GND_M1004_b N_Y_c_347_n 0.0152877f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.11
cc_62 N_GND_c_8_p N_Y_c_348_n 0.00127231f $X=1.05 $Y=0.755 $X2=1.55 $Y2=1.115
cc_63 N_GND_c_16_p N_Y_c_348_n 0.00245319f $X=1.895 $Y=0.152 $X2=1.55 $Y2=1.115
cc_64 N_GND_c_22_p N_Y_c_348_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=1.55 $Y2=1.115
cc_65 N_GND_M1004_b N_Y_c_351_n 0.00463624f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.995
cc_66 N_GND_M1004_b Y 0.0304285f $X=-0.045 $Y=0 $X2=1.555 $Y2=1.74
cc_67 N_GND_M1009_s N_Y_c_353_n 0.0100329f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1
cc_68 N_GND_c_16_p N_Y_c_353_n 0.0028844f $X=1.895 $Y=0.152 $X2=2.265 $Y2=1
cc_69 N_GND_c_22_p N_Y_c_353_n 0.0142303f $X=1.98 $Y=0.755 $X2=2.265 $Y2=1
cc_70 N_GND_c_30_p N_Y_c_353_n 0.0028844f $X=2.755 $Y=0.152 $X2=2.265 $Y2=1
cc_71 N_GND_M1004_b N_Y_c_357_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.11
cc_72 N_GND_c_22_p N_Y_c_358_n 7.53951e-19 $X=1.98 $Y=0.755 $X2=2.41 $Y2=1.115
cc_73 N_GND_c_30_p N_Y_c_358_n 0.00245319f $X=2.755 $Y=0.152 $X2=2.41 $Y2=1.115
cc_74 N_GND_c_36_p N_Y_c_358_n 0.00134236f $X=2.84 $Y=0.755 $X2=2.41 $Y2=1.115
cc_75 N_GND_M1004_b N_Y_c_361_n 0.0611971f $X=-0.045 $Y=0 $X2=2.41 $Y2=1.995
cc_76 N_VDD_M1000_b N_A_M1000_g 0.0189471f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_77 N_VDD_c_77_p N_A_M1000_g 0.00636672f $X=0.26 $Y=3.635 $X2=0.475 $Y2=3.235
cc_78 N_VDD_c_78_p N_A_M1000_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.475 $Y2=3.235
cc_79 N_VDD_c_79_p N_A_M1000_g 0.00468827f $X=2.38 $Y=4.25 $X2=0.475 $Y2=3.235
cc_80 N_VDD_M1000_b N_A_c_132_n 0.0111025f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=2.285
cc_81 N_VDD_M1000_s N_A_c_133_n 0.0127298f $X=0.135 $Y=2.605 $X2=0.27 $Y2=2.285
cc_82 N_VDD_M1000_b N_A_c_133_n 0.00612103f $X=-0.045 $Y=2.425 $X2=0.27
+ $Y2=2.285
cc_83 N_VDD_c_77_p N_A_c_133_n 0.00370742f $X=0.26 $Y=3.635 $X2=0.27 $Y2=2.285
cc_84 N_VDD_M1000_s A 0.00742066f $X=0.135 $Y=2.605 $X2=0.275 $Y2=2.85
cc_85 N_VDD_M1000_b A 0.00970321f $X=-0.045 $Y=2.425 $X2=0.275 $Y2=2.85
cc_86 N_VDD_c_77_p A 0.00434783f $X=0.26 $Y=3.635 $X2=0.275 $Y2=2.85
cc_87 N_VDD_M1000_b N_B_M1007_g 0.0187476f $X=-0.045 $Y=2.425 $X2=0.905
+ $Y2=3.235
cc_88 N_VDD_c_78_p N_B_M1007_g 0.00606474f $X=1.035 $Y=4.287 $X2=0.905 $Y2=3.235
cc_89 N_VDD_c_89_p N_B_M1007_g 0.00337744f $X=1.12 $Y=3.295 $X2=0.905 $Y2=3.235
cc_90 N_VDD_c_79_p N_B_M1007_g 0.00468827f $X=2.38 $Y=4.25 $X2=0.905 $Y2=3.235
cc_91 N_VDD_M1000_b N_B_c_167_n 0.00170274f $X=-0.045 $Y=2.425 $X2=0.95
+ $Y2=1.945
cc_92 N_VDD_M1000_b B 0.00856863f $X=-0.045 $Y=2.425 $X2=0.955 $Y2=2.48
cc_93 N_VDD_c_89_p B 0.00240671f $X=1.12 $Y=3.295 $X2=0.955 $Y2=2.48
cc_94 N_VDD_M1000_b N_A_27_115#_c_239_n 0.017104f $X=-0.045 $Y=2.425 $X2=1.335
+ $Y2=2.48
cc_95 N_VDD_c_89_p N_A_27_115#_c_239_n 0.00337744f $X=1.12 $Y=3.295 $X2=1.335
+ $Y2=2.48
cc_96 N_VDD_c_96_p N_A_27_115#_c_239_n 0.00606474f $X=1.895 $Y=4.287 $X2=1.335
+ $Y2=2.48
cc_97 N_VDD_c_79_p N_A_27_115#_c_239_n 0.00468827f $X=2.38 $Y=4.25 $X2=1.335
+ $Y2=2.48
cc_98 N_VDD_M1000_b N_A_27_115#_c_207_n 0.00428234f $X=-0.045 $Y=2.425 $X2=1.69
+ $Y2=2.405
cc_99 N_VDD_M1000_b N_A_27_115#_c_244_n 0.017006f $X=-0.045 $Y=2.425 $X2=1.765
+ $Y2=2.48
cc_100 N_VDD_c_89_p N_A_27_115#_c_244_n 3.67508e-19 $X=1.12 $Y=3.295 $X2=1.765
+ $Y2=2.48
cc_101 N_VDD_c_96_p N_A_27_115#_c_244_n 0.00610567f $X=1.895 $Y=4.287 $X2=1.765
+ $Y2=2.48
cc_102 N_VDD_c_102_p N_A_27_115#_c_244_n 0.0035715f $X=1.98 $Y=2.955 $X2=1.765
+ $Y2=2.48
cc_103 N_VDD_c_79_p N_A_27_115#_c_244_n 0.00470215f $X=2.38 $Y=4.25 $X2=1.765
+ $Y2=2.48
cc_104 N_VDD_M1000_b N_A_27_115#_c_215_n 0.00396043f $X=-0.045 $Y=2.425 $X2=2.12
+ $Y2=2.405
cc_105 N_VDD_c_102_p N_A_27_115#_c_215_n 0.00379272f $X=1.98 $Y=2.955 $X2=2.12
+ $Y2=2.405
cc_106 N_VDD_M1000_b N_A_27_115#_c_251_n 0.0166898f $X=-0.045 $Y=2.425 $X2=2.195
+ $Y2=2.48
cc_107 N_VDD_c_102_p N_A_27_115#_c_251_n 0.00337744f $X=1.98 $Y=2.955 $X2=2.195
+ $Y2=2.48
cc_108 N_VDD_c_108_p N_A_27_115#_c_251_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.195
+ $Y2=2.48
cc_109 N_VDD_c_79_p N_A_27_115#_c_251_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.195
+ $Y2=2.48
cc_110 N_VDD_M1000_b N_A_27_115#_c_221_n 0.00840215f $X=-0.045 $Y=2.425 $X2=2.55
+ $Y2=2.405
cc_111 N_VDD_M1000_b N_A_27_115#_c_256_n 0.0209036f $X=-0.045 $Y=2.425 $X2=2.625
+ $Y2=2.48
cc_112 N_VDD_c_108_p N_A_27_115#_c_256_n 0.00606474f $X=2.755 $Y=4.287 $X2=2.625
+ $Y2=2.48
cc_113 N_VDD_c_113_p N_A_27_115#_c_256_n 0.00636672f $X=2.84 $Y=2.955 $X2=2.625
+ $Y2=2.48
cc_114 N_VDD_c_79_p N_A_27_115#_c_256_n 0.00468827f $X=2.38 $Y=4.25 $X2=2.625
+ $Y2=2.48
cc_115 N_VDD_M1000_b N_A_27_115#_c_226_n 0.0021704f $X=-0.045 $Y=2.425 $X2=1.352
+ $Y2=2.405
cc_116 N_VDD_M1000_b N_A_27_115#_c_227_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=1.765 $Y2=2.405
cc_117 N_VDD_M1000_b N_A_27_115#_c_229_n 8.75564e-19 $X=-0.045 $Y=2.425
+ $X2=2.195 $Y2=2.405
cc_118 N_VDD_M1000_b N_A_27_115#_c_263_n 0.00155118f $X=-0.045 $Y=2.425 $X2=0.69
+ $Y2=3.295
cc_119 N_VDD_c_78_p N_A_27_115#_c_263_n 0.0075556f $X=1.035 $Y=4.287 $X2=0.69
+ $Y2=3.295
cc_120 N_VDD_c_79_p N_A_27_115#_c_263_n 0.00475776f $X=2.38 $Y=4.25 $X2=0.69
+ $Y2=3.295
cc_121 N_VDD_M1000_b N_A_27_115#_c_238_n 8.22047e-19 $X=-0.045 $Y=2.425 $X2=0.65
+ $Y2=3.065
cc_122 N_VDD_M1000_b N_Y_c_342_n 0.00344954f $X=-0.045 $Y=2.425 $X2=1.55
+ $Y2=2.11
cc_123 N_VDD_c_96_p N_Y_c_342_n 0.00737727f $X=1.895 $Y=4.287 $X2=1.55 $Y2=2.11
cc_124 N_VDD_c_79_p N_Y_c_342_n 0.00475776f $X=2.38 $Y=4.25 $X2=1.55 $Y2=2.11
cc_125 N_VDD_M1000_b N_Y_c_347_n 0.00380347f $X=-0.045 $Y=2.425 $X2=2.41
+ $Y2=2.11
cc_126 N_VDD_c_108_p N_Y_c_347_n 0.00734006f $X=2.755 $Y=4.287 $X2=2.41 $Y2=2.11
cc_127 N_VDD_c_79_p N_Y_c_347_n 0.00475776f $X=2.38 $Y=4.25 $X2=2.41 $Y2=2.11
cc_128 N_VDD_c_102_p N_Y_c_357_n 0.00634153f $X=1.98 $Y=2.955 $X2=2.265 $Y2=2.11
cc_129 N_A_M1004_g N_B_M1002_g 0.101204f $X=0.475 $Y=0.85 $X2=0.835 $Y2=0.85
cc_130 N_A_M1004_g N_B_M1007_g 0.048305f $X=0.475 $Y=0.85 $X2=0.905 $Y2=3.235
cc_131 N_A_M1004_g N_B_c_167_n 7.8234e-19 $X=0.475 $Y=0.85 $X2=0.95 $Y2=1.945
cc_132 N_A_M1004_g N_A_27_115#_c_230_n 0.0128217f $X=0.475 $Y=0.85 $X2=0.26
+ $Y2=0.755
cc_133 N_A_M1004_g N_A_27_115#_c_233_n 0.0160984f $X=0.475 $Y=0.85 $X2=0.525
+ $Y2=1.455
cc_134 N_A_c_132_n N_A_27_115#_c_233_n 0.00117122f $X=0.475 $Y=2.285 $X2=0.525
+ $Y2=1.455
cc_135 N_A_c_133_n N_A_27_115#_c_233_n 2.65873e-19 $X=0.27 $Y=2.285 $X2=0.525
+ $Y2=1.455
cc_136 N_A_c_132_n N_A_27_115#_c_234_n 0.00133457f $X=0.475 $Y=2.285 $X2=0.345
+ $Y2=1.455
cc_137 N_A_c_133_n N_A_27_115#_c_234_n 0.0055861f $X=0.27 $Y=2.285 $X2=0.345
+ $Y2=1.455
cc_138 N_A_M1004_g N_A_27_115#_c_237_n 0.00322084f $X=0.475 $Y=0.85 $X2=0.61
+ $Y2=1.455
cc_139 N_A_M1004_g N_A_27_115#_c_238_n 0.0265302f $X=0.475 $Y=0.85 $X2=0.65
+ $Y2=3.065
cc_140 N_A_M1000_g N_A_27_115#_c_238_n 0.0140172f $X=0.475 $Y=3.235 $X2=0.65
+ $Y2=3.065
cc_141 N_A_c_132_n N_A_27_115#_c_238_n 0.00766302f $X=0.475 $Y=2.285 $X2=0.65
+ $Y2=3.065
cc_142 N_A_c_133_n N_A_27_115#_c_238_n 0.0456533f $X=0.27 $Y=2.285 $X2=0.65
+ $Y2=3.065
cc_143 A N_A_27_115#_c_238_n 0.00758489f $X=0.275 $Y=2.85 $X2=0.65 $Y2=3.065
cc_144 N_A_M1000_g N_A_27_115#_c_279_n 0.00865855f $X=0.475 $Y=3.235 $X2=0.65
+ $Y2=3.235
cc_145 N_B_M1002_g N_A_27_115#_M1001_g 0.0272101f $X=0.835 $Y=0.85 $X2=1.335
+ $Y2=0.85
cc_146 N_B_M1007_g N_A_27_115#_c_206_n 0.00773101f $X=0.905 $Y=3.235 $X2=1.37
+ $Y2=2.33
cc_147 N_B_c_166_n N_A_27_115#_c_206_n 0.0206104f $X=0.95 $Y=1.945 $X2=1.37
+ $Y2=2.33
cc_148 N_B_c_167_n N_A_27_115#_c_206_n 0.0033451f $X=0.95 $Y=1.945 $X2=1.37
+ $Y2=2.33
cc_149 N_B_M1002_g N_A_27_115#_c_214_n 0.0104742f $X=0.835 $Y=0.85 $X2=1.84
+ $Y2=1.365
cc_150 N_B_M1007_g N_A_27_115#_c_226_n 0.0387792f $X=0.905 $Y=3.235 $X2=1.352
+ $Y2=2.405
cc_151 N_B_c_167_n N_A_27_115#_c_226_n 0.00173699f $X=0.95 $Y=1.945 $X2=1.352
+ $Y2=2.405
cc_152 B N_A_27_115#_c_226_n 0.00389258f $X=0.955 $Y=2.48 $X2=1.352 $Y2=2.405
cc_153 N_B_M1002_g N_A_27_115#_c_235_n 0.0182215f $X=0.835 $Y=0.85 $X2=1.43
+ $Y2=1.455
cc_154 N_B_c_166_n N_A_27_115#_c_235_n 0.00258465f $X=0.95 $Y=1.945 $X2=1.43
+ $Y2=1.455
cc_155 N_B_c_167_n N_A_27_115#_c_235_n 0.0101796f $X=0.95 $Y=1.945 $X2=1.43
+ $Y2=1.455
cc_156 N_B_M1002_g N_A_27_115#_c_238_n 0.00755919f $X=0.835 $Y=0.85 $X2=0.65
+ $Y2=3.065
cc_157 N_B_M1007_g N_A_27_115#_c_238_n 0.0133197f $X=0.905 $Y=3.235 $X2=0.65
+ $Y2=3.065
cc_158 N_B_c_167_n N_A_27_115#_c_238_n 0.0541375f $X=0.95 $Y=1.945 $X2=0.65
+ $Y2=3.065
cc_159 B N_A_27_115#_c_238_n 0.00866797f $X=0.955 $Y=2.48 $X2=0.65 $Y2=3.065
cc_160 B N_A_27_115#_c_279_n 0.00286715f $X=0.955 $Y=2.48 $X2=0.65 $Y2=3.235
cc_161 N_B_c_167_n N_Y_c_342_n 0.0149875f $X=0.95 $Y=1.945 $X2=1.55 $Y2=2.11
cc_162 B N_Y_c_342_n 0.00649253f $X=0.955 $Y=2.48 $X2=1.55 $Y2=2.11
cc_163 N_B_M1002_g N_Y_c_348_n 7.93934e-19 $X=0.835 $Y=0.85 $X2=1.55 $Y2=1.115
cc_164 N_B_c_166_n N_Y_c_351_n 5.85867e-19 $X=0.95 $Y=1.945 $X2=1.55 $Y2=1.995
cc_165 N_B_c_167_n N_Y_c_351_n 0.00592261f $X=0.95 $Y=1.945 $X2=1.55 $Y2=1.995
cc_166 N_B_M1002_g Y 6.71108e-19 $X=0.835 $Y=0.85 $X2=1.555 $Y2=1.74
cc_167 N_B_c_167_n Y 0.00695761f $X=0.95 $Y=1.945 $X2=1.555 $Y2=1.74
cc_168 N_A_27_115#_M1001_g N_Y_c_337_n 0.00184843f $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=0.755
cc_169 N_A_27_115#_M1009_g N_Y_c_337_n 0.00182852f $X=1.765 $Y=0.85 $X2=1.55
+ $Y2=0.755
cc_170 N_A_27_115#_c_214_n N_Y_c_337_n 0.0016986f $X=1.84 $Y=1.365 $X2=1.55
+ $Y2=0.755
cc_171 N_A_27_115#_c_235_n N_Y_c_337_n 0.00498892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=0.755
cc_172 N_A_27_115#_c_239_n N_Y_c_342_n 0.0026195f $X=1.335 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_173 N_A_27_115#_c_206_n N_Y_c_342_n 0.00744772f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=2.11
cc_174 N_A_27_115#_c_207_n N_Y_c_342_n 0.0167599f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=2.11
cc_175 N_A_27_115#_c_244_n N_Y_c_342_n 0.00375894f $X=1.765 $Y=2.48 $X2=1.55
+ $Y2=2.11
cc_176 N_A_27_115#_c_214_n N_Y_c_342_n 0.0013767f $X=1.84 $Y=1.365 $X2=1.55
+ $Y2=2.11
cc_177 N_A_27_115#_c_235_n N_Y_c_342_n 0.00273485f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=2.11
cc_178 N_A_27_115#_M1010_g N_Y_c_343_n 0.00182852f $X=2.195 $Y=0.85 $X2=2.41
+ $Y2=0.755
cc_179 N_A_27_115#_c_220_n N_Y_c_343_n 0.00274041f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=0.755
cc_180 N_A_27_115#_M1011_g N_Y_c_343_n 0.00182852f $X=2.625 $Y=0.85 $X2=2.41
+ $Y2=0.755
cc_181 N_A_27_115#_c_251_n N_Y_c_347_n 0.00375894f $X=2.195 $Y=2.48 $X2=2.41
+ $Y2=2.11
cc_182 N_A_27_115#_c_220_n N_Y_c_347_n 0.00250559f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=2.11
cc_183 N_A_27_115#_c_221_n N_Y_c_347_n 0.0206674f $X=2.55 $Y=2.405 $X2=2.41
+ $Y2=2.11
cc_184 N_A_27_115#_c_256_n N_Y_c_347_n 0.00375894f $X=2.625 $Y=2.48 $X2=2.41
+ $Y2=2.11
cc_185 N_A_27_115#_M1001_g N_Y_c_348_n 0.00493416f $X=1.335 $Y=0.85 $X2=1.55
+ $Y2=1.115
cc_186 N_A_27_115#_M1009_g N_Y_c_348_n 0.00198614f $X=1.765 $Y=0.85 $X2=1.55
+ $Y2=1.115
cc_187 N_A_27_115#_c_235_n N_Y_c_348_n 0.00238892f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1.115
cc_188 N_A_27_115#_c_206_n N_Y_c_351_n 0.00821104f $X=1.37 $Y=2.33 $X2=1.55
+ $Y2=1.995
cc_189 N_A_27_115#_c_207_n N_Y_c_351_n 0.00229755f $X=1.69 $Y=2.405 $X2=1.55
+ $Y2=1.995
cc_190 N_A_27_115#_c_214_n N_Y_c_351_n 0.00174847f $X=1.84 $Y=1.365 $X2=1.55
+ $Y2=1.995
cc_191 N_A_27_115#_c_235_n N_Y_c_351_n 0.00181779f $X=1.43 $Y=1.455 $X2=1.55
+ $Y2=1.995
cc_192 N_A_27_115#_M1001_g Y 0.00251111f $X=1.335 $Y=0.85 $X2=1.555 $Y2=1.74
cc_193 N_A_27_115#_c_206_n Y 0.00892438f $X=1.37 $Y=2.33 $X2=1.555 $Y2=1.74
cc_194 N_A_27_115#_M1009_g Y 0.00251111f $X=1.765 $Y=0.85 $X2=1.555 $Y2=1.74
cc_195 N_A_27_115#_c_214_n Y 0.0128645f $X=1.84 $Y=1.365 $X2=1.555 $Y2=1.74
cc_196 N_A_27_115#_c_235_n Y 0.0148238f $X=1.43 $Y=1.455 $X2=1.555 $Y2=1.74
cc_197 N_A_27_115#_M1009_g N_Y_c_353_n 0.00873177f $X=1.765 $Y=0.85 $X2=2.265
+ $Y2=1
cc_198 N_A_27_115#_c_212_n N_Y_c_353_n 0.00213861f $X=2.12 $Y=1.365 $X2=2.265
+ $Y2=1
cc_199 N_A_27_115#_M1010_g N_Y_c_353_n 0.00873177f $X=2.195 $Y=0.85 $X2=2.265
+ $Y2=1
cc_200 N_A_27_115#_c_214_n N_Y_c_357_n 0.0121767f $X=1.84 $Y=1.365 $X2=2.265
+ $Y2=2.11
cc_201 N_A_27_115#_c_227_n N_Y_c_357_n 0.0158479f $X=1.765 $Y=2.405 $X2=2.265
+ $Y2=2.11
cc_202 N_A_27_115#_M1010_g N_Y_c_358_n 0.00198614f $X=2.195 $Y=0.85 $X2=2.41
+ $Y2=1.115
cc_203 N_A_27_115#_M1011_g N_Y_c_358_n 0.00878256f $X=2.625 $Y=0.85 $X2=2.41
+ $Y2=1.115
cc_204 N_A_27_115#_M1010_g N_Y_c_361_n 0.00251111f $X=2.195 $Y=0.85 $X2=2.41
+ $Y2=1.995
cc_205 N_A_27_115#_c_220_n N_Y_c_361_n 0.0184054f $X=2.55 $Y=1.365 $X2=2.41
+ $Y2=1.995
cc_206 N_A_27_115#_M1011_g N_Y_c_361_n 0.00251111f $X=2.625 $Y=0.85 $X2=2.41
+ $Y2=1.995
cc_207 N_A_27_115#_c_228_n N_Y_c_361_n 0.00140336f $X=2.195 $Y=1.365 $X2=2.41
+ $Y2=1.995
cc_208 N_A_27_115#_c_229_n N_Y_c_361_n 0.00372651f $X=2.195 $Y=2.405 $X2=2.41
+ $Y2=1.995
