* File: sky130_osu_sc_18T_hs__ndlat_1.pex.spice
* Created: Thu Mar 10 17:10:18 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%GND 1 2 3 49 51 58 60 70 72 82 95 97 99
+ 101 103 107
c110 82 0 1.97615e-19 $X=4.365 $Y=0.825
r111 105 107 0.00465721 $w=3.05e-07 $l=1e-08 $layer=MET1_cond $X=4.42 $Y=0.152
+ $X2=4.43 $Y2=0.152
r112 103 105 0.323676 $w=3.05e-07 $l=6.95e-07 $layer=MET1_cond $X=3.725 $Y=0.152
+ $X2=4.42 $Y2=0.152
r113 101 103 0.312033 $w=3.05e-07 $l=6.7e-07 $layer=MET1_cond $X=3.055 $Y=0.152
+ $X2=3.725 $Y2=0.152
r114 99 101 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=2.375 $Y=0.152
+ $X2=3.055 $Y2=0.152
r115 97 99 0.321348 $w=3.05e-07 $l=6.9e-07 $layer=MET1_cond $X=1.685 $Y=0.152
+ $X2=2.375 $Y2=0.152
r116 95 97 0.309705 $w=3.05e-07 $l=6.65e-07 $layer=MET1_cond $X=1.02 $Y=0.152
+ $X2=1.685 $Y2=0.152
r117 80 82 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.365 $Y=0.305
+ $X2=4.365 $Y2=0.825
r118 73 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.152
+ $X2=2.895 $Y2=0.152
r119 68 87 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.895 $Y=0.305
+ $X2=2.895 $Y2=0.152
r120 68 70 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.895 $Y=0.305
+ $X2=2.895 $Y2=0.825
r121 61 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.152
+ $X2=1.145 $Y2=0.152
r122 60 87 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.152
+ $X2=2.895 $Y2=0.152
r123 56 86 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.145 $Y=0.305
+ $X2=1.145 $Y2=0.152
r124 56 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.145 $Y=0.305
+ $X2=1.145 $Y2=0.825
r125 51 86 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.152
+ $X2=1.145 $Y2=0.152
r126 49 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.42 $Y=0.19
+ $X2=4.42 $Y2=0.19
r127 49 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.02 $Y=0.19
+ $X2=1.02 $Y2=0.19
r128 49 80 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.365 $Y2=0.305
r129 49 72 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0.152
+ $X2=4.28 $Y2=0.152
r130 49 72 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.28 $Y2=0.152
r131 49 73 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=3.06 $Y=0.152 $X2=2.98
+ $Y2=0.152
r132 49 60 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.81 $Y2=0.152
r133 49 61 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.23 $Y2=0.152
r134 49 51 1.6 $w=3.05e-07 $l=4e-08 $layer=LI1_cond $X=1.02 $Y=0.152 $X2=1.06
+ $Y2=0.152
r135 3 82 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.225
+ $Y=0.575 $X2=4.365 $Y2=0.825
r136 2 70 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.575 $X2=2.895 $Y2=0.825
r137 1 58 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.575 $X2=1.145 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%VDD 1 2 3 37 41 47 51 59 63 71 80 86 88
+ 90 94
r61 92 94 0.00232861 $w=3.05e-07 $l=5e-09 $layer=MET1_cond $X=4.42 $Y=6.507
+ $X2=4.425 $Y2=6.507
r62 90 92 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=3.735 $Y=6.507
+ $X2=4.42 $Y2=6.507
r63 88 90 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=3.055 $Y=6.507
+ $X2=3.735 $Y2=6.507
r64 86 88 0.314362 $w=3.05e-07 $l=6.75e-07 $layer=MET1_cond $X=2.38 $Y=6.507
+ $X2=3.055 $Y2=6.507
r65 83 86 0.633381 $w=3.05e-07 $l=1.36e-06 $layer=MET1_cond $X=1.02 $Y=6.507
+ $X2=2.38 $Y2=6.507
r66 80 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.42 $Y=6.47
+ $X2=4.42 $Y2=6.47
r67 71 74 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.365 $Y=3.455
+ $X2=4.365 $Y2=5.835
r68 69 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.365 $Y=6.355
+ $X2=4.365 $Y2=6.507
r69 69 74 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.365 $Y=6.355
+ $X2=4.365 $Y2=5.835
r70 66 68 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=6.507
+ $X2=3.74 $Y2=6.507
r71 64 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=6.507
+ $X2=2.895 $Y2=6.507
r72 64 66 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=2.98 $Y=6.507 $X2=3.06
+ $Y2=6.507
r73 63 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=6.507
+ $X2=4.365 $Y2=6.507
r74 63 68 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=4.28 $Y=6.507
+ $X2=3.74 $Y2=6.507
r75 59 62 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.895 $Y=3.455
+ $X2=2.895 $Y2=5.835
r76 57 78 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.895 $Y=6.355
+ $X2=2.895 $Y2=6.507
r77 57 62 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.895 $Y=6.355
+ $X2=2.895 $Y2=5.835
r78 54 56 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=6.507
+ $X2=2.38 $Y2=6.507
r79 52 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=6.507
+ $X2=1.145 $Y2=6.507
r80 52 54 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.23 $Y=6.507 $X2=1.7
+ $Y2=6.507
r81 51 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=6.507
+ $X2=2.895 $Y2=6.507
r82 51 56 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.81 $Y=6.507
+ $X2=2.38 $Y2=6.507
r83 47 50 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.145 $Y=3.795
+ $X2=1.145 $Y2=5.835
r84 45 77 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.145 $Y=6.355
+ $X2=1.145 $Y2=6.507
r85 45 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.145 $Y=6.355
+ $X2=1.145 $Y2=5.835
r86 43 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.02 $Y=6.47
+ $X2=1.02 $Y2=6.47
r87 41 77 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=6.507
+ $X2=1.145 $Y2=6.507
r88 41 43 1.6 $w=3.05e-07 $l=4e-08 $layer=LI1_cond $X=1.06 $Y=6.507 $X2=1.02
+ $Y2=6.507
r89 37 80 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r90 37 68 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r91 37 66 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r92 37 56 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r93 37 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r94 37 43 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r95 3 74 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.225
+ $Y=3.085 $X2=4.365 $Y2=5.835
r96 3 71 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.225
+ $Y=3.085 $X2=4.365 $Y2=3.455
r97 2 62 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.755
+ $Y=3.085 $X2=2.895 $Y2=5.835
r98 2 59 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.755
+ $Y=3.085 $X2=2.895 $Y2=3.455
r99 1 50 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.005
+ $Y=3.085 $X2=1.145 $Y2=5.835
r100 1 47 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=1.005 $Y=3.085 $X2=1.145 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%A_161_337# 1 3 13 16 18 19 21 22 23 24
+ 25 27 28 30 31 32 35 39
r82 39 41 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=2.02 $Y=3.455
+ $X2=2.02 $Y2=5.835
r83 37 39 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=2.02 $Y=3.27
+ $X2=2.02 $Y2=3.455
r84 33 35 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=2.02 $Y=1.345
+ $X2=2.02 $Y2=0.825
r85 31 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.85 $Y=1.43
+ $X2=2.02 $Y2=1.345
r86 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.85 $Y=1.43
+ $X2=1.57 $Y2=1.43
r87 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=1.515
+ $X2=1.57 $Y2=1.43
r88 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.485 $Y=1.515
+ $X2=1.485 $Y2=1.765
r89 27 37 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.85 $Y=3.185
+ $X2=2.02 $Y2=3.27
r90 27 28 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.85 $Y=3.185
+ $X2=1.025 $Y2=3.185
r91 26 44 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.025 $Y=1.85
+ $X2=0.94 $Y2=1.81
r92 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.4 $Y=1.85
+ $X2=1.485 $Y2=1.765
r93 25 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.4 $Y=1.85
+ $X2=1.025 $Y2=1.85
r94 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.94 $Y=3.1
+ $X2=1.025 $Y2=3.185
r95 23 44 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=1.935
+ $X2=0.94 $Y2=1.81
r96 23 24 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=0.94 $Y=1.935
+ $X2=0.94 $Y2=3.1
r97 21 22 56.3681 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=0.905 $Y=2.805
+ $X2=0.905 $Y2=2.975
r98 20 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.88 $Y=2.015
+ $X2=0.88 $Y2=2.805
r99 18 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.85 $X2=0.94 $Y2=1.85
r100 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.85
+ $X2=0.94 $Y2=2.015
r101 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.85
+ $X2=0.94 $Y2=1.685
r102 16 22 517.347 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=0.93 $Y=4.585
+ $X2=0.93 $Y2=2.975
r103 13 19 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.93 $Y=1.075
+ $X2=0.93 $Y2=1.685
r104 3 41 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.795
+ $Y=3.085 $X2=2.02 $Y2=5.835
r105 3 39 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.795
+ $Y=3.085 $X2=2.02 $Y2=3.455
r106 1 35 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.795
+ $Y=0.575 $X2=2.02 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%D 3 7 10 14 20
c51 7 0 1.64001e-19 $X=1.36 $Y=4.585
c52 3 0 1.3839e-19 $X=1.36 $Y=1.075
r53 20 23 0.00169837 $w=3.68e-07 $l=5e-09 $layer=MET1_cond $X=1.352 $Y=2.59
+ $X2=1.352 $Y2=2.595
r54 17 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.3 $Y=2.595 $X2=1.3
+ $Y2=2.595
r55 14 17 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.3 $Y=2.425 $X2=1.3
+ $Y2=2.595
r56 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.3
+ $Y=2.425 $X2=1.3 $Y2=2.425
r57 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=2.425
+ $X2=1.3 $Y2=2.59
r58 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=2.425
+ $X2=1.3 $Y2=2.26
r59 7 12 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=1.36 $Y=4.585
+ $X2=1.36 $Y2=2.59
r60 3 11 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.36 $Y=1.075
+ $X2=1.36 $Y2=2.26
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%CK 3 7 8 10 13 15 18 22 23 25 26 30 31
+ 33 37 44 46 47 49
c123 44 0 9.95038e-20 $X=1.86 $Y=2.765
c124 31 0 1.3839e-19 $X=1.945 $Y=1.85
c125 30 0 1.64001e-19 $X=1.86 $Y=2.68
c126 25 0 1.9983e-19 $X=3.137 $Y=2.78
c127 18 0 1.47633e-20 $X=1.78 $Y=2.765
r128 47 49 0.0928211 $w=2.16e-07 $l=1.50997e-07 $layer=MET1_cond $X=2.41 $Y=1.85
+ $X2=2.26 $Y2=1.852
r129 46 53 0.101772 $w=2.27e-07 $l=1.71493e-07 $layer=MET1_cond $X=3.075 $Y=1.85
+ $X2=3.245 $Y2=1.847
r130 46 47 0.640317 $w=1.7e-07 $l=6.65e-07 $layer=MET1_cond $X=3.075 $Y=1.85
+ $X2=2.41 $Y2=1.85
r131 42 44 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.78 $Y=2.765
+ $X2=1.86 $Y2=2.765
r132 37 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.245 $Y=1.85
+ $X2=3.245 $Y2=1.85
r133 33 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.26 $Y=1.85
+ $X2=2.26 $Y2=1.85
r134 31 33 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.945 $Y=1.85
+ $X2=2.26 $Y2=1.85
r135 30 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=2.68
+ $X2=1.86 $Y2=2.765
r136 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.86 $Y=1.935
+ $X2=1.945 $Y2=1.85
r137 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.86 $Y=1.935
+ $X2=1.86 $Y2=2.68
r138 28 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.85 $X2=3.245 $Y2=1.85
r139 25 26 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=3.137 $Y=2.78
+ $X2=3.137 $Y2=2.93
r140 22 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.85 $X2=2.26 $Y2=1.85
r141 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.85
+ $X2=2.26 $Y2=1.685
r142 18 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=2.765 $X2=1.78 $Y2=2.765
r143 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=2.765
+ $X2=1.78 $Y2=2.93
r144 15 28 38.6212 $w=3.33e-07 $l=1.89222e-07 $layer=POLY_cond $X=3.165 $Y=2.015
+ $X2=3.217 $Y2=1.85
r145 15 25 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=3.165 $Y=2.015
+ $X2=3.165 $Y2=2.78
r146 13 26 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=3.11 $Y=4.585
+ $X2=3.11 $Y2=2.93
r147 8 28 41.516 $w=3.33e-07 $l=2.32422e-07 $layer=POLY_cond $X=3.11 $Y=1.665
+ $X2=3.217 $Y2=1.85
r148 8 10 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=1.075
r149 7 23 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.32 $Y=1.075
+ $X2=2.32 $Y2=1.685
r150 3 20 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.72 $Y=4.585
+ $X2=1.72 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%A_329_89# 1 3 11 13 14 19 22 23 26 33
+ 37 44 47 51 53 54 59
c125 54 0 1.47633e-20 $X=2.405 $Y=2.59
c126 22 0 1.2087e-19 $X=2.26 $Y=2.765
c127 13 0 9.95038e-20 $X=2.125 $Y=2.3
r128 54 56 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.405 $Y=2.59
+ $X2=2.26 $Y2=2.59
r129 53 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.18 $Y=2.59
+ $X2=3.325 $Y2=2.59
r130 53 54 0.746234 $w=1.7e-07 $l=7.75e-07 $layer=MET1_cond $X=3.18 $Y=2.59
+ $X2=2.405 $Y2=2.59
r131 49 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.325 $Y=2.27
+ $X2=3.595 $Y2=2.27
r132 45 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.325 $Y=1.42
+ $X2=3.595 $Y2=1.42
r133 44 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=2.185
+ $X2=3.595 $Y2=2.27
r134 43 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=1.505
+ $X2=3.595 $Y2=1.42
r135 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.595 $Y=1.505
+ $X2=3.595 $Y2=2.185
r136 39 41 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.325 $Y=3.455
+ $X2=3.325 $Y2=5.835
r137 37 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.325 $Y=2.59
+ $X2=3.325 $Y2=2.59
r138 37 39 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.325 $Y=2.59
+ $X2=3.325 $Y2=3.455
r139 35 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.355
+ $X2=3.325 $Y2=2.27
r140 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.325 $Y=2.355
+ $X2=3.325 $Y2=2.59
r141 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.335
+ $X2=3.325 $Y2=1.42
r142 31 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.325 $Y=1.335
+ $X2=3.325 $Y2=0.825
r143 26 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.26 $Y=2.59
+ $X2=2.26 $Y2=2.59
r144 26 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.26 $Y=2.59
+ $X2=2.26 $Y2=2.765
r145 22 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=2.765 $X2=2.26 $Y2=2.765
r146 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=2.765
+ $X2=2.26 $Y2=2.93
r147 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=2.765
+ $X2=2.26 $Y2=2.6
r148 19 24 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=2.32 $Y=4.585
+ $X2=2.32 $Y2=2.93
r149 15 23 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.2 $Y=2.375
+ $X2=2.2 $Y2=2.6
r150 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=2.3
+ $X2=2.2 $Y2=2.375
r151 13 14 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.125 $Y=2.3
+ $X2=1.795 $Y2=2.3
r152 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.72 $Y=2.225
+ $X2=1.795 $Y2=2.3
r153 9 11 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=1.72 $Y=2.225
+ $X2=1.72 $Y2=1.075
r154 3 41 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.185
+ $Y=3.085 $X2=3.325 $Y2=5.835
r155 3 39 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.185
+ $Y=3.085 $X2=3.325 $Y2=3.455
r156 1 33 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.185
+ $Y=0.575 $X2=3.325 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%A_118_115# 1 3 11 15 23 26 28 32 33 35
+ 36 37 38 42 45 49 54 59 65 68 73 74 78 81 83
c163 81 0 1.2087e-19 $X=2.595 $Y=2.22
c164 59 0 1.9983e-19 $X=4.035 $Y=2.22
c165 37 0 8.77106e-20 $X=4.125 $Y=2.855
c166 32 0 2.20611e-19 $X=4.035 $Y=2.22
r167 80 81 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.74 $Y=2.22
+ $X2=2.595 $Y2=2.22
r168 78 81 2.2896 $w=1.4e-07 $l=1.85e-06 $layer=MET1_cond $X=0.745 $Y=2.2
+ $X2=2.595 $Y2=2.2
r169 76 78 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.6 $Y=2.22
+ $X2=0.745 $Y2=2.22
r170 74 80 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=2.89 $Y=2.22
+ $X2=2.74 $Y2=2.22
r171 73 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.89 $Y=2.22
+ $X2=4.035 $Y2=2.22
r172 73 74 1.23762 $w=1.4e-07 $l=1e-06 $layer=MET1_cond $X=3.89 $Y=2.22 $X2=2.89
+ $Y2=2.22
r173 68 70 8.33135 $w=2.83e-07 $l=1.6e-07 $layer=LI1_cond $X=0.657 $Y=3.795
+ $X2=0.657 $Y2=3.955
r174 68 69 12.1728 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.657 $Y=3.795
+ $X2=0.657 $Y2=3.54
r175 63 65 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.6 $Y=1.395
+ $X2=0.715 $Y2=1.395
r176 59 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.035 $Y=2.22
+ $X2=4.035 $Y2=2.22
r177 54 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.74 $Y=2.22
+ $X2=2.74 $Y2=2.22
r178 49 51 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=5.835
r179 49 70 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.715 $Y=4.135
+ $X2=0.715 $Y2=3.955
r180 43 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=1.31
+ $X2=0.715 $Y2=1.395
r181 43 45 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.715 $Y=1.31
+ $X2=0.715 $Y2=0.825
r182 42 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.6 $Y=2.22 $X2=0.6
+ $Y2=2.22
r183 42 69 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.6 $Y=2.22
+ $X2=0.6 $Y2=3.54
r184 39 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=1.48 $X2=0.6
+ $Y2=1.395
r185 39 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.6 $Y=1.48 $X2=0.6
+ $Y2=2.22
r186 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=2.855
+ $X2=4.125 $Y2=3.005
r187 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.125 $Y=1.65
+ $X2=4.125 $Y2=1.8
r188 34 37 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.1 $Y=2.385 $X2=4.1
+ $Y2=2.855
r189 33 36 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.1 $Y=2.055
+ $X2=4.1 $Y2=1.8
r190 32 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=2.22 $X2=4.035 $Y2=2.22
r191 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.037 $Y=2.22
+ $X2=4.037 $Y2=2.385
r192 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.037 $Y=2.22
+ $X2=4.037 $Y2=2.055
r193 28 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=2.22 $X2=2.74 $Y2=2.22
r194 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=2.22
+ $X2=2.74 $Y2=2.385
r195 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=2.22
+ $X2=2.74 $Y2=2.055
r196 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=4.15 $Y=4.585
+ $X2=4.15 $Y2=3.005
r197 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.15 $Y=1.075
+ $X2=4.15 $Y2=1.65
r198 15 30 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=2.68 $Y=4.585
+ $X2=2.68 $Y2=2.385
r199 11 29 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.68 $Y=1.075
+ $X2=2.68 $Y2=2.055
r200 3 51 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.59
+ $Y=3.085 $X2=0.715 $Y2=5.835
r201 3 49 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.59
+ $Y=3.085 $X2=0.715 $Y2=4.135
r202 3 68 600 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=3.085 $X2=0.715 $Y2=3.795
r203 1 45 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.575 $X2=0.715 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%QN 1 3 11 15 18 23 27 33 34 35 36 40 44
c78 44 0 8.77106e-20 $X=3.94 $Y=2.96
c79 35 0 1.02575e-19 $X=4.435 $Y=2.765
c80 33 0 1.18035e-19 $X=4.435 $Y=1.85
c81 18 0 1.97615e-19 $X=4.52 $Y=2.22
r82 42 44 0.00296209 $w=2.11e-07 $l=5e-09 $layer=MET1_cond $X=3.935 $Y=2.96
+ $X2=3.94 $Y2=2.96
r83 38 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.52 $Y=2.68
+ $X2=4.52 $Y2=2.22
r84 37 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.52 $Y=1.935
+ $X2=4.52 $Y2=2.22
r85 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=2.765
+ $X2=4.52 $Y2=2.68
r86 35 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=2.765
+ $X2=4.02 $Y2=2.765
r87 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=1.85
+ $X2=4.52 $Y2=1.935
r88 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.435 $Y=1.85
+ $X2=4.02 $Y2=1.85
r89 29 31 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.935 $Y=3.455
+ $X2=3.935 $Y2=5.835
r90 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=2.96
+ $X2=3.935 $Y2=2.96
r91 27 29 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.935 $Y=2.96
+ $X2=3.935 $Y2=3.455
r92 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=2.85
+ $X2=4.02 $Y2=2.765
r93 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.935 $Y=2.85
+ $X2=3.935 $Y2=2.96
r94 21 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.935 $Y=1.765
+ $X2=4.02 $Y2=1.85
r95 21 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.935 $Y=1.765
+ $X2=3.935 $Y2=0.825
r96 18 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=2.22 $X2=4.52 $Y2=2.22
r97 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.22
+ $X2=4.52 $Y2=2.385
r98 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.22
+ $X2=4.52 $Y2=2.055
r99 15 20 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=4.58 $Y=4.585
+ $X2=4.58 $Y2=2.385
r100 11 19 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.58 $Y=1.075
+ $X2=4.58 $Y2=2.055
r101 3 31 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=3.81
+ $Y=3.085 $X2=3.935 $Y2=5.835
r102 3 29 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=3.81
+ $Y=3.085 $X2=3.935 $Y2=3.455
r103 1 23 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=3.81
+ $Y=0.575 $X2=3.935 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_HS__NDLAT_1%Q 1 3 11 15 17 24 25 28
r19 24 25 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=4.86 $Y=1.595
+ $X2=4.86 $Y2=3.16
r20 23 24 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.827 $Y=1.425
+ $X2=4.827 $Y2=1.595
r21 17 19 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.795 $Y=3.455
+ $X2=4.795 $Y2=5.835
r22 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.795 $Y=3.33
+ $X2=4.795 $Y2=3.33
r23 15 25 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.827 $Y=3.33
+ $X2=4.827 $Y2=3.16
r24 15 17 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.795 $Y=3.33
+ $X2=4.795 $Y2=3.455
r25 11 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.795 $Y=0.825
+ $X2=4.795 $Y2=1.425
r26 3 19 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.655
+ $Y=3.085 $X2=4.795 $Y2=5.835
r27 3 17 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.655
+ $Y=3.085 $X2=4.795 $Y2=3.455
r28 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.655
+ $Y=0.575 $X2=4.795 $Y2=0.825
.ends

