* File: sky130_osu_sc_12T_ms__dffr_l.spice
* Created: Fri Nov 12 15:22:47 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ms__dffr_l.pex.spice"
.subckt sky130_osu_sc_12T_ms__dffr_l  GND VDD RN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* RN	RN
* VDD	VDD
* GND	GND
MM1021 N_A_110_115#_M1021_d N_RN_M1021_g N_GND_M1021_s N_GND_M1021_b NSHORT
+ L=0.15 W=0.52 AD=0.1378 AS=0.1378 PD=1.57 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1018 N_A_217_605#_M1018_d N_A_110_115#_M1018_g N_GND_M1018_s N_GND_M1021_b
+ NSHORT L=0.15 W=0.36 AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75000.6 A=0.054 P=1.02 MULT=1
MM1005 N_GND_M1005_d N_A_342_442#_M1005_g N_A_217_605#_M1018_d N_GND_M1021_b
+ NSHORT L=0.15 W=0.36 AD=0.0954 AS=0.0504 PD=1.25 PS=0.64 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.6 SB=75000.2 A=0.054 P=1.02 MULT=1
MM1007 A_576_115# N_D_M1007_g N_GND_M1007_s N_GND_M1021_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75003.7 A=0.078 P=1.34 MULT=1
MM1031 N_A_342_442#_M1031_d N_A_618_89#_M1031_g A_576_115# N_GND_M1021_b NSHORT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75000.5 SB=75003.3 A=0.078 P=1.34 MULT=1
MM1026 A_768_115# N_CK_M1026_g N_A_342_442#_M1031_d N_GND_M1021_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.1 SB=75002.7 A=0.078 P=1.34 MULT=1
MM1027 N_GND_M1027_d N_A_217_605#_M1027_g A_768_115# N_GND_M1021_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.5 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1025 A_926_115# N_A_217_605#_M1025_g N_GND_M1027_d N_GND_M1021_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667
+ SA=75001.9 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1019 N_A_998_115#_M1019_d N_CK_M1019_g A_926_115# N_GND_M1021_b NSHORT L=0.15
+ W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75002.3 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1020 A_1118_115# N_A_618_89#_M1020_g N_A_998_115#_M1019_d N_GND_M1021_b NSHORT
+ L=0.15 W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1
+ R=3.46667 SA=75002.9 SB=75001 A=0.078 P=1.34 MULT=1
MM1023 N_GND_M1023_d N_A_1160_89#_M1023_g A_1118_115# N_GND_M1021_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1
+ R=3.46667 SA=75003.3 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1010 N_A_618_89#_M1010_d N_CK_M1010_g N_GND_M1023_d N_GND_M1021_b NSHORT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75003.7 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1012 N_A_1160_89#_M1012_d N_A_998_115#_M1012_g N_GND_M1012_s N_GND_M1021_b
+ NSHORT L=0.15 W=0.36 AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75000.6 A=0.054 P=1.02 MULT=1
MM1013 N_GND_M1013_d N_A_110_115#_M1013_g N_A_1160_89#_M1012_d N_GND_M1021_b
+ NSHORT L=0.15 W=0.36 AD=0.0954 AS=0.0504 PD=1.25 PS=0.64 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.6 SB=75000.2 A=0.054 P=1.02 MULT=1
MM1016 N_GND_M1016_d N_A_1160_89#_M1016_g N_QN_M1016_s N_GND_M1021_b NSHORT
+ L=0.15 W=0.36 AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75000.6 A=0.054 P=1.02 MULT=1
MM1008 N_Q_M1008_d N_QN_M1008_g N_GND_M1016_d N_GND_M1021_b NSHORT L=0.15 W=0.36
+ AD=0.0954 AS=0.0504 PD=1.25 PS=0.64 NRD=0 NRS=0 M=1 R=2.4 SA=75000.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1004 N_A_110_115#_M1004_d N_RN_M1004_g N_VDD_M1004_s N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1015 A_300_605# N_A_110_115#_M1015_g N_A_217_605#_M1015_s N_VDD_M1004_b PSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_VDD_M1002_d N_A_342_442#_M1002_g A_300_605# N_VDD_M1004_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1028 A_576_521# N_D_M1028_g N_VDD_M1028_s N_VDD_M1004_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1024 N_A_342_442#_M1024_d N_CK_M1024_g A_576_521# N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1017 A_768_521# N_A_618_89#_M1017_g N_A_342_442#_M1024_d N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1022 N_VDD_M1022_d N_A_217_605#_M1022_g A_768_521# N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1014 A_926_521# N_A_217_605#_M1014_g N_VDD_M1022_d N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_998_115#_M1003_d N_A_618_89#_M1003_g A_926_521# N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 A_1118_521# N_CK_M1000_g N_A_998_115#_M1003_d N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1009 N_VDD_M1009_d N_A_1160_89#_M1009_g A_1118_521# N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_A_618_89#_M1029_d N_CK_M1029_g N_VDD_M1009_d N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 A_1466_605# N_A_998_115#_M1006_g N_A_1160_89#_M1006_s N_VDD_M1004_b
+ PSHORT L=0.15 W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_VDD_M1030_d N_A_110_115#_M1030_g A_1466_605# N_VDD_M1004_b PSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VDD_M1011_d N_A_1160_89#_M1011_g N_QN_M1011_s N_VDD_M1004_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_Q_M1001_d N_QN_M1001_g N_VDD_M1011_d N_VDD_M1004_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX32_noxref N_GND_M1021_b N_VDD_M1004_b NWDIODE A=19.8481 P=23.39
pX33_noxref noxref_24 RN RN PROBETYPE=1
pX34_noxref noxref_25 D D PROBETYPE=1
pX35_noxref noxref_26 CK CK PROBETYPE=1
pX36_noxref noxref_27 QN QN PROBETYPE=1
pX37_noxref noxref_28 Q Q PROBETYPE=1
c_1769 A_926_521# 0 1.57671e-19 $X=4.63 $Y=2.605
*
.include "sky130_osu_sc_12T_ms__dffr_l.pxi.spice"
*
.ends
*
*
