* File: sky130_osu_sc_12T_hs__nor2_1.pxi.spice
* Created: Fri Nov 12 15:12:01 2021
* 
x_PM_SKY130_OSU_SC_12T_HS__NOR2_1%GND N_GND_M1002_s N_GND_M1001_d N_GND_M1002_b
+ N_GND_c_2_p N_GND_c_3_p N_GND_c_14_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_12T_HS__NOR2_1%GND
x_PM_SKY130_OSU_SC_12T_HS__NOR2_1%VDD N_VDD_M1003_d N_VDD_M1000_b N_VDD_c_29_p
+ N_VDD_c_35_p VDD N_VDD_c_30_p PM_SKY130_OSU_SC_12T_HS__NOR2_1%VDD
x_PM_SKY130_OSU_SC_12T_HS__NOR2_1%B N_B_M1002_g N_B_M1000_g N_B_c_51_n
+ N_B_c_53_n N_B_c_55_n B PM_SKY130_OSU_SC_12T_HS__NOR2_1%B
x_PM_SKY130_OSU_SC_12T_HS__NOR2_1%A N_A_M1003_g N_A_M1001_g N_A_c_99_n
+ N_A_c_100_n A PM_SKY130_OSU_SC_12T_HS__NOR2_1%A
x_PM_SKY130_OSU_SC_12T_HS__NOR2_1%Y N_Y_M1002_d N_Y_M1000_s N_Y_c_131_n
+ N_Y_c_132_n N_Y_c_135_n N_Y_c_136_n Y N_Y_c_138_n
+ PM_SKY130_OSU_SC_12T_HS__NOR2_1%Y
cc_1 N_GND_M1002_b N_B_M1002_g 0.0373962f $X=-0.045 $Y=0 $X2=0.475 $Y2=0.85
cc_2 N_GND_c_2_p N_B_M1002_g 0.00502587f $X=0.26 $Y=0.755 $X2=0.475 $Y2=0.85
cc_3 N_GND_c_3_p N_B_M1002_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=0.85
cc_4 N_GND_c_4_p N_B_M1002_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.475 $Y2=0.85
cc_5 N_GND_M1002_b N_B_M1000_g 0.0432223f $X=-0.045 $Y=0 $X2=0.475 $Y2=3.235
cc_6 N_GND_M1002_b N_B_c_51_n 0.0362021f $X=-0.045 $Y=0 $X2=0.415 $Y2=1.61
cc_7 N_GND_c_2_p N_B_c_51_n 0.00122211f $X=0.26 $Y=0.755 $X2=0.415 $Y2=1.61
cc_8 N_GND_M1002_b N_B_c_53_n 0.0115466f $X=-0.045 $Y=0 $X2=0.565 $Y2=1.61
cc_9 N_GND_c_2_p N_B_c_53_n 0.00289632f $X=0.26 $Y=0.755 $X2=0.565 $Y2=1.61
cc_10 N_GND_M1002_b N_B_c_55_n 0.0148611f $X=-0.045 $Y=0 $X2=0.65 $Y2=2.48
cc_11 N_GND_M1002_b B 5.75357e-19 $X=-0.045 $Y=0 $X2=0.65 $Y2=2.48
cc_12 N_GND_M1002_b N_A_M1001_g 0.0918519f $X=-0.045 $Y=0 $X2=0.905 $Y2=0.85
cc_13 N_GND_c_3_p N_A_M1001_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=0.85
cc_14 N_GND_c_14_p N_A_M1001_g 0.00502587f $X=1.12 $Y=0.755 $X2=0.905 $Y2=0.85
cc_15 N_GND_c_4_p N_A_M1001_g 0.00468827f $X=1.02 $Y=0.19 $X2=0.905 $Y2=0.85
cc_16 N_GND_M1002_b N_A_c_99_n 0.0416705f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.275
cc_17 N_GND_M1002_b N_A_c_100_n 0.00382838f $X=-0.045 $Y=0 $X2=0.99 $Y2=2.275
cc_18 N_GND_M1002_b N_Y_c_131_n 0.0154673f $X=-0.045 $Y=0 $X2=0.26 $Y2=2.11
cc_19 N_GND_M1002_b N_Y_c_132_n 0.00154299f $X=-0.045 $Y=0 $X2=0.69 $Y2=0.755
cc_20 N_GND_c_3_p N_Y_c_132_n 0.00740081f $X=1.035 $Y=0.152 $X2=0.69 $Y2=0.755
cc_21 N_GND_c_4_p N_Y_c_132_n 0.0047139f $X=1.02 $Y=0.19 $X2=0.69 $Y2=0.755
cc_22 N_GND_M1002_b N_Y_c_135_n 0.00182421f $X=-0.045 $Y=0 $X2=0.605 $Y2=2.11
cc_23 N_GND_M1002_b N_Y_c_136_n 0.0197856f $X=-0.045 $Y=0 $X2=0.405 $Y2=2.11
cc_24 N_GND_M1002_b Y 0.0193014f $X=-0.045 $Y=0 $X2=0.685 $Y2=1.485
cc_25 N_GND_c_2_p N_Y_c_138_n 0.00125659f $X=0.26 $Y=0.755 $X2=0.69 $Y2=1
cc_26 N_GND_c_3_p N_Y_c_138_n 0.00245319f $X=1.035 $Y=0.152 $X2=0.69 $Y2=1
cc_27 N_GND_c_14_p N_Y_c_138_n 0.00125659f $X=1.12 $Y=0.755 $X2=0.69 $Y2=1
cc_28 N_VDD_M1000_b N_B_M1000_g 0.0246289f $X=-0.045 $Y=2.425 $X2=0.475
+ $Y2=3.235
cc_29 N_VDD_c_29_p N_B_M1000_g 0.00606474f $X=0.965 $Y=4.287 $X2=0.475 $Y2=3.235
cc_30 N_VDD_c_30_p N_B_M1000_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.475 $Y2=3.235
cc_31 N_VDD_M1000_b N_B_c_55_n 0.00408216f $X=-0.045 $Y=2.425 $X2=0.65 $Y2=2.48
cc_32 N_VDD_M1000_b B 0.00838127f $X=-0.045 $Y=2.425 $X2=0.65 $Y2=2.48
cc_33 N_VDD_M1000_b N_A_M1003_g 0.0199366f $X=-0.045 $Y=2.425 $X2=0.835
+ $Y2=3.235
cc_34 N_VDD_c_29_p N_A_M1003_g 0.00606474f $X=0.965 $Y=4.287 $X2=0.835 $Y2=3.235
cc_35 N_VDD_c_35_p N_A_M1003_g 0.00636672f $X=1.05 $Y=3.635 $X2=0.835 $Y2=3.235
cc_36 N_VDD_c_30_p N_A_M1003_g 0.00468827f $X=1.02 $Y=4.25 $X2=0.835 $Y2=3.235
cc_37 N_VDD_M1000_b N_A_c_99_n 0.00807651f $X=-0.045 $Y=2.425 $X2=0.99 $Y2=2.275
cc_38 N_VDD_M1003_d N_A_c_100_n 0.00953431f $X=0.91 $Y=2.605 $X2=0.99 $Y2=2.275
cc_39 N_VDD_M1000_b N_A_c_100_n 0.00566834f $X=-0.045 $Y=2.425 $X2=0.99
+ $Y2=2.275
cc_40 N_VDD_c_35_p N_A_c_100_n 0.00252874f $X=1.05 $Y=3.635 $X2=0.99 $Y2=2.275
cc_41 N_VDD_M1003_d A 0.0150141f $X=0.91 $Y=2.605 $X2=0.99 $Y2=2.85
cc_42 N_VDD_c_35_p A 0.00522047f $X=1.05 $Y=3.635 $X2=0.99 $Y2=2.85
cc_43 N_VDD_M1000_b N_Y_c_131_n 0.00981538f $X=-0.045 $Y=2.425 $X2=0.26 $Y2=2.11
cc_44 N_VDD_c_29_p N_Y_c_131_n 0.00736239f $X=0.965 $Y=4.287 $X2=0.26 $Y2=2.11
cc_45 N_VDD_c_30_p N_Y_c_131_n 0.00476261f $X=1.02 $Y=4.25 $X2=0.26 $Y2=2.11
cc_46 B N_A_M1003_g 0.00231474f $X=0.65 $Y=2.48 $X2=0.835 $Y2=3.235
cc_47 N_B_M1002_g N_A_M1001_g 0.0548658f $X=0.475 $Y=0.85 $X2=0.905 $Y2=0.85
cc_48 N_B_c_53_n N_A_M1001_g 0.00368334f $X=0.565 $Y=1.61 $X2=0.905 $Y2=0.85
cc_49 N_B_c_55_n N_A_M1001_g 0.00805543f $X=0.65 $Y=2.48 $X2=0.905 $Y2=0.85
cc_50 N_B_M1000_g N_A_c_99_n 0.115892f $X=0.475 $Y=3.235 $X2=0.99 $Y2=2.275
cc_51 N_B_c_55_n N_A_c_99_n 0.00287728f $X=0.65 $Y=2.48 $X2=0.99 $Y2=2.275
cc_52 B N_A_c_99_n 0.00187972f $X=0.65 $Y=2.48 $X2=0.99 $Y2=2.275
cc_53 N_B_M1000_g N_A_c_100_n 0.00136939f $X=0.475 $Y=3.235 $X2=0.99 $Y2=2.275
cc_54 N_B_c_55_n N_A_c_100_n 0.029766f $X=0.65 $Y=2.48 $X2=0.99 $Y2=2.275
cc_55 B N_A_c_100_n 0.00643447f $X=0.65 $Y=2.48 $X2=0.99 $Y2=2.275
cc_56 N_B_M1000_g A 0.00297933f $X=0.475 $Y=3.235 $X2=0.99 $Y2=2.85
cc_57 B A 0.0050603f $X=0.65 $Y=2.48 $X2=0.99 $Y2=2.85
cc_58 N_B_M1000_g N_Y_c_131_n 0.0158498f $X=0.475 $Y=3.235 $X2=0.26 $Y2=2.11
cc_59 N_B_c_51_n N_Y_c_131_n 0.00138434f $X=0.415 $Y=1.61 $X2=0.26 $Y2=2.11
cc_60 N_B_c_53_n N_Y_c_131_n 0.00308264f $X=0.565 $Y=1.61 $X2=0.26 $Y2=2.11
cc_61 N_B_c_55_n N_Y_c_131_n 0.0294278f $X=0.65 $Y=2.48 $X2=0.26 $Y2=2.11
cc_62 B N_Y_c_131_n 0.00774605f $X=0.65 $Y=2.48 $X2=0.26 $Y2=2.11
cc_63 N_B_M1002_g N_Y_c_132_n 0.00182852f $X=0.475 $Y=0.85 $X2=0.69 $Y2=0.755
cc_64 N_B_c_53_n N_Y_c_132_n 0.00335445f $X=0.565 $Y=1.61 $X2=0.69 $Y2=0.755
cc_65 N_B_M1000_g N_Y_c_135_n 0.00382028f $X=0.475 $Y=3.235 $X2=0.605 $Y2=2.11
cc_66 N_B_c_53_n N_Y_c_135_n 0.00523952f $X=0.565 $Y=1.61 $X2=0.605 $Y2=2.11
cc_67 N_B_c_55_n N_Y_c_135_n 0.0116239f $X=0.65 $Y=2.48 $X2=0.605 $Y2=2.11
cc_68 B N_Y_c_135_n 0.0327205f $X=0.65 $Y=2.48 $X2=0.605 $Y2=2.11
cc_69 N_B_M1000_g N_Y_c_136_n 0.00327819f $X=0.475 $Y=3.235 $X2=0.405 $Y2=2.11
cc_70 N_B_c_51_n N_Y_c_136_n 0.00301446f $X=0.415 $Y=1.61 $X2=0.405 $Y2=2.11
cc_71 N_B_c_53_n N_Y_c_136_n 0.00469337f $X=0.565 $Y=1.61 $X2=0.405 $Y2=2.11
cc_72 N_B_c_55_n N_Y_c_136_n 0.00157282f $X=0.65 $Y=2.48 $X2=0.405 $Y2=2.11
cc_73 B N_Y_c_136_n 9.25684e-19 $X=0.65 $Y=2.48 $X2=0.405 $Y2=2.11
cc_74 N_B_M1002_g Y 0.00594872f $X=0.475 $Y=0.85 $X2=0.685 $Y2=1.485
cc_75 N_B_c_53_n Y 0.0124433f $X=0.565 $Y=1.61 $X2=0.685 $Y2=1.485
cc_76 N_B_c_55_n Y 0.0178687f $X=0.65 $Y=2.48 $X2=0.685 $Y2=1.485
cc_77 N_B_M1002_g N_Y_c_138_n 0.00837334f $X=0.475 $Y=0.85 $X2=0.69 $Y2=1
cc_78 N_B_c_53_n N_Y_c_138_n 0.00244196f $X=0.565 $Y=1.61 $X2=0.69 $Y2=1
cc_79 N_A_c_100_n N_Y_c_131_n 0.00350166f $X=0.99 $Y=2.275 $X2=0.26 $Y2=2.11
cc_80 A N_Y_c_131_n 0.00623956f $X=0.99 $Y=2.85 $X2=0.26 $Y2=2.11
cc_81 N_A_M1001_g N_Y_c_132_n 0.00182852f $X=0.905 $Y=0.85 $X2=0.69 $Y2=0.755
cc_82 N_A_c_99_n N_Y_c_135_n 0.00155621f $X=0.99 $Y=2.275 $X2=0.605 $Y2=2.11
cc_83 N_A_c_100_n N_Y_c_135_n 0.00255034f $X=0.99 $Y=2.275 $X2=0.605 $Y2=2.11
cc_84 N_A_M1001_g Y 0.0148599f $X=0.905 $Y=0.85 $X2=0.685 $Y2=1.485
cc_85 N_A_M1001_g N_Y_c_138_n 0.00852585f $X=0.905 $Y=0.85 $X2=0.69 $Y2=1
cc_86 A A_110_521# 0.00289505f $X=0.99 $Y=2.85 $X2=0.55 $Y2=2.605
