* File: sky130_osu_sc_12T_ls__dffs_1.spice
* Created: Fri Nov 12 15:36:23 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ls__dffs_1.pex.spice"
.subckt sky130_osu_sc_12T_ls__dffs_1  GND VDD SN D CK QN Q
* 
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* VDD	VDD
* GND	GND
MM1012 A_110_115# N_SN_M1012_g N_A_27_115#_M1012_s N_GND_M1012_b NSHORT L=0.15
+ W=0.36 AD=0.0378 AS=0.0954 PD=0.57 PS=1.25 NRD=16.656 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75000.6 A=0.054 P=1.02 MULT=1
MM1000 N_GND_M1000_d N_A_152_89#_M1000_g A_110_115# N_GND_M1012_b NSHORT L=0.15
+ W=0.36 AD=0.0954 AS=0.0378 PD=1.25 PS=0.57 NRD=0 NRS=16.656 M=1 R=2.4
+ SA=75000.6 SB=75000.2 A=0.054 P=1.02 MULT=1
MM1001 A_386_115# N_D_M1001_g N_GND_M1001_s N_GND_M1012_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75003.7 A=0.078 P=1.34 MULT=1
MM1023 N_A_152_89#_M1023_d N_A_428_89#_M1023_g A_386_115# N_GND_M1012_b NSHORT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75000.5 SB=75003.3 A=0.078 P=1.34 MULT=1
MM1018 A_578_115# N_CK_M1018_g N_A_152_89#_M1023_d N_GND_M1012_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.1 SB=75002.7 A=0.078 P=1.34 MULT=1
MM1021 N_GND_M1021_d N_A_27_115#_M1021_g A_578_115# N_GND_M1012_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.5 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1013 A_736_115# N_A_27_115#_M1013_g N_GND_M1021_d N_GND_M1012_b NSHORT L=0.15
+ W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667
+ SA=75001.9 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1010 N_A_808_115#_M1010_d N_CK_M1010_g A_736_115# N_GND_M1012_b NSHORT L=0.15
+ W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75002.3 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1002 A_928_115# N_A_428_89#_M1002_g N_A_808_115#_M1010_d N_GND_M1012_b NSHORT
+ L=0.15 W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1
+ R=3.46667 SA=75002.9 SB=75001 A=0.078 P=1.34 MULT=1
MM1006 N_GND_M1006_d N_A_970_89#_M1006_g A_928_115# N_GND_M1012_b NSHORT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75003.3 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1003 N_A_428_89#_M1003_d N_CK_M1003_g N_GND_M1006_d N_GND_M1012_b NSHORT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75003.7 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1004 A_1276_115# N_A_808_115#_M1004_g N_A_970_89#_M1004_s N_GND_M1012_b NSHORT
+ L=0.15 W=0.36 AD=0.0378 AS=0.0954 PD=0.57 PS=1.25 NRD=16.656 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75000.6 A=0.054 P=1.02 MULT=1
MM1025 N_GND_M1025_d N_SN_M1025_g A_1276_115# N_GND_M1012_b NSHORT L=0.15 W=0.36
+ AD=0.0954 AS=0.0378 PD=1.25 PS=0.57 NRD=0 NRS=16.656 M=1 R=2.4 SA=75000.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1008 N_GND_M1008_d N_A_970_89#_M1008_g N_QN_M1008_s N_GND_M1012_b NSHORT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1027 N_Q_M1027_d N_QN_M1027_g N_GND_M1008_d N_GND_M1012_b NSHORT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1009 N_A_27_115#_M1009_d N_SN_M1009_g N_VDD_M1009_s N_VDD_M1009_b PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_VDD_M1020_d N_A_152_89#_M1020_g N_A_27_115#_M1009_d N_VDD_M1009_b
+ PHIGHVT L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 A_386_521# N_D_M1007_g N_VDD_M1007_s N_VDD_M1009_b PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1011 N_A_152_89#_M1011_d N_CK_M1011_g A_386_521# N_VDD_M1009_b PHIGHVT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1015 A_578_521# N_A_428_89#_M1015_g N_A_152_89#_M1011_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1014 N_VDD_M1014_d N_A_27_115#_M1014_g A_578_521# N_VDD_M1009_b PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1005 A_736_521# N_A_27_115#_M1005_g N_VDD_M1014_d N_VDD_M1009_b PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1022 N_A_808_115#_M1022_d N_A_428_89#_M1022_g A_736_521# N_VDD_M1009_b PHIGHVT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1028 A_928_521# N_CK_M1028_g N_A_808_115#_M1022_d N_VDD_M1009_b PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1026 N_VDD_M1026_d N_A_970_89#_M1026_g A_928_521# N_VDD_M1009_b PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_A_428_89#_M1017_d N_CK_M1017_g N_VDD_M1026_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1024 N_A_970_89#_M1024_d N_A_808_115#_M1024_g N_VDD_M1024_s N_VDD_M1009_b
+ PHIGHVT L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_VDD_M1016_d N_SN_M1016_g N_A_970_89#_M1024_d N_VDD_M1009_b PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1029 N_VDD_M1029_d N_A_970_89#_M1029_g N_QN_M1029_s N_VDD_M1009_b PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_Q_M1019_d N_QN_M1019_g N_VDD_M1029_d N_VDD_M1009_b PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX30_noxref N_GND_M1012_b N_VDD_M1009_b NWDIODE A=18.0409 P=21.64
pX31_noxref noxref_23 SN SN PROBETYPE=1
pX32_noxref noxref_24 D D PROBETYPE=1
pX33_noxref noxref_25 CK CK PROBETYPE=1
pX34_noxref noxref_26 QN QN PROBETYPE=1
pX35_noxref noxref_27 Q Q PROBETYPE=1
c_1609 A_736_521# 0 1.57671e-19 $X=3.68 $Y=2.605
*
.include "sky130_osu_sc_12T_ls__dffs_1.pxi.spice"
*
.ends
*
*
