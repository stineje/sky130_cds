* File: sky130_osu_sc_18T_ms__or2_8.pxi.spice
* Created: Thu Oct 29 17:31:22 2020
* 
x_PM_SKY130_OSU_SC_18T_MS__OR2_8%GND N_GND_M1004_s N_GND_M1000_d N_GND_M1005_s
+ N_GND_M1010_s N_GND_M1014_s N_GND_M1018_s N_GND_M1004_b N_GND_c_2_p
+ N_GND_c_3_p N_GND_c_11_p N_GND_c_18_p N_GND_c_24_p N_GND_c_32_p N_GND_c_38_p
+ N_GND_c_45_p N_GND_c_52_p N_GND_c_64_p N_GND_c_59_p GND N_GND_c_4_p
+ PM_SKY130_OSU_SC_18T_MS__OR2_8%GND
x_PM_SKY130_OSU_SC_18T_MS__OR2_8%VDD N_VDD_M1001_d N_VDD_M1007_s N_VDD_M1011_s
+ N_VDD_M1015_s N_VDD_M1019_s N_VDD_M1006_b N_VDD_c_142_p N_VDD_c_150_p
+ N_VDD_c_156_p N_VDD_c_162_p N_VDD_c_167_p N_VDD_c_173_p N_VDD_c_178_p
+ N_VDD_c_188_p N_VDD_c_137_p N_VDD_c_184_p VDD N_VDD_c_138_p
+ PM_SKY130_OSU_SC_18T_MS__OR2_8%VDD
x_PM_SKY130_OSU_SC_18T_MS__OR2_8%B N_B_M1004_g N_B_M1006_g B N_B_c_223_n
+ N_B_c_224_n PM_SKY130_OSU_SC_18T_MS__OR2_8%B
x_PM_SKY130_OSU_SC_18T_MS__OR2_8%A N_A_M1000_g N_A_M1001_g A N_A_c_250_n
+ N_A_c_251_n PM_SKY130_OSU_SC_18T_MS__OR2_8%A
x_PM_SKY130_OSU_SC_18T_MS__OR2_8%A_27_617# N_A_27_617#_M1004_d
+ N_A_27_617#_M1006_s N_A_27_617#_M1002_g N_A_27_617#_c_359_n
+ N_A_27_617#_M1003_g N_A_27_617#_c_293_n N_A_27_617#_c_294_n
+ N_A_27_617#_M1005_g N_A_27_617#_c_364_n N_A_27_617#_M1007_g
+ N_A_27_617#_c_299_n N_A_27_617#_c_301_n N_A_27_617#_c_302_n
+ N_A_27_617#_M1008_g N_A_27_617#_c_371_n N_A_27_617#_M1009_g
+ N_A_27_617#_c_307_n N_A_27_617#_c_308_n N_A_27_617#_M1010_g
+ N_A_27_617#_c_376_n N_A_27_617#_M1011_g N_A_27_617#_c_313_n
+ N_A_27_617#_c_315_n N_A_27_617#_M1012_g N_A_27_617#_c_320_n
+ N_A_27_617#_c_382_n N_A_27_617#_M1013_g N_A_27_617#_c_321_n
+ N_A_27_617#_c_322_n N_A_27_617#_M1014_g N_A_27_617#_c_387_n
+ N_A_27_617#_M1015_g N_A_27_617#_c_327_n N_A_27_617#_c_329_n
+ N_A_27_617#_M1016_g N_A_27_617#_c_393_n N_A_27_617#_M1017_g
+ N_A_27_617#_c_334_n N_A_27_617#_c_335_n N_A_27_617#_M1018_g
+ N_A_27_617#_c_398_n N_A_27_617#_M1019_g N_A_27_617#_c_340_n
+ N_A_27_617#_c_341_n N_A_27_617#_c_342_n N_A_27_617#_c_343_n
+ N_A_27_617#_c_344_n N_A_27_617#_c_345_n N_A_27_617#_c_346_n
+ N_A_27_617#_c_347_n N_A_27_617#_c_348_n N_A_27_617#_c_349_n
+ N_A_27_617#_c_350_n N_A_27_617#_c_351_n N_A_27_617#_c_409_n
+ N_A_27_617#_c_413_n N_A_27_617#_c_415_n N_A_27_617#_c_352_n
+ N_A_27_617#_c_353_n N_A_27_617#_c_356_n N_A_27_617#_c_358_n
+ PM_SKY130_OSU_SC_18T_MS__OR2_8%A_27_617#
x_PM_SKY130_OSU_SC_18T_MS__OR2_8%Y N_Y_M1002_d N_Y_M1008_d N_Y_M1012_d
+ N_Y_M1016_d N_Y_M1003_d N_Y_M1009_d N_Y_M1013_d N_Y_M1017_d N_Y_c_535_n
+ N_Y_c_538_n Y N_Y_c_540_n N_Y_c_542_n N_Y_c_543_n N_Y_c_544_n N_Y_c_546_n
+ N_Y_c_549_n N_Y_c_550_n N_Y_c_551_n N_Y_c_554_n N_Y_c_555_n N_Y_c_556_n
+ N_Y_c_557_n N_Y_c_560_n N_Y_c_561_n N_Y_c_562_n N_Y_c_563_n N_Y_c_564_n
+ N_Y_c_566_n N_Y_c_567_n N_Y_c_571_n N_Y_c_576_n N_Y_c_581_n
+ PM_SKY130_OSU_SC_18T_MS__OR2_8%Y
cc_1 N_GND_M1004_b N_B_M1004_g 0.083817f $X=-0.045 $Y=0 $X2=0.475 $Y2=1.075
cc_2 N_GND_c_2_p N_B_M1004_g 0.00713292f $X=0.26 $Y=0.825 $X2=0.475 $Y2=1.075
cc_3 N_GND_c_3_p N_B_M1004_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.475 $Y2=1.075
cc_4 N_GND_c_4_p N_B_M1004_g 0.00468827f $X=4.42 $Y=0.17 $X2=0.475 $Y2=1.075
cc_5 N_GND_M1004_b N_B_M1006_g 0.0039012f $X=-0.045 $Y=0 $X2=0.475 $Y2=4.585
cc_6 N_GND_M1004_b B 0.00409308f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.96
cc_7 N_GND_M1004_b N_B_c_223_n 0.00781915f $X=-0.045 $Y=0 $X2=0.27 $Y2=2.675
cc_8 N_GND_M1004_b N_B_c_224_n 0.0541719f $X=-0.045 $Y=0 $X2=0.475 $Y2=2.675
cc_9 N_GND_M1004_b N_A_M1000_g 0.0440597f $X=-0.045 $Y=0 $X2=0.905 $Y2=1.075
cc_10 N_GND_c_3_p N_A_M1000_g 0.00606474f $X=1.035 $Y=0.152 $X2=0.905 $Y2=1.075
cc_11 N_GND_c_11_p N_A_M1000_g 0.00354579f $X=1.12 $Y=0.825 $X2=0.905 $Y2=1.075
cc_12 N_GND_c_4_p N_A_M1000_g 0.00468827f $X=4.42 $Y=0.17 $X2=0.905 $Y2=1.075
cc_13 N_GND_M1004_b N_A_M1001_g 0.0174023f $X=-0.045 $Y=0 $X2=0.905 $Y2=4.585
cc_14 N_GND_M1004_b N_A_c_250_n 0.0034276f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.385
cc_15 N_GND_M1004_b N_A_c_251_n 0.0291701f $X=-0.045 $Y=0 $X2=0.95 $Y2=2.385
cc_16 N_GND_M1004_b N_A_27_617#_M1002_g 0.0207501f $X=-0.045 $Y=0 $X2=1.335
+ $Y2=1.075
cc_17 N_GND_c_11_p N_A_27_617#_M1002_g 0.00354579f $X=1.12 $Y=0.825 $X2=1.335
+ $Y2=1.075
cc_18 N_GND_c_18_p N_A_27_617#_M1002_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.335
+ $Y2=1.075
cc_19 N_GND_c_4_p N_A_27_617#_M1002_g 0.00468827f $X=4.42 $Y=0.17 $X2=1.335
+ $Y2=1.075
cc_20 N_GND_M1004_b N_A_27_617#_c_293_n 0.0466273f $X=-0.045 $Y=0 $X2=1.37
+ $Y2=2.81
cc_21 N_GND_M1004_b N_A_27_617#_c_294_n 0.00727817f $X=-0.045 $Y=0 $X2=1.69
+ $Y2=2.885
cc_22 N_GND_M1004_b N_A_27_617#_M1005_g 0.020212f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=1.075
cc_23 N_GND_c_18_p N_A_27_617#_M1005_g 0.00606474f $X=1.895 $Y=0.152 $X2=1.765
+ $Y2=1.075
cc_24 N_GND_c_24_p N_A_27_617#_M1005_g 0.00356864f $X=1.98 $Y=0.825 $X2=1.765
+ $Y2=1.075
cc_25 N_GND_c_4_p N_A_27_617#_M1005_g 0.00468827f $X=4.42 $Y=0.17 $X2=1.765
+ $Y2=1.075
cc_26 N_GND_M1004_b N_A_27_617#_c_299_n 0.0181078f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=1.845
cc_27 N_GND_c_24_p N_A_27_617#_c_299_n 0.00256938f $X=1.98 $Y=0.825 $X2=2.12
+ $Y2=1.845
cc_28 N_GND_M1004_b N_A_27_617#_c_301_n 0.0447518f $X=-0.045 $Y=0 $X2=1.84
+ $Y2=1.845
cc_29 N_GND_M1004_b N_A_27_617#_c_302_n 0.013058f $X=-0.045 $Y=0 $X2=2.12
+ $Y2=2.885
cc_30 N_GND_M1004_b N_A_27_617#_M1008_g 0.020212f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.075
cc_31 N_GND_c_24_p N_A_27_617#_M1008_g 0.00356864f $X=1.98 $Y=0.825 $X2=2.195
+ $Y2=1.075
cc_32 N_GND_c_32_p N_A_27_617#_M1008_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.195
+ $Y2=1.075
cc_33 N_GND_c_4_p N_A_27_617#_M1008_g 0.00468827f $X=4.42 $Y=0.17 $X2=2.195
+ $Y2=1.075
cc_34 N_GND_M1004_b N_A_27_617#_c_307_n 0.0180386f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=1.845
cc_35 N_GND_M1004_b N_A_27_617#_c_308_n 0.0118833f $X=-0.045 $Y=0 $X2=2.55
+ $Y2=2.885
cc_36 N_GND_M1004_b N_A_27_617#_M1010_g 0.020212f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.075
cc_37 N_GND_c_32_p N_A_27_617#_M1010_g 0.00606474f $X=2.755 $Y=0.152 $X2=2.625
+ $Y2=1.075
cc_38 N_GND_c_38_p N_A_27_617#_M1010_g 0.00356864f $X=2.84 $Y=0.825 $X2=2.625
+ $Y2=1.075
cc_39 N_GND_c_4_p N_A_27_617#_M1010_g 0.00468827f $X=4.42 $Y=0.17 $X2=2.625
+ $Y2=1.075
cc_40 N_GND_M1004_b N_A_27_617#_c_313_n 0.0181078f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=1.845
cc_41 N_GND_c_38_p N_A_27_617#_c_313_n 0.00256938f $X=2.84 $Y=0.825 $X2=2.98
+ $Y2=1.845
cc_42 N_GND_M1004_b N_A_27_617#_c_315_n 0.00959015f $X=-0.045 $Y=0 $X2=2.98
+ $Y2=2.885
cc_43 N_GND_M1004_b N_A_27_617#_M1012_g 0.020212f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.075
cc_44 N_GND_c_38_p N_A_27_617#_M1012_g 0.00356864f $X=2.84 $Y=0.825 $X2=3.055
+ $Y2=1.075
cc_45 N_GND_c_45_p N_A_27_617#_M1012_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.055
+ $Y2=1.075
cc_46 N_GND_c_4_p N_A_27_617#_M1012_g 0.00468827f $X=4.42 $Y=0.17 $X2=3.055
+ $Y2=1.075
cc_47 N_GND_M1004_b N_A_27_617#_c_320_n 0.0620214f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.81
cc_48 N_GND_M1004_b N_A_27_617#_c_321_n 0.0180386f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=1.845
cc_49 N_GND_M1004_b N_A_27_617#_c_322_n 0.0118833f $X=-0.045 $Y=0 $X2=3.41
+ $Y2=2.885
cc_50 N_GND_M1004_b N_A_27_617#_M1014_g 0.020212f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.075
cc_51 N_GND_c_45_p N_A_27_617#_M1014_g 0.00606474f $X=3.615 $Y=0.152 $X2=3.485
+ $Y2=1.075
cc_52 N_GND_c_52_p N_A_27_617#_M1014_g 0.00356864f $X=3.7 $Y=0.825 $X2=3.485
+ $Y2=1.075
cc_53 N_GND_c_4_p N_A_27_617#_M1014_g 0.00468827f $X=4.42 $Y=0.17 $X2=3.485
+ $Y2=1.075
cc_54 N_GND_M1004_b N_A_27_617#_c_327_n 0.0181078f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=1.845
cc_55 N_GND_c_52_p N_A_27_617#_c_327_n 0.00256938f $X=3.7 $Y=0.825 $X2=3.84
+ $Y2=1.845
cc_56 N_GND_M1004_b N_A_27_617#_c_329_n 0.013058f $X=-0.045 $Y=0 $X2=3.84
+ $Y2=2.885
cc_57 N_GND_M1004_b N_A_27_617#_M1016_g 0.020212f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=1.075
cc_58 N_GND_c_52_p N_A_27_617#_M1016_g 0.00356864f $X=3.7 $Y=0.825 $X2=3.915
+ $Y2=1.075
cc_59 N_GND_c_59_p N_A_27_617#_M1016_g 0.00606474f $X=4.475 $Y=0.152 $X2=3.915
+ $Y2=1.075
cc_60 N_GND_c_4_p N_A_27_617#_M1016_g 0.00468827f $X=4.42 $Y=0.17 $X2=3.915
+ $Y2=1.075
cc_61 N_GND_M1004_b N_A_27_617#_c_334_n 0.0369419f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=1.845
cc_62 N_GND_M1004_b N_A_27_617#_c_335_n 0.0268552f $X=-0.045 $Y=0 $X2=4.27
+ $Y2=2.885
cc_63 N_GND_M1004_b N_A_27_617#_M1018_g 0.0264941f $X=-0.045 $Y=0 $X2=4.345
+ $Y2=1.075
cc_64 N_GND_c_64_p N_A_27_617#_M1018_g 0.00713292f $X=4.56 $Y=0.825 $X2=4.345
+ $Y2=1.075
cc_65 N_GND_c_59_p N_A_27_617#_M1018_g 0.00606474f $X=4.475 $Y=0.152 $X2=4.345
+ $Y2=1.075
cc_66 N_GND_c_4_p N_A_27_617#_M1018_g 0.00468827f $X=4.42 $Y=0.17 $X2=4.345
+ $Y2=1.075
cc_67 N_GND_M1004_b N_A_27_617#_c_340_n 0.00568338f $X=-0.045 $Y=0 $X2=1.352
+ $Y2=2.885
cc_68 N_GND_M1004_b N_A_27_617#_c_341_n 0.00735657f $X=-0.045 $Y=0 $X2=1.765
+ $Y2=2.885
cc_69 N_GND_M1004_b N_A_27_617#_c_342_n 0.00873941f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=1.845
cc_70 N_GND_M1004_b N_A_27_617#_c_343_n 0.00735657f $X=-0.045 $Y=0 $X2=2.195
+ $Y2=2.885
cc_71 N_GND_M1004_b N_A_27_617#_c_344_n 0.00873941f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=1.845
cc_72 N_GND_M1004_b N_A_27_617#_c_345_n 0.00735657f $X=-0.045 $Y=0 $X2=2.625
+ $Y2=2.885
cc_73 N_GND_M1004_b N_A_27_617#_c_346_n 0.0023879f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=1.845
cc_74 N_GND_M1004_b N_A_27_617#_c_347_n 0.00151234f $X=-0.045 $Y=0 $X2=3.055
+ $Y2=2.885
cc_75 N_GND_M1004_b N_A_27_617#_c_348_n 0.00873941f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=1.845
cc_76 N_GND_M1004_b N_A_27_617#_c_349_n 0.00735657f $X=-0.045 $Y=0 $X2=3.485
+ $Y2=2.885
cc_77 N_GND_M1004_b N_A_27_617#_c_350_n 0.00873941f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=1.845
cc_78 N_GND_M1004_b N_A_27_617#_c_351_n 0.00735657f $X=-0.045 $Y=0 $X2=3.915
+ $Y2=2.885
cc_79 N_GND_M1004_b N_A_27_617#_c_352_n 0.00591391f $X=-0.045 $Y=0 $X2=0.61
+ $Y2=3.545
cc_80 N_GND_M1004_b N_A_27_617#_c_353_n 0.00710171f $X=-0.045 $Y=0 $X2=0.69
+ $Y2=0.825
cc_81 N_GND_c_3_p N_A_27_617#_c_353_n 0.0075556f $X=1.035 $Y=0.152 $X2=0.69
+ $Y2=0.825
cc_82 N_GND_c_4_p N_A_27_617#_c_353_n 0.00475776f $X=4.42 $Y=0.17 $X2=0.69
+ $Y2=0.825
cc_83 N_GND_M1004_b N_A_27_617#_c_356_n 0.0190355f $X=-0.045 $Y=0 $X2=1.43
+ $Y2=1.935
cc_84 N_GND_c_11_p N_A_27_617#_c_356_n 0.00702738f $X=1.12 $Y=0.825 $X2=1.43
+ $Y2=1.935
cc_85 N_GND_M1004_b N_A_27_617#_c_358_n 0.00549821f $X=-0.045 $Y=0 $X2=0.65
+ $Y2=1.935
cc_86 N_GND_M1004_b N_Y_c_535_n 0.00248416f $X=-0.045 $Y=0 $X2=1.55 $Y2=1.595
cc_87 N_GND_c_11_p N_Y_c_535_n 0.00134236f $X=1.12 $Y=0.825 $X2=1.55 $Y2=1.595
cc_88 N_GND_c_24_p N_Y_c_535_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=1.595
cc_89 N_GND_M1004_b N_Y_c_538_n 0.00509006f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.475
cc_90 N_GND_M1004_b Y 0.0305055f $X=-0.045 $Y=0 $X2=1.555 $Y2=2.22
cc_91 N_GND_M1005_s N_Y_c_540_n 0.0127884f $X=1.84 $Y=0.575 $X2=2.265 $Y2=1.48
cc_92 N_GND_c_24_p N_Y_c_540_n 0.0142303f $X=1.98 $Y=0.825 $X2=2.265 $Y2=1.48
cc_93 N_GND_M1004_b N_Y_c_542_n 0.018807f $X=-0.045 $Y=0 $X2=2.265 $Y2=2.59
cc_94 N_GND_M1004_b N_Y_c_543_n 0.0367149f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.475
cc_95 N_GND_M1010_s N_Y_c_544_n 0.0127884f $X=2.7 $Y=0.575 $X2=3.125 $Y2=1.48
cc_96 N_GND_c_38_p N_Y_c_544_n 0.0142303f $X=2.84 $Y=0.825 $X2=3.125 $Y2=1.48
cc_97 N_GND_M1004_b N_Y_c_546_n 0.00409378f $X=-0.045 $Y=0 $X2=2.555 $Y2=1.48
cc_98 N_GND_c_24_p N_Y_c_546_n 7.53951e-19 $X=1.98 $Y=0.825 $X2=2.555 $Y2=1.48
cc_99 N_GND_c_38_p N_Y_c_546_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=2.555 $Y2=1.48
cc_100 N_GND_M1004_b N_Y_c_549_n 0.0144211f $X=-0.045 $Y=0 $X2=3.125 $Y2=2.59
cc_101 N_GND_M1004_b N_Y_c_550_n 0.0069606f $X=-0.045 $Y=0 $X2=2.555 $Y2=2.59
cc_102 N_GND_M1004_b N_Y_c_551_n 0.00409378f $X=-0.045 $Y=0 $X2=3.27 $Y2=1.595
cc_103 N_GND_c_38_p N_Y_c_551_n 7.53951e-19 $X=2.84 $Y=0.825 $X2=3.27 $Y2=1.595
cc_104 N_GND_c_52_p N_Y_c_551_n 8.22956e-19 $X=3.7 $Y=0.825 $X2=3.27 $Y2=1.595
cc_105 N_GND_M1004_b N_Y_c_554_n 0.0358528f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.475
cc_106 N_GND_M1004_b N_Y_c_555_n 0.018807f $X=-0.045 $Y=0 $X2=3.985 $Y2=2.59
cc_107 N_GND_M1004_b N_Y_c_556_n 0.00584404f $X=-0.045 $Y=0 $X2=3.415 $Y2=2.59
cc_108 N_GND_M1004_b N_Y_c_557_n 0.00409378f $X=-0.045 $Y=0 $X2=4.13 $Y2=1.595
cc_109 N_GND_c_52_p N_Y_c_557_n 7.53951e-19 $X=3.7 $Y=0.825 $X2=4.13 $Y2=1.595
cc_110 N_GND_c_64_p N_Y_c_557_n 0.00134792f $X=4.56 $Y=0.825 $X2=4.13 $Y2=1.595
cc_111 N_GND_M1004_b N_Y_c_560_n 0.06145f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.475
cc_112 N_GND_M1004_b N_Y_c_561_n 0.0107267f $X=-0.045 $Y=0 $X2=1.55 $Y2=2.59
cc_113 N_GND_M1004_b N_Y_c_562_n 0.0149623f $X=-0.045 $Y=0 $X2=2.41 $Y2=2.59
cc_114 N_GND_M1004_b N_Y_c_563_n 0.0149086f $X=-0.045 $Y=0 $X2=3.27 $Y2=2.59
cc_115 N_GND_M1014_s N_Y_c_564_n 0.0129565f $X=3.56 $Y=0.575 $X2=4.13 $Y2=1.48
cc_116 N_GND_c_52_p N_Y_c_564_n 0.0140638f $X=3.7 $Y=0.825 $X2=4.13 $Y2=1.48
cc_117 N_GND_M1004_b N_Y_c_566_n 0.0152877f $X=-0.045 $Y=0 $X2=4.13 $Y2=2.59
cc_118 N_GND_M1004_b N_Y_c_567_n 0.00155118f $X=-0.045 $Y=0 $X2=1.55 $Y2=0.825
cc_119 N_GND_c_18_p N_Y_c_567_n 0.00737727f $X=1.895 $Y=0.152 $X2=1.55 $Y2=0.825
cc_120 N_GND_c_24_p N_Y_c_567_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=1.55 $Y2=0.825
cc_121 N_GND_c_4_p N_Y_c_567_n 0.00475776f $X=4.42 $Y=0.17 $X2=1.55 $Y2=0.825
cc_122 N_GND_M1004_b N_Y_c_571_n 0.00155118f $X=-0.045 $Y=0 $X2=2.41 $Y2=0.825
cc_123 N_GND_c_24_p N_Y_c_571_n 8.14297e-19 $X=1.98 $Y=0.825 $X2=2.41 $Y2=0.825
cc_124 N_GND_c_32_p N_Y_c_571_n 0.00734006f $X=2.755 $Y=0.152 $X2=2.41 $Y2=0.825
cc_125 N_GND_c_38_p N_Y_c_571_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=2.41 $Y2=0.825
cc_126 N_GND_c_4_p N_Y_c_571_n 0.00475776f $X=4.42 $Y=0.17 $X2=2.41 $Y2=0.825
cc_127 N_GND_M1004_b N_Y_c_576_n 0.00155118f $X=-0.045 $Y=0 $X2=3.27 $Y2=0.825
cc_128 N_GND_c_38_p N_Y_c_576_n 8.14297e-19 $X=2.84 $Y=0.825 $X2=3.27 $Y2=0.825
cc_129 N_GND_c_45_p N_Y_c_576_n 0.00745425f $X=3.615 $Y=0.152 $X2=3.27 $Y2=0.825
cc_130 N_GND_c_52_p N_Y_c_576_n 8.14297e-19 $X=3.7 $Y=0.825 $X2=3.27 $Y2=0.825
cc_131 N_GND_c_4_p N_Y_c_576_n 0.00475776f $X=4.42 $Y=0.17 $X2=3.27 $Y2=0.825
cc_132 N_GND_M1004_b N_Y_c_581_n 0.00155118f $X=-0.045 $Y=0 $X2=4.13 $Y2=0.825
cc_133 N_GND_c_52_p N_Y_c_581_n 8.14297e-19 $X=3.7 $Y=0.825 $X2=4.13 $Y2=0.825
cc_134 N_GND_c_59_p N_Y_c_581_n 0.0075556f $X=4.475 $Y=0.152 $X2=4.13 $Y2=0.825
cc_135 N_GND_c_4_p N_Y_c_581_n 0.00475776f $X=4.42 $Y=0.17 $X2=4.13 $Y2=0.825
cc_136 N_VDD_M1006_b N_B_M1006_g 0.0260091f $X=-0.045 $Y=2.905 $X2=0.475
+ $Y2=4.585
cc_137 N_VDD_c_137_p N_B_M1006_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.475
+ $Y2=4.585
cc_138 N_VDD_c_138_p N_B_M1006_g 0.00468827f $X=4.42 $Y=6.49 $X2=0.475 $Y2=4.585
cc_139 N_VDD_M1006_b B 0.0108395f $X=-0.045 $Y=2.905 $X2=0.27 $Y2=2.96
cc_140 N_VDD_M1006_b N_B_c_223_n 0.00375034f $X=-0.045 $Y=2.905 $X2=0.27
+ $Y2=2.675
cc_141 N_VDD_M1006_b N_A_M1001_g 0.0195137f $X=-0.045 $Y=2.905 $X2=0.905
+ $Y2=4.585
cc_142 N_VDD_c_142_p N_A_M1001_g 0.00354579f $X=1.12 $Y=4.135 $X2=0.905
+ $Y2=4.585
cc_143 N_VDD_c_137_p N_A_M1001_g 0.00606474f $X=1.035 $Y=6.507 $X2=0.905
+ $Y2=4.585
cc_144 N_VDD_c_138_p N_A_M1001_g 0.00468827f $X=4.42 $Y=6.49 $X2=0.905 $Y2=4.585
cc_145 N_VDD_M1001_d A 0.0077995f $X=0.98 $Y=3.085 $X2=0.95 $Y2=3.33
cc_146 N_VDD_c_142_p A 0.00247404f $X=1.12 $Y=4.135 $X2=0.95 $Y2=3.33
cc_147 N_VDD_M1006_b N_A_c_250_n 0.00153494f $X=-0.045 $Y=2.905 $X2=0.95
+ $Y2=2.385
cc_148 N_VDD_M1006_b N_A_27_617#_c_359_n 0.0170965f $X=-0.045 $Y=2.905 $X2=1.335
+ $Y2=2.96
cc_149 N_VDD_c_142_p N_A_27_617#_c_359_n 0.00354579f $X=1.12 $Y=4.135 $X2=1.335
+ $Y2=2.96
cc_150 N_VDD_c_150_p N_A_27_617#_c_359_n 0.00606474f $X=1.895 $Y=6.507 $X2=1.335
+ $Y2=2.96
cc_151 N_VDD_c_138_p N_A_27_617#_c_359_n 0.00468827f $X=4.42 $Y=6.49 $X2=1.335
+ $Y2=2.96
cc_152 N_VDD_M1006_b N_A_27_617#_c_294_n 0.00427883f $X=-0.045 $Y=2.905 $X2=1.69
+ $Y2=2.885
cc_153 N_VDD_M1006_b N_A_27_617#_c_364_n 0.017006f $X=-0.045 $Y=2.905 $X2=1.765
+ $Y2=2.96
cc_154 N_VDD_c_142_p N_A_27_617#_c_364_n 3.67508e-19 $X=1.12 $Y=4.135 $X2=1.765
+ $Y2=2.96
cc_155 N_VDD_c_150_p N_A_27_617#_c_364_n 0.00610567f $X=1.895 $Y=6.507 $X2=1.765
+ $Y2=2.96
cc_156 N_VDD_c_156_p N_A_27_617#_c_364_n 0.00373985f $X=1.98 $Y=3.455 $X2=1.765
+ $Y2=2.96
cc_157 N_VDD_c_138_p N_A_27_617#_c_364_n 0.00470215f $X=4.42 $Y=6.49 $X2=1.765
+ $Y2=2.96
cc_158 N_VDD_M1006_b N_A_27_617#_c_302_n 0.00396043f $X=-0.045 $Y=2.905 $X2=2.12
+ $Y2=2.885
cc_159 N_VDD_c_156_p N_A_27_617#_c_302_n 0.00379272f $X=1.98 $Y=3.455 $X2=2.12
+ $Y2=2.885
cc_160 N_VDD_M1006_b N_A_27_617#_c_371_n 0.0166898f $X=-0.045 $Y=2.905 $X2=2.195
+ $Y2=2.96
cc_161 N_VDD_c_156_p N_A_27_617#_c_371_n 0.00354579f $X=1.98 $Y=3.455 $X2=2.195
+ $Y2=2.96
cc_162 N_VDD_c_162_p N_A_27_617#_c_371_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.195
+ $Y2=2.96
cc_163 N_VDD_c_138_p N_A_27_617#_c_371_n 0.00468827f $X=4.42 $Y=6.49 $X2=2.195
+ $Y2=2.96
cc_164 N_VDD_M1006_b N_A_27_617#_c_308_n 0.00448664f $X=-0.045 $Y=2.905 $X2=2.55
+ $Y2=2.885
cc_165 N_VDD_M1006_b N_A_27_617#_c_376_n 0.0166898f $X=-0.045 $Y=2.905 $X2=2.625
+ $Y2=2.96
cc_166 N_VDD_c_162_p N_A_27_617#_c_376_n 0.00606474f $X=2.755 $Y=6.507 $X2=2.625
+ $Y2=2.96
cc_167 N_VDD_c_167_p N_A_27_617#_c_376_n 0.00354579f $X=2.84 $Y=3.455 $X2=2.625
+ $Y2=2.96
cc_168 N_VDD_c_138_p N_A_27_617#_c_376_n 0.00468827f $X=4.42 $Y=6.49 $X2=2.625
+ $Y2=2.96
cc_169 N_VDD_M1006_b N_A_27_617#_c_315_n 0.00396043f $X=-0.045 $Y=2.905 $X2=2.98
+ $Y2=2.885
cc_170 N_VDD_c_167_p N_A_27_617#_c_315_n 0.00379272f $X=2.84 $Y=3.455 $X2=2.98
+ $Y2=2.885
cc_171 N_VDD_M1006_b N_A_27_617#_c_382_n 0.0166898f $X=-0.045 $Y=2.905 $X2=3.055
+ $Y2=2.96
cc_172 N_VDD_c_167_p N_A_27_617#_c_382_n 0.00354579f $X=2.84 $Y=3.455 $X2=3.055
+ $Y2=2.96
cc_173 N_VDD_c_173_p N_A_27_617#_c_382_n 0.00606474f $X=3.615 $Y=6.507 $X2=3.055
+ $Y2=2.96
cc_174 N_VDD_c_138_p N_A_27_617#_c_382_n 0.00468827f $X=4.42 $Y=6.49 $X2=3.055
+ $Y2=2.96
cc_175 N_VDD_M1006_b N_A_27_617#_c_322_n 0.00448664f $X=-0.045 $Y=2.905 $X2=3.41
+ $Y2=2.885
cc_176 N_VDD_M1006_b N_A_27_617#_c_387_n 0.0166898f $X=-0.045 $Y=2.905 $X2=3.485
+ $Y2=2.96
cc_177 N_VDD_c_173_p N_A_27_617#_c_387_n 0.00606474f $X=3.615 $Y=6.507 $X2=3.485
+ $Y2=2.96
cc_178 N_VDD_c_178_p N_A_27_617#_c_387_n 0.00354579f $X=3.7 $Y=3.455 $X2=3.485
+ $Y2=2.96
cc_179 N_VDD_c_138_p N_A_27_617#_c_387_n 0.00468827f $X=4.42 $Y=6.49 $X2=3.485
+ $Y2=2.96
cc_180 N_VDD_M1006_b N_A_27_617#_c_329_n 0.00396043f $X=-0.045 $Y=2.905 $X2=3.84
+ $Y2=2.885
cc_181 N_VDD_c_178_p N_A_27_617#_c_329_n 0.00379272f $X=3.7 $Y=3.455 $X2=3.84
+ $Y2=2.885
cc_182 N_VDD_M1006_b N_A_27_617#_c_393_n 0.0166898f $X=-0.045 $Y=2.905 $X2=3.915
+ $Y2=2.96
cc_183 N_VDD_c_178_p N_A_27_617#_c_393_n 0.00354579f $X=3.7 $Y=3.455 $X2=3.915
+ $Y2=2.96
cc_184 N_VDD_c_184_p N_A_27_617#_c_393_n 0.00606474f $X=4.475 $Y=6.507 $X2=3.915
+ $Y2=2.96
cc_185 N_VDD_c_138_p N_A_27_617#_c_393_n 0.00468827f $X=4.42 $Y=6.49 $X2=3.915
+ $Y2=2.96
cc_186 N_VDD_M1006_b N_A_27_617#_c_335_n 0.00840215f $X=-0.045 $Y=2.905 $X2=4.27
+ $Y2=2.885
cc_187 N_VDD_M1006_b N_A_27_617#_c_398_n 0.0209036f $X=-0.045 $Y=2.905 $X2=4.345
+ $Y2=2.96
cc_188 N_VDD_c_188_p N_A_27_617#_c_398_n 0.00713292f $X=4.56 $Y=3.455 $X2=4.345
+ $Y2=2.96
cc_189 N_VDD_c_184_p N_A_27_617#_c_398_n 0.00606474f $X=4.475 $Y=6.507 $X2=4.345
+ $Y2=2.96
cc_190 N_VDD_c_138_p N_A_27_617#_c_398_n 0.00468827f $X=4.42 $Y=6.49 $X2=4.345
+ $Y2=2.96
cc_191 N_VDD_M1006_b N_A_27_617#_c_340_n 0.0021704f $X=-0.045 $Y=2.905 $X2=1.352
+ $Y2=2.885
cc_192 N_VDD_M1006_b N_A_27_617#_c_341_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=1.765 $Y2=2.885
cc_193 N_VDD_M1006_b N_A_27_617#_c_343_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.195 $Y2=2.885
cc_194 N_VDD_M1006_b N_A_27_617#_c_345_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=2.625 $Y2=2.885
cc_195 N_VDD_M1006_b N_A_27_617#_c_347_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=3.055 $Y2=2.885
cc_196 N_VDD_M1006_b N_A_27_617#_c_349_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=3.485 $Y2=2.885
cc_197 N_VDD_M1006_b N_A_27_617#_c_351_n 8.75564e-19 $X=-0.045 $Y=2.905
+ $X2=3.915 $Y2=2.885
cc_198 N_VDD_M1006_b N_A_27_617#_c_409_n 0.00156053f $X=-0.045 $Y=2.905 $X2=0.26
+ $Y2=3.795
cc_199 N_VDD_c_137_p N_A_27_617#_c_409_n 0.00736239f $X=1.035 $Y=6.507 $X2=0.26
+ $Y2=3.795
cc_200 N_VDD_c_138_p N_A_27_617#_c_409_n 0.00476261f $X=4.42 $Y=6.49 $X2=0.26
+ $Y2=3.795
cc_201 N_VDD_M1006_b N_A_27_617#_c_352_n 0.00106577f $X=-0.045 $Y=2.905 $X2=0.61
+ $Y2=3.545
cc_202 N_VDD_c_156_p N_Y_c_542_n 0.00634153f $X=1.98 $Y=3.455 $X2=2.265 $Y2=2.59
cc_203 N_VDD_c_167_p N_Y_c_549_n 0.00634153f $X=2.84 $Y=3.455 $X2=3.125 $Y2=2.59
cc_204 N_VDD_c_178_p N_Y_c_555_n 0.00634153f $X=3.7 $Y=3.455 $X2=3.985 $Y2=2.59
cc_205 N_VDD_M1006_b N_Y_c_561_n 0.00367096f $X=-0.045 $Y=2.905 $X2=1.55
+ $Y2=2.59
cc_206 N_VDD_c_150_p N_Y_c_561_n 0.00737727f $X=1.895 $Y=6.507 $X2=1.55 $Y2=2.59
cc_207 N_VDD_c_138_p N_Y_c_561_n 0.00475776f $X=4.42 $Y=6.49 $X2=1.55 $Y2=2.59
cc_208 N_VDD_M1006_b N_Y_c_562_n 0.00380347f $X=-0.045 $Y=2.905 $X2=2.41
+ $Y2=2.59
cc_209 N_VDD_c_162_p N_Y_c_562_n 0.00734006f $X=2.755 $Y=6.507 $X2=2.41 $Y2=2.59
cc_210 N_VDD_c_138_p N_Y_c_562_n 0.00475776f $X=4.42 $Y=6.49 $X2=2.41 $Y2=2.59
cc_211 N_VDD_M1006_b N_Y_c_563_n 0.00380347f $X=-0.045 $Y=2.905 $X2=3.27
+ $Y2=2.59
cc_212 N_VDD_c_173_p N_Y_c_563_n 0.00745425f $X=3.615 $Y=6.507 $X2=3.27 $Y2=2.59
cc_213 N_VDD_c_138_p N_Y_c_563_n 0.00475776f $X=4.42 $Y=6.49 $X2=3.27 $Y2=2.59
cc_214 N_VDD_M1006_b N_Y_c_566_n 0.00380347f $X=-0.045 $Y=2.905 $X2=4.13
+ $Y2=2.59
cc_215 N_VDD_c_184_p N_Y_c_566_n 0.0075556f $X=4.475 $Y=6.507 $X2=4.13 $Y2=2.59
cc_216 N_VDD_c_138_p N_Y_c_566_n 0.00475776f $X=4.42 $Y=6.49 $X2=4.13 $Y2=2.59
cc_217 N_B_M1004_g N_A_M1000_g 0.0402111f $X=0.475 $Y=1.075 $X2=0.905 $Y2=1.075
cc_218 N_B_c_224_n N_A_M1001_g 0.154838f $X=0.475 $Y=2.675 $X2=0.905 $Y2=4.585
cc_219 N_B_M1004_g N_A_c_250_n 0.00121111f $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.385
cc_220 N_B_M1004_g N_A_c_251_n 0.0148656f $X=0.475 $Y=1.075 $X2=0.95 $Y2=2.385
cc_221 N_B_M1006_g N_A_27_617#_c_413_n 0.0140282f $X=0.475 $Y=4.585 $X2=0.525
+ $Y2=3.63
cc_222 B N_A_27_617#_c_413_n 0.00520961f $X=0.27 $Y=2.96 $X2=0.525 $Y2=3.63
cc_223 B N_A_27_617#_c_415_n 0.00431991f $X=0.27 $Y=2.96 $X2=0.345 $Y2=3.63
cc_224 N_B_c_223_n N_A_27_617#_c_415_n 0.00369517f $X=0.27 $Y=2.675 $X2=0.345
+ $Y2=3.63
cc_225 N_B_M1004_g N_A_27_617#_c_352_n 0.0231435f $X=0.475 $Y=1.075 $X2=0.61
+ $Y2=3.545
cc_226 N_B_M1006_g N_A_27_617#_c_352_n 0.026563f $X=0.475 $Y=4.585 $X2=0.61
+ $Y2=3.545
cc_227 B N_A_27_617#_c_352_n 0.00758489f $X=0.27 $Y=2.96 $X2=0.61 $Y2=3.545
cc_228 N_B_c_223_n N_A_27_617#_c_352_n 0.0350086f $X=0.27 $Y=2.675 $X2=0.61
+ $Y2=3.545
cc_229 N_B_c_224_n N_A_27_617#_c_352_n 0.00764878f $X=0.475 $Y=2.675 $X2=0.61
+ $Y2=3.545
cc_230 N_B_M1004_g N_A_27_617#_c_353_n 0.00765999f $X=0.475 $Y=1.075 $X2=0.69
+ $Y2=0.825
cc_231 N_B_M1004_g N_A_27_617#_c_358_n 0.0113001f $X=0.475 $Y=1.075 $X2=0.65
+ $Y2=1.935
cc_232 N_A_M1000_g N_A_27_617#_M1002_g 0.0310007f $X=0.905 $Y=1.075 $X2=1.335
+ $Y2=1.075
cc_233 A N_A_27_617#_c_359_n 0.00374181f $X=0.95 $Y=3.33 $X2=1.335 $Y2=2.96
cc_234 N_A_M1001_g N_A_27_617#_c_293_n 0.00914307f $X=0.905 $Y=4.585 $X2=1.37
+ $Y2=2.81
cc_235 N_A_c_250_n N_A_27_617#_c_293_n 0.00375034f $X=0.95 $Y=2.385 $X2=1.37
+ $Y2=2.81
cc_236 N_A_c_251_n N_A_27_617#_c_293_n 0.0204279f $X=0.95 $Y=2.385 $X2=1.37
+ $Y2=2.81
cc_237 N_A_M1000_g N_A_27_617#_c_301_n 0.0119161f $X=0.905 $Y=1.075 $X2=1.84
+ $Y2=1.845
cc_238 N_A_M1001_g N_A_27_617#_c_340_n 0.0547156f $X=0.905 $Y=4.585 $X2=1.352
+ $Y2=2.885
cc_239 N_A_c_250_n N_A_27_617#_c_340_n 0.00358357f $X=0.95 $Y=2.385 $X2=1.352
+ $Y2=2.885
cc_240 N_A_M1001_g N_A_27_617#_c_413_n 0.00457566f $X=0.905 $Y=4.585 $X2=0.525
+ $Y2=3.63
cc_241 N_A_M1000_g N_A_27_617#_c_352_n 0.00429604f $X=0.905 $Y=1.075 $X2=0.61
+ $Y2=3.545
cc_242 N_A_M1001_g N_A_27_617#_c_352_n 0.00776428f $X=0.905 $Y=4.585 $X2=0.61
+ $Y2=3.545
cc_243 A N_A_27_617#_c_352_n 0.00866797f $X=0.95 $Y=3.33 $X2=0.61 $Y2=3.545
cc_244 N_A_c_250_n N_A_27_617#_c_352_n 0.0822139f $X=0.95 $Y=2.385 $X2=0.61
+ $Y2=3.545
cc_245 N_A_c_251_n N_A_27_617#_c_352_n 0.0021255f $X=0.95 $Y=2.385 $X2=0.61
+ $Y2=3.545
cc_246 N_A_M1000_g N_A_27_617#_c_353_n 0.00765999f $X=0.905 $Y=1.075 $X2=0.69
+ $Y2=0.825
cc_247 N_A_M1000_g N_A_27_617#_c_356_n 0.0163305f $X=0.905 $Y=1.075 $X2=1.43
+ $Y2=1.935
cc_248 N_A_c_250_n N_A_27_617#_c_356_n 0.0114342f $X=0.95 $Y=2.385 $X2=1.43
+ $Y2=1.935
cc_249 N_A_c_251_n N_A_27_617#_c_356_n 0.00276813f $X=0.95 $Y=2.385 $X2=1.43
+ $Y2=1.935
cc_250 A A_110_617# 0.0123256f $X=0.95 $Y=3.33 $X2=0.55 $Y2=3.085
cc_251 N_A_M1000_g N_Y_c_535_n 8.23842e-19 $X=0.905 $Y=1.075 $X2=1.55 $Y2=1.595
cc_252 N_A_c_250_n N_Y_c_538_n 0.0059581f $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.475
cc_253 N_A_c_251_n N_Y_c_538_n 3.73261e-19 $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.475
cc_254 N_A_M1000_g Y 6.73508e-19 $X=0.905 $Y=1.075 $X2=1.555 $Y2=2.22
cc_255 N_A_c_250_n Y 0.00825539f $X=0.95 $Y=2.385 $X2=1.555 $Y2=2.22
cc_256 A N_Y_c_561_n 0.00659455f $X=0.95 $Y=3.33 $X2=1.55 $Y2=2.59
cc_257 N_A_c_250_n N_Y_c_561_n 0.0206732f $X=0.95 $Y=2.385 $X2=1.55 $Y2=2.59
cc_258 N_A_27_617#_c_413_n A_110_617# 0.00613297f $X=0.525 $Y=3.63 $X2=0.55
+ $Y2=3.085
cc_259 N_A_27_617#_c_352_n A_110_617# 0.00377193f $X=0.61 $Y=3.545 $X2=0.55
+ $Y2=3.085
cc_260 N_A_27_617#_M1002_g N_Y_c_535_n 0.00542903f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_261 N_A_27_617#_M1005_g N_Y_c_535_n 0.00259902f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=1.595
cc_262 N_A_27_617#_c_356_n N_Y_c_535_n 0.00238892f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=1.595
cc_263 N_A_27_617#_c_293_n N_Y_c_538_n 0.00821104f $X=1.37 $Y=2.81 $X2=1.55
+ $Y2=2.475
cc_264 N_A_27_617#_c_294_n N_Y_c_538_n 0.00186325f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.475
cc_265 N_A_27_617#_c_301_n N_Y_c_538_n 0.00194187f $X=1.84 $Y=1.845 $X2=1.55
+ $Y2=2.475
cc_266 N_A_27_617#_c_356_n N_Y_c_538_n 0.00181779f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.475
cc_267 N_A_27_617#_M1002_g Y 0.00251111f $X=1.335 $Y=1.075 $X2=1.555 $Y2=2.22
cc_268 N_A_27_617#_c_293_n Y 0.00892438f $X=1.37 $Y=2.81 $X2=1.555 $Y2=2.22
cc_269 N_A_27_617#_M1005_g Y 0.00251111f $X=1.765 $Y=1.075 $X2=1.555 $Y2=2.22
cc_270 N_A_27_617#_c_301_n Y 0.0131034f $X=1.84 $Y=1.845 $X2=1.555 $Y2=2.22
cc_271 N_A_27_617#_c_356_n Y 0.0147088f $X=1.43 $Y=1.935 $X2=1.555 $Y2=2.22
cc_272 N_A_27_617#_M1005_g N_Y_c_540_n 0.0130095f $X=1.765 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_273 N_A_27_617#_c_299_n N_Y_c_540_n 0.00213861f $X=2.12 $Y=1.845 $X2=2.265
+ $Y2=1.48
cc_274 N_A_27_617#_M1008_g N_Y_c_540_n 0.0130095f $X=2.195 $Y=1.075 $X2=2.265
+ $Y2=1.48
cc_275 N_A_27_617#_c_301_n N_Y_c_542_n 0.0121767f $X=1.84 $Y=1.845 $X2=2.265
+ $Y2=2.59
cc_276 N_A_27_617#_c_341_n N_Y_c_542_n 0.0158479f $X=1.765 $Y=2.885 $X2=2.265
+ $Y2=2.59
cc_277 N_A_27_617#_M1008_g N_Y_c_543_n 0.00251111f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_278 N_A_27_617#_c_307_n N_Y_c_543_n 0.0177725f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.475
cc_279 N_A_27_617#_M1010_g N_Y_c_543_n 0.00251111f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=2.475
cc_280 N_A_27_617#_c_320_n N_Y_c_543_n 0.00843025f $X=3.055 $Y=2.81 $X2=2.41
+ $Y2=2.475
cc_281 N_A_27_617#_M1010_g N_Y_c_544_n 0.0130095f $X=2.625 $Y=1.075 $X2=3.125
+ $Y2=1.48
cc_282 N_A_27_617#_c_313_n N_Y_c_544_n 0.00213861f $X=2.98 $Y=1.845 $X2=3.125
+ $Y2=1.48
cc_283 N_A_27_617#_M1012_g N_Y_c_544_n 0.0136594f $X=3.055 $Y=1.075 $X2=3.125
+ $Y2=1.48
cc_284 N_A_27_617#_M1008_g N_Y_c_546_n 0.00259902f $X=2.195 $Y=1.075 $X2=2.555
+ $Y2=1.48
cc_285 N_A_27_617#_M1010_g N_Y_c_546_n 0.00259902f $X=2.625 $Y=1.075 $X2=2.555
+ $Y2=1.48
cc_286 N_A_27_617#_c_320_n N_Y_c_549_n 0.0155956f $X=3.055 $Y=2.81 $X2=3.125
+ $Y2=2.59
cc_287 N_A_27_617#_c_344_n N_Y_c_549_n 0.00894336f $X=2.625 $Y=1.845 $X2=3.125
+ $Y2=2.59
cc_288 N_A_27_617#_c_345_n N_Y_c_549_n 0.00903839f $X=2.625 $Y=2.885 $X2=3.125
+ $Y2=2.59
cc_289 N_A_27_617#_c_307_n N_Y_c_550_n 0.00140336f $X=2.55 $Y=1.845 $X2=2.555
+ $Y2=2.59
cc_290 N_A_27_617#_c_320_n N_Y_c_550_n 0.0012308f $X=3.055 $Y=2.81 $X2=2.555
+ $Y2=2.59
cc_291 N_A_27_617#_c_342_n N_Y_c_550_n 0.00140336f $X=2.195 $Y=1.845 $X2=2.555
+ $Y2=2.59
cc_292 N_A_27_617#_c_343_n N_Y_c_550_n 0.00372651f $X=2.195 $Y=2.885 $X2=2.555
+ $Y2=2.59
cc_293 N_A_27_617#_M1012_g N_Y_c_551_n 0.00262362f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_294 N_A_27_617#_M1014_g N_Y_c_551_n 0.00394441f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_295 N_A_27_617#_M1016_g N_Y_c_551_n 2.43068e-19 $X=3.915 $Y=1.075 $X2=3.27
+ $Y2=1.595
cc_296 N_A_27_617#_M1012_g N_Y_c_554_n 0.00251111f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=2.475
cc_297 N_A_27_617#_c_320_n N_Y_c_554_n 0.0108556f $X=3.055 $Y=2.81 $X2=3.27
+ $Y2=2.475
cc_298 N_A_27_617#_c_321_n N_Y_c_554_n 0.0177725f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=2.475
cc_299 N_A_27_617#_M1014_g N_Y_c_554_n 0.00251111f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=2.475
cc_300 N_A_27_617#_c_348_n N_Y_c_555_n 0.0121767f $X=3.485 $Y=1.845 $X2=3.985
+ $Y2=2.59
cc_301 N_A_27_617#_c_349_n N_Y_c_555_n 0.0158479f $X=3.485 $Y=2.885 $X2=3.985
+ $Y2=2.59
cc_302 N_A_27_617#_c_320_n N_Y_c_556_n 0.00618817f $X=3.055 $Y=2.81 $X2=3.415
+ $Y2=2.59
cc_303 N_A_27_617#_c_321_n N_Y_c_556_n 0.00268861f $X=3.41 $Y=1.845 $X2=3.415
+ $Y2=2.59
cc_304 N_A_27_617#_c_322_n N_Y_c_556_n 0.00357274f $X=3.41 $Y=2.885 $X2=3.415
+ $Y2=2.59
cc_305 N_A_27_617#_M1016_g N_Y_c_557_n 0.00259902f $X=3.915 $Y=1.075 $X2=4.13
+ $Y2=1.595
cc_306 N_A_27_617#_M1018_g N_Y_c_557_n 0.00954936f $X=4.345 $Y=1.075 $X2=4.13
+ $Y2=1.595
cc_307 N_A_27_617#_M1016_g N_Y_c_560_n 0.00251111f $X=3.915 $Y=1.075 $X2=4.13
+ $Y2=2.475
cc_308 N_A_27_617#_c_334_n N_Y_c_560_n 0.0184054f $X=4.27 $Y=1.845 $X2=4.13
+ $Y2=2.475
cc_309 N_A_27_617#_M1018_g N_Y_c_560_n 0.00251111f $X=4.345 $Y=1.075 $X2=4.13
+ $Y2=2.475
cc_310 N_A_27_617#_c_350_n N_Y_c_560_n 0.00140336f $X=3.915 $Y=1.845 $X2=4.13
+ $Y2=2.475
cc_311 N_A_27_617#_c_351_n N_Y_c_560_n 0.00372651f $X=3.915 $Y=2.885 $X2=4.13
+ $Y2=2.475
cc_312 N_A_27_617#_c_359_n N_Y_c_561_n 0.00226504f $X=1.335 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_313 N_A_27_617#_c_293_n N_Y_c_561_n 0.00744772f $X=1.37 $Y=2.81 $X2=1.55
+ $Y2=2.59
cc_314 N_A_27_617#_c_294_n N_Y_c_561_n 0.0156814f $X=1.69 $Y=2.885 $X2=1.55
+ $Y2=2.59
cc_315 N_A_27_617#_c_364_n N_Y_c_561_n 0.00392729f $X=1.765 $Y=2.96 $X2=1.55
+ $Y2=2.59
cc_316 N_A_27_617#_c_301_n N_Y_c_561_n 0.00182797f $X=1.84 $Y=1.845 $X2=1.55
+ $Y2=2.59
cc_317 N_A_27_617#_c_356_n N_Y_c_561_n 0.00273485f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=2.59
cc_318 N_A_27_617#_c_371_n N_Y_c_562_n 0.00392729f $X=2.195 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_319 N_A_27_617#_c_307_n N_Y_c_562_n 0.00250559f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=2.59
cc_320 N_A_27_617#_c_308_n N_Y_c_562_n 0.021445f $X=2.55 $Y=2.885 $X2=2.41
+ $Y2=2.59
cc_321 N_A_27_617#_c_376_n N_Y_c_562_n 0.00392729f $X=2.625 $Y=2.96 $X2=2.41
+ $Y2=2.59
cc_322 N_A_27_617#_c_320_n N_Y_c_562_n 0.00361281f $X=3.055 $Y=2.81 $X2=2.41
+ $Y2=2.59
cc_323 N_A_27_617#_c_320_n N_Y_c_563_n 0.00721971f $X=3.055 $Y=2.81 $X2=3.27
+ $Y2=2.59
cc_324 N_A_27_617#_c_382_n N_Y_c_563_n 0.00392729f $X=3.055 $Y=2.96 $X2=3.27
+ $Y2=2.59
cc_325 N_A_27_617#_c_321_n N_Y_c_563_n 0.00250559f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=2.59
cc_326 N_A_27_617#_c_322_n N_Y_c_563_n 0.021445f $X=3.41 $Y=2.885 $X2=3.27
+ $Y2=2.59
cc_327 N_A_27_617#_c_387_n N_Y_c_563_n 0.00392729f $X=3.485 $Y=2.96 $X2=3.27
+ $Y2=2.59
cc_328 N_A_27_617#_M1014_g N_Y_c_564_n 8.84842e-19 $X=3.485 $Y=1.075 $X2=4.13
+ $Y2=1.48
cc_329 N_A_27_617#_c_327_n N_Y_c_564_n 0.00213861f $X=3.84 $Y=1.845 $X2=4.13
+ $Y2=1.48
cc_330 N_A_27_617#_M1016_g N_Y_c_564_n 0.0130426f $X=3.915 $Y=1.075 $X2=4.13
+ $Y2=1.48
cc_331 N_A_27_617#_c_393_n N_Y_c_566_n 0.00392729f $X=3.915 $Y=2.96 $X2=4.13
+ $Y2=2.59
cc_332 N_A_27_617#_c_334_n N_Y_c_566_n 0.00250559f $X=4.27 $Y=1.845 $X2=4.13
+ $Y2=2.59
cc_333 N_A_27_617#_c_335_n N_Y_c_566_n 0.0206674f $X=4.27 $Y=2.885 $X2=4.13
+ $Y2=2.59
cc_334 N_A_27_617#_c_398_n N_Y_c_566_n 0.00392729f $X=4.345 $Y=2.96 $X2=4.13
+ $Y2=2.59
cc_335 N_A_27_617#_M1002_g N_Y_c_567_n 0.00231637f $X=1.335 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_336 N_A_27_617#_M1005_g N_Y_c_567_n 0.00231637f $X=1.765 $Y=1.075 $X2=1.55
+ $Y2=0.825
cc_337 N_A_27_617#_c_301_n N_Y_c_567_n 0.00171364f $X=1.84 $Y=1.845 $X2=1.55
+ $Y2=0.825
cc_338 N_A_27_617#_c_356_n N_Y_c_567_n 0.00500271f $X=1.43 $Y=1.935 $X2=1.55
+ $Y2=0.825
cc_339 N_A_27_617#_M1008_g N_Y_c_571_n 0.00231637f $X=2.195 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_340 N_A_27_617#_c_307_n N_Y_c_571_n 0.00280419f $X=2.55 $Y=1.845 $X2=2.41
+ $Y2=0.825
cc_341 N_A_27_617#_M1010_g N_Y_c_571_n 0.00231637f $X=2.625 $Y=1.075 $X2=2.41
+ $Y2=0.825
cc_342 N_A_27_617#_M1012_g N_Y_c_576_n 0.00231637f $X=3.055 $Y=1.075 $X2=3.27
+ $Y2=0.825
cc_343 N_A_27_617#_c_321_n N_Y_c_576_n 0.00280419f $X=3.41 $Y=1.845 $X2=3.27
+ $Y2=0.825
cc_344 N_A_27_617#_M1014_g N_Y_c_576_n 0.00231637f $X=3.485 $Y=1.075 $X2=3.27
+ $Y2=0.825
cc_345 N_A_27_617#_M1016_g N_Y_c_581_n 0.00231637f $X=3.915 $Y=1.075 $X2=4.13
+ $Y2=0.825
cc_346 N_A_27_617#_c_334_n N_Y_c_581_n 0.00280419f $X=4.27 $Y=1.845 $X2=4.13
+ $Y2=0.825
cc_347 N_A_27_617#_M1018_g N_Y_c_581_n 0.00231637f $X=4.345 $Y=1.075 $X2=4.13
+ $Y2=0.825
