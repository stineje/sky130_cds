magic
tech sky130A
magscale 1 2
timestamp 1612373804
<< nwell >>
rect -9 529 199 1119
<< nmoslvt >>
rect 80 115 110 243
<< pmos >>
rect 80 565 110 965
<< ndiff >>
rect 27 215 80 243
rect 27 131 35 215
rect 69 131 80 215
rect 27 115 80 131
rect 110 215 163 243
rect 110 131 121 215
rect 155 131 163 215
rect 110 115 163 131
<< pdiff >>
rect 27 949 80 965
rect 27 605 35 949
rect 69 605 80 949
rect 27 565 80 605
rect 110 949 163 965
rect 110 605 121 949
rect 155 605 163 949
rect 110 565 163 605
<< ndiffc >>
rect 35 131 69 215
rect 121 131 155 215
<< pdiffc >>
rect 35 605 69 949
rect 121 605 155 949
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 1049 51 1083
rect 85 1049 109 1083
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 1049 85 1083
<< poly >>
rect 80 965 110 991
rect 80 381 110 565
rect 80 365 134 381
rect 80 331 90 365
rect 124 331 134 365
rect 80 315 134 331
rect 80 243 110 315
rect 80 89 110 115
<< polycont >>
rect 90 331 124 365
<< locali >>
rect 0 1089 198 1110
rect 0 1049 51 1089
rect 85 1049 198 1089
rect 35 949 69 1049
rect 35 589 69 605
rect 121 949 155 965
rect 121 557 155 605
rect 74 331 90 365
rect 124 331 155 365
rect 35 215 69 231
rect 35 61 69 131
rect 121 215 155 331
rect 121 115 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 1083 85 1089
rect 51 1055 85 1083
rect 121 523 155 557
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 1089 198 1110
rect 0 1055 51 1089
rect 85 1055 198 1089
rect 0 1049 198 1055
rect 94 557 167 563
rect 94 523 121 557
rect 155 523 167 557
rect 94 517 167 523
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel viali 138 540 138 540 1 Y
port 1 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 1062 68 1062 1 vdd
<< end >>
