* File: sky130_osu_sc_18T_ls__pcgate_1.pex.spice
* Created: Thu Mar 10 13:46:56 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%GND 1 2 3 4 5 6 85 89 91 98 100 107
+ 109 119 121 131 133 140 159 164 166 168 170 172 174 176 178 181
c180 131 0 1.97615e-19 $X=3.99 $Y=0.825
r181 178 181 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=5.02 $Y=0.152
+ $X2=5.7 $Y2=0.152
r182 176 178 0.454078 $w=3.05e-07 $l=9.75e-07 $layer=MET1_cond $X=4.045 $Y=0.152
+ $X2=5.02 $Y2=0.152
r183 174 176 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=3.365 $Y=0.152
+ $X2=4.045 $Y2=0.152
r184 172 174 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=2.685 $Y=0.152
+ $X2=3.365 $Y2=0.152
r185 170 172 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=2.005 $Y=0.152
+ $X2=2.685 $Y2=0.152
r186 168 170 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=1.32 $Y=0.152
+ $X2=2.005 $Y2=0.152
r187 166 168 0.314362 $w=3.05e-07 $l=6.75e-07 $layer=MET1_cond $X=0.645 $Y=0.152
+ $X2=1.32 $Y2=0.152
r188 164 166 0.430792 $w=3.05e-07 $l=9.25e-07 $layer=MET1_cond $X=-0.28 $Y=0.152
+ $X2=0.645 $Y2=0.152
r189 162 164 0.316225 $w=3.05e-07 $l=6.79e-07 $layer=MET1_cond $X=-0.959
+ $Y=0.152 $X2=-0.28 $Y2=0.152
r190 159 162 0.000465721 $w=3.05e-07 $l=1e-09 $layer=MET1_cond $X=-0.96 $Y=0.152
+ $X2=-0.959 $Y2=0.152
r191 138 140 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.73 $Y=0.305
+ $X2=5.73 $Y2=0.825
r192 129 131 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.99 $Y=0.305
+ $X2=3.99 $Y2=0.825
r193 122 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.152
+ $X2=2.52 $Y2=0.152
r194 117 150 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.52 $Y=0.305
+ $X2=2.52 $Y2=0.152
r195 117 119 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.52 $Y=0.305
+ $X2=2.52 $Y2=0.825
r196 110 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.152
+ $X2=0.77 $Y2=0.152
r197 109 150 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.152
+ $X2=2.52 $Y2=0.152
r198 105 149 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.77 $Y=0.305
+ $X2=0.77 $Y2=0.152
r199 105 107 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.77 $Y=0.305
+ $X2=0.77 $Y2=0.825
r200 101 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.095 $Y=0.152
+ $X2=-0.18 $Y2=0.152
r201 100 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.152
+ $X2=0.77 $Y2=0.152
r202 96 148 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=-0.18 $Y=0.305
+ $X2=-0.18 $Y2=0.152
r203 96 98 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=-0.18 $Y=0.305
+ $X2=-0.18 $Y2=0.825
r204 91 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.265 $Y=0.152
+ $X2=-0.18 $Y2=0.152
r205 87 89 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=-1.04 $Y=0.305
+ $X2=-1.04 $Y2=0.825
r206 85 181 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.7 $Y=0.19
+ $X2=5.7 $Y2=0.19
r207 85 162 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=-0.959 $Y=0.19
+ $X2=-0.959 $Y2=0.19
r208 85 138 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.73 $Y=0.152
+ $X2=5.73 $Y2=0.305
r209 85 133 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=0.152
+ $X2=5.645 $Y2=0.152
r210 85 129 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.99 $Y=0.152
+ $X2=3.99 $Y2=0.305
r211 85 121 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=0.152
+ $X2=3.905 $Y2=0.152
r212 85 134 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=0.152
+ $X2=4.075 $Y2=0.152
r213 85 87 4.35274 $w=1.7e-07 $l=1.98681e-07 $layer=LI1_cond $X=-1.145 $Y=0.152
+ $X2=-1.04 $Y2=0.305
r214 85 92 3.2055 $w=3.05e-07 $l=1.9e-07 $layer=LI1_cond $X=-1.145 $Y=0.152
+ $X2=-0.955 $Y2=0.152
r215 85 133 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=5.02 $Y=0.152
+ $X2=5.645 $Y2=0.152
r216 85 134 35.7068 $w=3.03e-07 $l=9.45e-07 $layer=LI1_cond $X=5.02 $Y=0.152
+ $X2=4.075 $Y2=0.152
r217 85 121 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.365 $Y=0.152
+ $X2=3.905 $Y2=0.152
r218 85 122 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=2.685 $Y=0.152
+ $X2=2.605 $Y2=0.152
r219 85 109 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.005 $Y=0.152
+ $X2=2.435 $Y2=0.152
r220 85 110 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.325 $Y=0.152
+ $X2=0.855 $Y2=0.152
r221 85 100 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=0.645 $Y=0.152
+ $X2=0.685 $Y2=0.152
r222 85 101 27.9609 $w=3.03e-07 $l=7.4e-07 $layer=LI1_cond $X=0.645 $Y=0.152
+ $X2=-0.095 $Y2=0.152
r223 85 91 0.52899 $w=3.03e-07 $l=1.4e-08 $layer=LI1_cond $X=-0.279 $Y=0.152
+ $X2=-0.265 $Y2=0.152
r224 85 92 25.5427 $w=3.03e-07 $l=6.76e-07 $layer=LI1_cond $X=-0.279 $Y=0.152
+ $X2=-0.955 $Y2=0.152
r225 6 140 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.59
+ $Y=0.575 $X2=5.73 $Y2=0.825
r226 5 131 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.85
+ $Y=0.575 $X2=3.99 $Y2=0.825
r227 4 119 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.38
+ $Y=0.575 $X2=2.52 $Y2=0.825
r228 3 107 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.575 $X2=0.77 $Y2=0.825
r229 2 98 91 $w=1.7e-07 $l=3.1265e-07 $layer=licon1_NDIFF $count=2 $X=-0.32
+ $Y=0.575 $X2=-0.179 $Y2=0.825
r230 1 89 91 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=2 $X=-1.165
+ $Y=0.575 $X2=-1.039 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%VDD 1 2 3 4 5 6 65 67 74 78 84 88 96
+ 100 108 112 116 120 127 141 143 148 150 152 154 156 158 160 162 166
r119 164 166 0.00232861 $w=3.05e-07 $l=5e-09 $layer=MET1_cond $X=5.7 $Y=6.507
+ $X2=5.705 $Y2=6.507
r120 162 164 0.314362 $w=3.05e-07 $l=6.75e-07 $layer=MET1_cond $X=5.025 $Y=6.507
+ $X2=5.7 $Y2=6.507
r121 160 162 0.456407 $w=3.05e-07 $l=9.8e-07 $layer=MET1_cond $X=4.045 $Y=6.507
+ $X2=5.025 $Y2=6.507
r122 158 160 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=3.365 $Y=6.507
+ $X2=4.045 $Y2=6.507
r123 156 158 0.314362 $w=3.05e-07 $l=6.75e-07 $layer=MET1_cond $X=2.69 $Y=6.507
+ $X2=3.365 $Y2=6.507
r124 154 156 0.319019 $w=3.05e-07 $l=6.85e-07 $layer=MET1_cond $X=2.005 $Y=6.507
+ $X2=2.69 $Y2=6.507
r125 152 154 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=1.325 $Y=6.507
+ $X2=2.005 $Y2=6.507
r126 150 152 0.316691 $w=3.05e-07 $l=6.8e-07 $layer=MET1_cond $X=0.645 $Y=6.507
+ $X2=1.325 $Y2=6.507
r127 148 150 0.428464 $w=3.05e-07 $l=9.2e-07 $layer=MET1_cond $X=-0.275 $Y=6.507
+ $X2=0.645 $Y2=6.507
r128 146 148 0.318553 $w=3.05e-07 $l=6.84e-07 $layer=MET1_cond $X=-0.959
+ $Y=6.507 $X2=-0.275 $Y2=6.507
r129 143 146 0.000465721 $w=3.05e-07 $l=1e-09 $layer=MET1_cond $X=-0.96 $Y=6.507
+ $X2=-0.959 $Y2=6.507
r130 127 130 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=5.8 $Y=3.795
+ $X2=5.8 $Y2=5.835
r131 125 141 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.8 $Y=6.355
+ $X2=5.8 $Y2=6.507
r132 125 130 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.8 $Y=6.355
+ $X2=5.8 $Y2=5.835
r133 123 164 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.7 $Y=6.47
+ $X2=5.7 $Y2=6.47
r134 121 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=6.507
+ $X2=4.94 $Y2=6.507
r135 121 123 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=5.025 $Y=6.507
+ $X2=5.7 $Y2=6.507
r136 120 141 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=6.507
+ $X2=5.8 $Y2=6.507
r137 120 123 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=5.715 $Y=6.507
+ $X2=5.7 $Y2=6.507
r138 116 119 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=4.94 $Y=4.135
+ $X2=4.94 $Y2=5.835
r139 114 140 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.94 $Y=6.355
+ $X2=4.94 $Y2=6.507
r140 114 119 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.94 $Y=6.355
+ $X2=4.94 $Y2=5.835
r141 113 138 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=6.507
+ $X2=3.99 $Y2=6.507
r142 112 140 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=6.507
+ $X2=4.94 $Y2=6.507
r143 112 113 29.4723 $w=3.03e-07 $l=7.8e-07 $layer=LI1_cond $X=4.855 $Y=6.507
+ $X2=4.075 $Y2=6.507
r144 108 111 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.99 $Y=3.455
+ $X2=3.99 $Y2=5.835
r145 106 138 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.99 $Y=6.355
+ $X2=3.99 $Y2=6.507
r146 106 111 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.99 $Y=6.355
+ $X2=3.99 $Y2=5.835
r147 103 105 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=2.685 $Y=6.507
+ $X2=3.365 $Y2=6.507
r148 101 136 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=6.507
+ $X2=2.52 $Y2=6.507
r149 101 103 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=2.605 $Y=6.507
+ $X2=2.685 $Y2=6.507
r150 100 138 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=6.507
+ $X2=3.99 $Y2=6.507
r151 100 105 20.4039 $w=3.03e-07 $l=5.4e-07 $layer=LI1_cond $X=3.905 $Y=6.507
+ $X2=3.365 $Y2=6.507
r152 96 99 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.52 $Y=3.455
+ $X2=2.52 $Y2=5.835
r153 94 136 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.52 $Y=6.355
+ $X2=2.52 $Y2=6.507
r154 94 99 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.52 $Y=6.355
+ $X2=2.52 $Y2=5.835
r155 91 93 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.325 $Y=6.507
+ $X2=2.005 $Y2=6.507
r156 89 135 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=6.507
+ $X2=0.77 $Y2=6.507
r157 89 91 17.759 $w=3.03e-07 $l=4.7e-07 $layer=LI1_cond $X=0.855 $Y=6.507
+ $X2=1.325 $Y2=6.507
r158 88 136 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=6.507
+ $X2=2.52 $Y2=6.507
r159 88 93 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.435 $Y=6.507
+ $X2=2.005 $Y2=6.507
r160 84 87 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.77 $Y=3.795
+ $X2=0.77 $Y2=5.835
r161 82 135 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.77 $Y=6.355
+ $X2=0.77 $Y2=6.507
r162 82 87 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.77 $Y=6.355
+ $X2=0.77 $Y2=5.835
r163 79 134 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.165 $Y=6.507
+ $X2=-0.25 $Y2=6.507
r164 79 81 30.6059 $w=3.03e-07 $l=8.1e-07 $layer=LI1_cond $X=-0.165 $Y=6.507
+ $X2=0.645 $Y2=6.507
r165 78 135 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=6.507
+ $X2=0.77 $Y2=6.507
r166 78 81 1.5114 $w=3.03e-07 $l=4e-08 $layer=LI1_cond $X=0.685 $Y=6.507
+ $X2=0.645 $Y2=6.507
r167 74 77 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=-0.25 $Y=4.135
+ $X2=-0.25 $Y2=5.835
r168 72 134 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=-0.25 $Y=6.355
+ $X2=-0.25 $Y2=6.507
r169 72 77 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=-0.25 $Y=6.355
+ $X2=-0.25 $Y2=5.835
r170 69 146 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=-0.959 $Y=6.47
+ $X2=-0.959 $Y2=6.47
r171 67 134 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=-0.335 $Y=6.507
+ $X2=-0.25 $Y2=6.507
r172 67 69 23.5779 $w=3.03e-07 $l=6.24e-07 $layer=LI1_cond $X=-0.335 $Y=6.507
+ $X2=-0.959 $Y2=6.507
r173 65 123 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.495 $Y=6.355 $X2=5.7 $Y2=6.44
r174 65 140 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.815 $Y=6.355 $X2=5.02 $Y2=6.44
r175 65 138 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.84 $Y=6.355 $X2=4.045 $Y2=6.44
r176 65 105 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.16 $Y=6.355 $X2=3.365 $Y2=6.44
r177 65 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.48 $Y=6.355 $X2=2.685 $Y2=6.44
r178 65 93 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.8 $Y=6.355 $X2=2.005 $Y2=6.44
r179 65 91 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.12 $Y=6.355 $X2=1.325 $Y2=6.44
r180 65 81 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.44 $Y=6.355 $X2=0.645 $Y2=6.44
r181 65 134 182 $w=1.7e-07 $l=2.44839e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=-0.485 $Y=6.355 $X2=-0.279 $Y2=6.44
r182 65 69 182 $w=1.7e-07 $l=2.44839e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=-1.165 $Y=6.355 $X2=-0.959 $Y2=6.44
r183 6 130 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3
+ $X=5.66 $Y=3.085 $X2=5.8 $Y2=5.835
r184 6 127 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3
+ $X=5.66 $Y=3.085 $X2=5.8 $Y2=3.795
r185 5 119 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=4.815
+ $Y=3.085 $X2=4.94 $Y2=5.835
r186 5 116 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=4.815
+ $Y=3.085 $X2=4.94 $Y2=4.135
r187 4 111 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.85
+ $Y=3.085 $X2=3.99 $Y2=5.835
r188 4 108 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.85
+ $Y=3.085 $X2=3.99 $Y2=3.455
r189 3 99 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.38
+ $Y=3.085 $X2=2.52 $Y2=5.835
r190 3 96 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.38
+ $Y=3.085 $X2=2.52 $Y2=3.455
r191 2 87 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.63
+ $Y=3.085 $X2=0.77 $Y2=5.835
r192 2 84 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.63
+ $Y=3.085 $X2=0.77 $Y2=3.795
r193 1 77 200 $w=1.7e-07 $l=2.81962e-06 $layer=licon1_PDIFF $count=3 $X=-0.39
+ $Y=3.085 $X2=-0.249 $Y2=5.835
r194 1 74 200 $w=1.7e-07 $l=1.11828e-06 $layer=licon1_PDIFF $count=3 $X=-0.39
+ $Y=3.085 $X2=-0.249 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%SE 3 7 10 13 19 22 24
r51 24 26 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=-0.654 $Y=2.96
+ $X2=-0.649 $Y2=2.96
r52 22 24 0.000586854 $w=2.13e-07 $l=1e-09 $layer=MET1_cond $X=-0.655 $Y=2.96
+ $X2=-0.654 $Y2=2.96
r53 19 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-0.649 $Y=2.96
+ $X2=-0.649 $Y2=2.96
r54 17 19 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=-0.65 $Y=2.175
+ $X2=-0.65 $Y2=2.96
r55 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=-0.735 $Y=2.09
+ $X2=-0.65 $Y2=2.175
r56 13 15 9.72086 $w=1.68e-07 $l=1.49e-07 $layer=LI1_cond $X=-0.735 $Y=2.09
+ $X2=-0.884 $Y2=2.09
r57 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=-0.884
+ $Y=2.09 $X2=-0.884 $Y2=2.09
r58 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.885 $Y=2.09
+ $X2=-0.885 $Y2=2.255
r59 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.885 $Y=2.09
+ $X2=-0.885 $Y2=1.925
r60 7 12 1194.74 $w=1.5e-07 $l=2.33e-06 $layer=POLY_cond $X=-0.825 $Y=4.585
+ $X2=-0.825 $Y2=2.255
r61 3 11 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=-0.825 $Y=1.075
+ $X2=-0.825 $Y2=1.925
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%E 3 7 10 14 22
r47 20 22 0.001703 $w=3.67e-07 $l=5e-09 $layer=MET1_cond $X=-0.362 $Y=3.33
+ $X2=-0.362 $Y2=3.335
r48 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-0.309 $Y=3.33
+ $X2=-0.309 $Y2=3.33
r49 14 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=-0.31 $Y=2.755
+ $X2=-0.31 $Y2=3.33
r50 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=-0.309
+ $Y=2.755 $X2=-0.309 $Y2=2.755
r51 10 12 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.357 $Y=2.755
+ $X2=-0.357 $Y2=2.92
r52 10 11 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=-0.357 $Y=2.755
+ $X2=-0.357 $Y2=2.59
r53 7 11 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=-0.395 $Y=1.075
+ $X2=-0.395 $Y2=2.59
r54 3 12 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=-0.465 $Y=4.585
+ $X2=-0.465 $Y2=2.92
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_86_337# 1 3 13 16 18 19 21 22 23 24
+ 25 27 28 30 31 32 35 39
r86 39 41 80.671 $w=3.38e-07 $l=2.38e-06 $layer=LI1_cond $X=1.645 $Y=3.455
+ $X2=1.645 $Y2=5.835
r87 37 39 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=1.645 $Y=3.27
+ $X2=1.645 $Y2=3.455
r88 33 35 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=1.645 $Y=1.345
+ $X2=1.645 $Y2=0.825
r89 31 33 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.475 $Y=1.43
+ $X2=1.645 $Y2=1.345
r90 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.475 $Y=1.43
+ $X2=1.195 $Y2=1.43
r91 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.11 $Y=1.515
+ $X2=1.195 $Y2=1.43
r92 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.11 $Y=1.515
+ $X2=1.11 $Y2=1.765
r93 27 37 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.475 $Y=3.185
+ $X2=1.645 $Y2=3.27
r94 27 28 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.475 $Y=3.185
+ $X2=0.65 $Y2=3.185
r95 26 44 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.65 $Y=1.85
+ $X2=0.565 $Y2=1.81
r96 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.025 $Y=1.85
+ $X2=1.11 $Y2=1.765
r97 25 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.025 $Y=1.85
+ $X2=0.65 $Y2=1.85
r98 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=3.1
+ $X2=0.65 $Y2=3.185
r99 23 44 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=1.935
+ $X2=0.565 $Y2=1.81
r100 23 24 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=0.565 $Y=1.935
+ $X2=0.565 $Y2=3.1
r101 21 22 56.3681 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=0.53 $Y=2.805
+ $X2=0.53 $Y2=2.975
r102 20 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.505 $Y=2.015
+ $X2=0.505 $Y2=2.805
r103 18 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.85 $X2=0.565 $Y2=1.85
r104 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.85
+ $X2=0.565 $Y2=2.015
r105 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.85
+ $X2=0.565 $Y2=1.685
r106 16 22 517.347 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=0.555 $Y=4.585
+ $X2=0.555 $Y2=2.975
r107 13 19 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.555 $Y=1.075
+ $X2=0.555 $Y2=1.685
r108 3 41 150 $w=1.7e-07 $l=2.86029e-06 $layer=licon1_PDIFF $count=4 $X=1.42
+ $Y=3.085 $X2=1.645 $Y2=5.835
r109 3 39 150 $w=1.7e-07 $l=4.69201e-07 $layer=licon1_PDIFF $count=4 $X=1.42
+ $Y=3.085 $X2=1.645 $Y2=3.455
r110 1 35 91 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.575 $X2=1.645 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_N233_617# 1 3 11 15 18 22 30 36 41
+ 42 44 51 53 55 56
c111 36 0 1.69728e-19 $X=0.925 $Y=2.425
c112 15 0 1.88247e-19 $X=0.985 $Y=4.585
c113 11 0 1.38221e-19 $X=0.985 $Y=1.075
r114 55 56 0.10183 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.925 $Y=2.595
+ $X2=0.78 $Y2=2.595
r115 46 53 0.0522905 $w=1.72e-07 $l=9.2e-08 $layer=MET1_cond $X=-0.525 $Y=2.592
+ $X2=-0.617 $Y2=2.592
r116 46 56 1.18114 $w=1.75e-07 $l=1.305e-06 $layer=MET1_cond $X=-0.525 $Y=2.592
+ $X2=0.78 $Y2=2.592
r117 44 53 0.0142949 $w=1.7e-07 $l=9.04323e-08 $layer=MET1_cond $X=-0.61
+ $Y=2.505 $X2=-0.617 $Y2=2.592
r118 43 51 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=-0.61 $Y=1.595
+ $X2=-0.61 $Y2=1.48
r119 43 44 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=-0.61 $Y=1.595
+ $X2=-0.61 $Y2=2.505
r120 42 48 0.102734 $w=2.3e-07 $l=1.44e-07 $layer=MET1_cond $X=-0.895 $Y=2.59
+ $X2=-1.039 $Y2=2.59
r121 41 53 0.0522905 $w=1.72e-07 $l=9.39947e-08 $layer=MET1_cond $X=-0.71
+ $Y=2.59 $X2=-0.617 $Y2=2.592
r122 41 42 0.178133 $w=1.7e-07 $l=1.85e-07 $layer=MET1_cond $X=-0.71 $Y=2.59
+ $X2=-0.895 $Y2=2.59
r123 39 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.925 $Y=2.595
+ $X2=0.925 $Y2=2.595
r124 36 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.925 $Y=2.425
+ $X2=0.925 $Y2=2.595
r125 33 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-0.609 $Y=1.48
+ $X2=-0.609 $Y2=1.48
r126 30 33 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=-0.61 $Y=0.825
+ $X2=-0.61 $Y2=1.48
r127 25 27 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=-1.04 $Y=3.455
+ $X2=-1.04 $Y2=5.835
r128 22 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=-1.039 $Y=2.59
+ $X2=-1.039 $Y2=2.59
r129 22 25 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=-1.04 $Y=2.59
+ $X2=-1.04 $Y2=3.455
r130 18 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.425 $X2=0.925 $Y2=2.425
r131 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.425
+ $X2=0.925 $Y2=2.59
r132 18 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.425
+ $X2=0.925 $Y2=2.26
r133 15 20 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=0.985 $Y=4.585
+ $X2=0.985 $Y2=2.59
r134 11 19 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.985 $Y=1.075
+ $X2=0.985 $Y2=2.26
r135 3 27 150 $w=1.7e-07 $l=2.81229e-06 $layer=licon1_PDIFF $count=4 $X=-1.165
+ $Y=3.085 $X2=-1.039 $Y2=5.835
r136 3 25 150 $w=1.7e-07 $l=4.28392e-07 $layer=licon1_PDIFF $count=4 $X=-1.165
+ $Y=3.085 $X2=-1.039 $Y2=3.455
r137 1 30 91 $w=1.7e-07 $l=3.1265e-07 $layer=licon1_NDIFF $count=2 $X=-0.75
+ $Y=0.575 $X2=-0.609 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%CK 3 7 8 10 13 15 19 23 26 30 31 33 34
+ 38 42 43 44 48 57 61 64 67 70 74
c194 67 0 1.69728e-19 $X=1.405 $Y=2.765
c195 57 0 2.90509e-19 $X=1.485 $Y=2.765
c196 44 0 1.38221e-19 $X=1.57 $Y=1.85
c197 42 0 1.88247e-19 $X=1.485 $Y=2.68
c198 33 0 1.9983e-19 $X=2.762 $Y=2.78
c199 26 0 3.61476e-21 $X=1.405 $Y=2.765
r200 67 68 0.0923295 $w=2.64e-07 $l=1.95e-07 $layer=MET1_cond $X=1.405 $Y=2.765
+ $X2=1.405 $Y2=2.96
r201 65 68 0.0339426 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.55 $Y=2.96
+ $X2=1.405 $Y2=2.96
r202 64 74 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.485 $Y=2.96
+ $X2=5.63 $Y2=2.96
r203 64 65 3.78894 $w=1.7e-07 $l=3.935e-06 $layer=MET1_cond $X=5.485 $Y=2.96
+ $X2=1.55 $Y2=2.96
r204 61 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.87 $Y=1.85
+ $X2=2.87 $Y2=1.85
r205 54 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.405 $Y=2.765
+ $X2=1.405 $Y2=2.765
r206 54 57 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.405 $Y=2.765
+ $X2=1.485 $Y2=2.765
r207 51 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.63 $Y=2.96
+ $X2=5.63 $Y2=2.96
r208 48 51 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.63 $Y=2.425
+ $X2=5.63 $Y2=2.96
r209 44 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.57 $Y=1.85
+ $X2=1.885 $Y2=1.85
r210 43 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.85
+ $X2=2.87 $Y2=1.85
r211 43 46 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.785 $Y=1.85
+ $X2=1.885 $Y2=1.85
r212 42 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=2.68
+ $X2=1.485 $Y2=2.765
r213 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=1.935
+ $X2=1.57 $Y2=1.85
r214 41 42 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.485 $Y=1.935
+ $X2=1.485 $Y2=2.68
r215 38 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=2.425 $X2=5.63 $Y2=2.425
r216 38 40 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=5.602 $Y=2.425
+ $X2=5.602 $Y2=2.59
r217 38 39 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=5.602 $Y=2.425
+ $X2=5.602 $Y2=2.26
r218 36 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.85 $X2=2.87 $Y2=1.85
r219 33 34 50.1409 $w=2.05e-07 $l=1.55e-07 $layer=POLY_cond $X=2.762 $Y=2.78
+ $X2=2.762 $Y2=2.935
r220 30 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=1.85 $X2=1.885 $Y2=1.85
r221 30 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.85
+ $X2=1.885 $Y2=1.685
r222 26 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=2.765 $X2=1.405 $Y2=2.765
r223 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=2.765
+ $X2=1.405 $Y2=2.93
r224 23 40 1022.97 $w=1.5e-07 $l=1.995e-06 $layer=POLY_cond $X=5.585 $Y=4.585
+ $X2=5.585 $Y2=2.59
r225 19 39 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=5.515 $Y=1.075
+ $X2=5.515 $Y2=2.26
r226 15 36 38.5334 $w=3.13e-07 $l=1.84811e-07 $layer=POLY_cond $X=2.79 $Y=2.015
+ $X2=2.832 $Y2=1.85
r227 15 33 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.79 $Y=2.015
+ $X2=2.79 $Y2=2.78
r228 13 34 846.064 $w=1.5e-07 $l=1.65e-06 $layer=POLY_cond $X=2.735 $Y=4.585
+ $X2=2.735 $Y2=2.935
r229 8 36 41.6133 $w=3.13e-07 $l=2.28408e-07 $layer=POLY_cond $X=2.735 $Y=1.665
+ $X2=2.832 $Y2=1.85
r230 8 10 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.735 $Y=1.665
+ $X2=2.735 $Y2=1.075
r231 7 31 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.945 $Y=1.075
+ $X2=1.945 $Y2=1.685
r232 3 28 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.345 $Y=4.585
+ $X2=1.345 $Y2=2.93
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_254_89# 1 3 11 13 14 19 22 23 26 33
+ 37 44 47 51 53 54 59
c133 54 0 1.94649e-19 $X=2.03 $Y=2.59
c134 22 0 1.2087e-19 $X=1.885 $Y=2.765
c135 13 0 9.94742e-20 $X=1.75 $Y=2.3
r136 54 56 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.03 $Y=2.59
+ $X2=1.885 $Y2=2.59
r137 53 59 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.805 $Y=2.59
+ $X2=2.95 $Y2=2.59
r138 53 54 0.746234 $w=1.7e-07 $l=7.75e-07 $layer=MET1_cond $X=2.805 $Y=2.59
+ $X2=2.03 $Y2=2.59
r139 49 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.95 $Y=2.27
+ $X2=3.22 $Y2=2.27
r140 45 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.95 $Y=1.43
+ $X2=3.22 $Y2=1.43
r141 44 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.185
+ $X2=3.22 $Y2=2.27
r142 43 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.515
+ $X2=3.22 $Y2=1.43
r143 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.22 $Y=1.515
+ $X2=3.22 $Y2=2.185
r144 39 41 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.95 $Y=3.455
+ $X2=2.95 $Y2=5.835
r145 37 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.95 $Y=2.59
+ $X2=2.95 $Y2=2.59
r146 37 39 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.95 $Y=2.59
+ $X2=2.95 $Y2=3.455
r147 35 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=2.355
+ $X2=2.95 $Y2=2.27
r148 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.95 $Y=2.355
+ $X2=2.95 $Y2=2.59
r149 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=1.345
+ $X2=2.95 $Y2=1.43
r150 31 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.95 $Y=1.345
+ $X2=2.95 $Y2=0.825
r151 26 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.885 $Y=2.59
+ $X2=1.885 $Y2=2.59
r152 26 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.885 $Y=2.59
+ $X2=1.885 $Y2=2.765
r153 22 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=2.765 $X2=1.885 $Y2=2.765
r154 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=2.765
+ $X2=1.885 $Y2=2.93
r155 22 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=2.765
+ $X2=1.885 $Y2=2.6
r156 19 24 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=1.945 $Y=4.585
+ $X2=1.945 $Y2=2.93
r157 15 23 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.825 $Y=2.375
+ $X2=1.825 $Y2=2.6
r158 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.75 $Y=2.3
+ $X2=1.825 $Y2=2.375
r159 13 14 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.75 $Y=2.3
+ $X2=1.42 $Y2=2.3
r160 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=2.225
+ $X2=1.42 $Y2=2.3
r161 9 11 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=1.345 $Y=2.225
+ $X2=1.345 $Y2=1.075
r162 3 41 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.81
+ $Y=3.085 $X2=2.95 $Y2=5.835
r163 3 39 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.81
+ $Y=3.085 $X2=2.95 $Y2=3.455
r164 1 33 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.81
+ $Y=0.575 $X2=2.95 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_43_115# 1 3 11 15 23 26 28 32 33 35
+ 36 37 38 42 45 49 54 59 65 68 73 74 78 81 83
c181 81 0 1.2087e-19 $X=2.22 $Y=2.22
c182 59 0 1.9983e-19 $X=3.66 $Y=2.22
c183 32 0 2.20611e-19 $X=3.66 $Y=2.22
r184 80 81 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.365 $Y=2.22
+ $X2=2.22 $Y2=2.22
r185 78 81 2.2896 $w=1.4e-07 $l=1.85e-06 $layer=MET1_cond $X=0.37 $Y=2.2
+ $X2=2.22 $Y2=2.2
r186 76 78 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.225 $Y=2.22
+ $X2=0.37 $Y2=2.22
r187 74 80 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=2.515 $Y=2.22
+ $X2=2.365 $Y2=2.22
r188 73 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.515 $Y=2.22
+ $X2=3.66 $Y2=2.22
r189 73 74 1.23762 $w=1.4e-07 $l=1e-06 $layer=MET1_cond $X=3.515 $Y=2.22
+ $X2=2.515 $Y2=2.22
r190 68 70 8.33135 $w=2.83e-07 $l=1.6e-07 $layer=LI1_cond $X=0.282 $Y=3.795
+ $X2=0.282 $Y2=3.955
r191 68 69 12.1728 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.282 $Y=3.795
+ $X2=0.282 $Y2=3.54
r192 63 65 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.225 $Y=1.395
+ $X2=0.34 $Y2=1.395
r193 59 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.66 $Y=2.22
+ $X2=3.66 $Y2=2.22
r194 54 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.365 $Y=2.22
+ $X2=2.365 $Y2=2.22
r195 49 51 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.34 $Y=4.135
+ $X2=0.34 $Y2=5.835
r196 49 70 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.34 $Y=4.135
+ $X2=0.34 $Y2=3.955
r197 43 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=1.31
+ $X2=0.34 $Y2=1.395
r198 43 45 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.34 $Y=1.31
+ $X2=0.34 $Y2=0.825
r199 42 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.225 $Y=2.22
+ $X2=0.225 $Y2=2.22
r200 42 69 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.225 $Y=2.22
+ $X2=0.225 $Y2=3.54
r201 39 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=1.48
+ $X2=0.225 $Y2=1.395
r202 39 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.225 $Y=1.48
+ $X2=0.225 $Y2=2.22
r203 37 38 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.75 $Y=2.855
+ $X2=3.75 $Y2=3.005
r204 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.75 $Y=1.65 $X2=3.75
+ $Y2=1.8
r205 34 37 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.725 $Y=2.385
+ $X2=3.725 $Y2=2.855
r206 33 36 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.725 $Y=2.055
+ $X2=3.725 $Y2=1.8
r207 32 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=2.22 $X2=3.66 $Y2=2.22
r208 32 34 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.662 $Y=2.22
+ $X2=3.662 $Y2=2.385
r209 32 33 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.662 $Y=2.22
+ $X2=3.662 $Y2=2.055
r210 28 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=2.22 $X2=2.365 $Y2=2.22
r211 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=2.22
+ $X2=2.365 $Y2=2.385
r212 28 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=2.22
+ $X2=2.365 $Y2=2.055
r213 26 38 507.707 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=3.775 $Y=4.585
+ $X2=3.775 $Y2=3.005
r214 23 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.775 $Y=1.075
+ $X2=3.775 $Y2=1.65
r215 15 30 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=2.305 $Y=4.585
+ $X2=2.305 $Y2=2.385
r216 11 29 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.305 $Y=1.075
+ $X2=2.305 $Y2=2.055
r217 3 51 200 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.215
+ $Y=3.085 $X2=0.34 $Y2=5.835
r218 3 49 200 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=3 $X=0.215
+ $Y=3.085 $X2=0.34 $Y2=4.135
r219 3 68 600 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=3.085 $X2=0.34 $Y2=3.795
r220 1 45 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.575 $X2=0.34 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_687_115# 1 3 11 15 19 23 26 32 36 40
+ 46 47 48 49 53 55 60 61
c128 48 0 1.02575e-19 $X=4.06 $Y=2.765
c129 46 0 1.18035e-19 $X=4.06 $Y=1.85
c130 26 0 1.97615e-19 $X=4.145 $Y=2.22
r131 61 63 0.100167 $w=2.3e-07 $l=1.4e-07 $layer=MET1_cond $X=3.7 $Y=3.33
+ $X2=3.56 $Y2=3.33
r132 60 66 0.0905464 $w=2.13e-07 $l=1.45e-07 $layer=MET1_cond $X=4.805 $Y=3.33
+ $X2=4.95 $Y2=3.33
r133 60 61 1.06398 $w=1.7e-07 $l=1.105e-06 $layer=MET1_cond $X=4.805 $Y=3.33
+ $X2=3.7 $Y2=3.33
r134 58 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.95 $Y=3.33
+ $X2=4.95 $Y2=3.33
r135 55 58 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.95 $Y=2.765
+ $X2=4.95 $Y2=3.33
r136 51 53 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.145 $Y=2.68
+ $X2=4.145 $Y2=2.22
r137 50 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.145 $Y=1.935
+ $X2=4.145 $Y2=2.22
r138 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=2.765
+ $X2=4.145 $Y2=2.68
r139 48 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.06 $Y=2.765
+ $X2=3.645 $Y2=2.765
r140 46 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=1.85
+ $X2=4.145 $Y2=1.935
r141 46 47 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.06 $Y=1.85
+ $X2=3.645 $Y2=1.85
r142 42 44 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.56 $Y=3.455
+ $X2=3.56 $Y2=5.835
r143 40 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.56 $Y=3.33
+ $X2=3.56 $Y2=3.33
r144 40 42 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=3.33
+ $X2=3.56 $Y2=3.455
r145 38 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=2.85
+ $X2=3.645 $Y2=2.765
r146 38 40 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.56 $Y=2.85
+ $X2=3.56 $Y2=3.33
r147 34 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=1.765
+ $X2=3.645 $Y2=1.85
r148 34 36 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.56 $Y=1.765
+ $X2=3.56 $Y2=0.825
r149 30 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.95
+ $Y=2.765 $X2=4.95 $Y2=2.765
r150 30 32 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.95 $Y=2.765
+ $X2=5.155 $Y2=2.765
r151 26 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=2.22 $X2=4.145 $Y2=2.22
r152 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.145 $Y=2.22
+ $X2=4.145 $Y2=2.385
r153 26 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.145 $Y=2.22
+ $X2=4.145 $Y2=2.055
r154 21 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=2.93
+ $X2=5.155 $Y2=2.765
r155 21 23 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=5.155 $Y=2.93
+ $X2=5.155 $Y2=4.585
r156 17 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=2.6
+ $X2=5.155 $Y2=2.765
r157 17 19 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=5.155 $Y=2.6
+ $X2=5.155 $Y2=1.075
r158 15 28 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=4.205 $Y=4.585
+ $X2=4.205 $Y2=2.385
r159 11 27 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.205 $Y=1.075
+ $X2=4.205 $Y2=2.055
r160 3 44 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=3.435
+ $Y=3.085 $X2=3.56 $Y2=5.835
r161 3 42 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=3.435
+ $Y=3.085 $X2=3.56 $Y2=3.455
r162 1 36 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.575 $X2=3.56 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_963_115# 1 3 11 15 16 18 19 24 26 27
+ 32 36 38 39 40 43
r76 39 40 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.33 $Y=3.545
+ $X2=5.33 $Y2=3.715
r77 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=1.935
+ $X2=5.29 $Y2=1.935
r78 36 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=1.935
+ $X2=6.11 $Y2=1.935
r79 36 37 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.025 $Y=1.935
+ $X2=5.375 $Y2=1.935
r80 32 34 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=5.37 $Y=3.795
+ $X2=5.37 $Y2=5.835
r81 32 40 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=5.37 $Y=3.795 $X2=5.37
+ $Y2=3.715
r82 28 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=2.02 $X2=5.29
+ $Y2=1.935
r83 28 39 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=5.29 $Y=2.02
+ $X2=5.29 $Y2=3.545
r84 26 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=1.935
+ $X2=5.29 $Y2=1.935
r85 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.205 $Y=1.935
+ $X2=5.025 $Y2=1.935
r86 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.94 $Y=1.85
+ $X2=5.025 $Y2=1.935
r87 22 24 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=4.94 $Y=1.85
+ $X2=4.94 $Y2=0.825
r88 21 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.935 $X2=6.11 $Y2=1.935
r89 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=6.032 $Y=2.81
+ $X2=6.032 $Y2=2.96
r90 16 21 38.666 $w=2.85e-07 $l=1.84811e-07 $layer=POLY_cond $X=6.05 $Y=2.1
+ $X2=6.092 $Y2=1.935
r91 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.05 $Y=2.1 $X2=6.05
+ $Y2=2.81
r92 15 19 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=6.015 $Y=4.585
+ $X2=6.015 $Y2=2.96
r93 9 21 38.666 $w=2.85e-07 $l=1.99825e-07 $layer=POLY_cond $X=6.015 $Y=1.77
+ $X2=6.092 $Y2=1.935
r94 9 11 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.015 $Y=1.77
+ $X2=6.015 $Y2=1.075
r95 3 34 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=5.23
+ $Y=3.085 $X2=5.37 $Y2=5.835
r96 3 32 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=5.23
+ $Y=3.085 $X2=5.37 $Y2=3.795
r97 1 24 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=4.815
+ $Y=0.575 $X2=4.94 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%A_856_115# 1 3 11 15 22 24 26
r34 25 26 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.452 $Y=3.16
+ $X2=4.452 $Y2=3.33
r35 23 24 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.452 $Y=1.425
+ $X2=4.452 $Y2=1.595
r36 22 25 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=4.485 $Y=1.85
+ $X2=4.485 $Y2=3.16
r37 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.485 $Y=1.85
+ $X2=4.485 $Y2=1.595
r38 15 17 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.42 $Y=3.455
+ $X2=4.42 $Y2=5.835
r39 15 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.42 $Y=3.455
+ $X2=4.42 $Y2=3.33
r40 11 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.42 $Y=0.825 $X2=4.42
+ $Y2=1.425
r41 3 17 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=4.28
+ $Y=3.085 $X2=4.42 $Y2=5.835
r42 3 15 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=4.28
+ $Y=3.085 $X2=4.42 $Y2=3.455
r43 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=4.28
+ $Y=0.575 $X2=4.42 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__PCGATE_1%ECK 1 3 10 16 26 29 32
r33 24 32 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=6.23 $Y=2.475
+ $X2=6.23 $Y2=2.59
r34 24 26 0.250349 $w=1.7e-07 $l=2.6e-07 $layer=MET1_cond $X=6.23 $Y=2.475
+ $X2=6.23 $Y2=2.215
r35 23 29 0.0804477 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=6.23 $Y=1.595
+ $X2=6.23 $Y2=1.48
r36 23 26 0.596987 $w=1.7e-07 $l=6.2e-07 $layer=MET1_cond $X=6.23 $Y=1.595
+ $X2=6.23 $Y2=2.215
r37 19 21 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.23 $Y=3.455
+ $X2=6.23 $Y2=5.835
r38 16 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.23 $Y=2.59
+ $X2=6.23 $Y2=2.59
r39 16 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.23 $Y=2.59
+ $X2=6.23 $Y2=3.455
r40 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.23 $Y=1.48
+ $X2=6.23 $Y2=1.48
r41 10 13 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.23 $Y=0.825
+ $X2=6.23 $Y2=1.48
r42 3 21 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.09
+ $Y=3.085 $X2=6.23 $Y2=5.835
r43 3 19 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.09
+ $Y=3.085 $X2=6.23 $Y2=3.455
r44 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.09
+ $Y=0.575 $X2=6.23 $Y2=0.825
.ends

