* File: sky130_osu_sc_18T_ls__addf_1.pex.spice
* Created: Fri Nov 12 14:12:46 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%GND 1 2 3 4 5 81 83 91 93 103 105 112
+ 114 127 129 136 153 155
c182 127 0 1.91914e-19 $X=5.31 $Y=0.825
c183 103 0 1.85877e-19 $X=2.34 $Y=0.825
r184 153 155 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=6.46 $Y2=0.152
r185 138 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=0.152
+ $X2=6.32 $Y2=0.152
r186 134 149 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.152
r187 134 136 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.32 $Y=0.305
+ $X2=6.32 $Y2=0.825
r188 130 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.152
+ $X2=5.31 $Y2=0.152
r189 129 149 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.152
+ $X2=6.32 $Y2=0.152
r190 125 148 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.152
r191 125 127 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.31 $Y=0.305
+ $X2=5.31 $Y2=0.825
r192 115 147 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0.152
+ $X2=3.2 $Y2=0.152
r193 114 148 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=0.152
+ $X2=5.31 $Y2=0.152
r194 110 147 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.152
r195 110 112 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.2 $Y=0.305
+ $X2=3.2 $Y2=0.825
r196 105 147 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.152
+ $X2=3.2 $Y2=0.152
r197 101 103 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.34 $Y=0.305
+ $X2=2.34 $Y2=0.825
r198 94 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r199 89 143 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r200 89 91 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r201 83 143 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r202 81 155 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=0.19
+ $X2=6.46 $Y2=0.19
r203 81 153 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r204 81 101 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.34 $Y2=0.305
r205 81 93 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.255 $Y2=0.152
r206 81 106 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.152
+ $X2=2.425 $Y2=0.152
r207 81 138 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.46 $Y=0.152
+ $X2=6.405 $Y2=0.152
r208 81 129 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=6.235 $Y2=0.152
r209 81 130 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.78 $Y=0.152
+ $X2=5.395 $Y2=0.152
r210 81 114 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=0.152
+ $X2=5.225 $Y2=0.152
r211 81 115 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.285 $Y2=0.152
r212 81 105 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.115 $Y2=0.152
r213 81 106 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.425 $Y2=0.152
r214 81 93 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.255 $Y2=0.152
r215 81 94 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r216 81 83 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r217 5 136 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=6.195
+ $Y=0.575 $X2=6.32 $Y2=0.825
r218 4 127 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.17
+ $Y=0.575 $X2=5.31 $Y2=0.825
r219 3 112 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.575 $X2=3.2 $Y2=0.825
r220 2 103 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.2
+ $Y=0.575 $X2=2.34 $Y2=0.825
r221 1 91 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%VDD 1 2 3 4 5 61 63 70 74 82 86 92 96
+ 106 110 116 122 131 135
r110 131 135 2.85021 $w=3.05e-07 $l=6.12e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=6.46 $Y2=6.507
r111 122 135 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.46 $Y=6.47
+ $X2=6.46 $Y2=6.47
r112 120 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=6.507
+ $X2=6.32 $Y2=6.507
r113 120 122 2.2 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=6.405 $Y=6.507
+ $X2=6.46 $Y2=6.507
r114 116 119 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.32 $Y=3.455
+ $X2=6.32 $Y2=5.835
r115 114 129 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.32 $Y=6.355
+ $X2=6.32 $Y2=6.507
r116 114 119 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.32 $Y=6.355
+ $X2=6.32 $Y2=5.835
r117 111 128 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=6.507
+ $X2=5.31 $Y2=6.507
r118 111 113 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=5.395 $Y=6.507
+ $X2=5.78 $Y2=6.507
r119 110 129 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=6.507
+ $X2=6.32 $Y2=6.507
r120 110 113 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=6.235 $Y=6.507
+ $X2=5.78 $Y2=6.507
r121 106 109 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=5.31 $Y=4.135
+ $X2=5.31 $Y2=5.835
r122 104 128 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.31 $Y=6.355
+ $X2=5.31 $Y2=6.507
r123 104 109 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.31 $Y=6.355
+ $X2=5.31 $Y2=5.835
r124 101 103 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=4.42 $Y=6.507
+ $X2=5.1 $Y2=6.507
r125 99 101 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=3.74 $Y=6.507
+ $X2=4.42 $Y2=6.507
r126 97 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=6.507
+ $X2=3.2 $Y2=6.507
r127 97 99 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=3.285 $Y=6.507
+ $X2=3.74 $Y2=6.507
r128 96 128 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.31 $Y2=6.507
r129 96 103 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=5.225 $Y=6.507
+ $X2=5.1 $Y2=6.507
r130 92 95 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=3.2 $Y=4.135
+ $X2=3.2 $Y2=5.835
r131 90 127 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.2 $Y=6.355
+ $X2=3.2 $Y2=6.507
r132 90 95 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.2 $Y=6.355
+ $X2=3.2 $Y2=5.835
r133 87 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=6.507
+ $X2=2.34 $Y2=6.507
r134 87 89 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=2.425 $Y=6.507
+ $X2=3.06 $Y2=6.507
r135 86 127 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=6.507
+ $X2=3.2 $Y2=6.507
r136 86 89 2.07818 $w=3.03e-07 $l=5.5e-08 $layer=LI1_cond $X=3.115 $Y=6.507
+ $X2=3.06 $Y2=6.507
r137 82 85 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.34 $Y=3.795
+ $X2=2.34 $Y2=5.835
r138 80 126 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.34 $Y=6.355
+ $X2=2.34 $Y2=6.507
r139 80 85 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.34 $Y=6.355
+ $X2=2.34 $Y2=5.835
r140 77 79 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.02 $Y=6.507
+ $X2=1.7 $Y2=6.507
r141 75 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r142 75 77 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r143 74 126 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=6.507
+ $X2=2.34 $Y2=6.507
r144 74 79 20.9707 $w=3.03e-07 $l=5.55e-07 $layer=LI1_cond $X=2.255 $Y=6.507
+ $X2=1.7 $Y2=6.507
r145 70 73 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r146 68 124 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r147 68 73 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r148 65 131 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.34 $Y=6.47
+ $X2=0.34 $Y2=6.47
r149 63 124 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r150 63 65 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r151 61 122 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=6.255 $Y=6.355 $X2=6.46 $Y2=6.44
r152 61 113 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=5.575 $Y=6.355 $X2=5.78 $Y2=6.44
r153 61 103 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.895 $Y=6.355 $X2=5.1 $Y2=6.44
r154 61 101 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=4.215 $Y=6.355 $X2=4.42 $Y2=6.44
r155 61 99 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r156 61 89 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r157 61 126 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r158 61 79 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r159 61 77 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r160 61 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r161 5 119 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=6.195
+ $Y=3.085 $X2=6.32 $Y2=5.835
r162 5 116 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=6.195
+ $Y=3.085 $X2=6.32 $Y2=3.455
r163 4 109 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=5.17
+ $Y=3.085 $X2=5.31 $Y2=5.835
r164 4 106 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=5.17
+ $Y=3.085 $X2=5.31 $Y2=4.135
r165 3 95 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.06
+ $Y=3.085 $X2=3.2 $Y2=5.835
r166 3 92 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=3.06
+ $Y=3.085 $X2=3.2 $Y2=4.135
r167 2 85 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.2
+ $Y=3.085 $X2=2.34 $Y2=5.835
r168 2 82 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=2.2
+ $Y=3.085 $X2=2.34 $Y2=3.795
r169 1 73 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r170 1 70 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%A 3 6 8 10 11 13 14 15 16 17 19 22 23 25
+ 28 31 36 37 39 40 45 48 49 51 52 54 59 64 68 69 70 71 73 80
c207 80 0 1.91914e-19 $X=5.155 $Y=1.85
c208 71 0 1.85877e-19 $X=2.64 $Y=1.85
c209 69 0 1.24216e-19 $X=0.63 $Y=1.85
c210 68 0 1.77566e-19 $X=2.35 $Y=1.85
c211 52 0 2.67871e-19 $X=5.13 $Y=2.925
c212 31 0 1.32911e-19 $X=5.095 $Y=4.585
c213 19 0 1.74961e-19 $X=2.435 $Y=2.81
c214 14 0 9.53445e-20 $X=2.36 $Y=1.76
r215 71 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.64 $Y=1.85
+ $X2=2.495 $Y2=1.85
r216 70 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.01 $Y=1.85
+ $X2=5.155 $Y2=1.85
r217 70 71 2.28203 $w=1.7e-07 $l=2.37e-06 $layer=MET1_cond $X=5.01 $Y=1.85
+ $X2=2.64 $Y2=1.85
r218 69 73 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=1.85
+ $X2=0.485 $Y2=1.85
r219 68 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.35 $Y=1.85
+ $X2=2.495 $Y2=1.85
r220 68 69 1.65616 $w=1.7e-07 $l=1.72e-06 $layer=MET1_cond $X=2.35 $Y=1.85
+ $X2=0.63 $Y2=1.85
r221 64 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.155 $Y=1.85
+ $X2=5.155 $Y2=1.85
r222 59 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.495 $Y=1.85
+ $X2=2.495 $Y2=1.85
r223 54 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=1.85
r224 51 52 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=5.13 $Y=2.775
+ $X2=5.13 $Y2=2.925
r225 50 51 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.165 $Y=2.015
+ $X2=5.165 $Y2=2.775
r226 48 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.85 $X2=5.155 $Y2=1.85
r227 48 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.85
+ $X2=5.155 $Y2=2.015
r228 48 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.85
+ $X2=5.155 $Y2=1.685
r229 44 45 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.435 $Y=2.885
+ $X2=2.555 $Y2=2.885
r230 42 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.85 $X2=2.495 $Y2=1.85
r231 42 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.85
+ $X2=2.495 $Y2=2.015
r232 39 42 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.495 $Y=1.76
+ $X2=2.495 $Y2=1.85
r233 39 40 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.495 $Y=1.76
+ $X2=2.495 $Y2=1.685
r234 36 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.85 $X2=0.485 $Y2=1.85
r235 36 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=2.015
r236 36 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=1.685
r237 31 52 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=5.095 $Y=4.585
+ $X2=5.095 $Y2=2.925
r238 28 49 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.095 $Y=1.075
+ $X2=5.095 $Y2=1.685
r239 23 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.555 $Y=2.96
+ $X2=2.555 $Y2=2.885
r240 23 25 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.555 $Y=2.96
+ $X2=2.555 $Y2=4.585
r241 22 40 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.555 $Y=1.075
+ $X2=2.555 $Y2=1.685
r242 19 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=2.81
+ $X2=2.435 $Y2=2.885
r243 19 43 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.435 $Y=2.81
+ $X2=2.435 $Y2=2.015
r244 16 44 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=2.885
+ $X2=2.435 $Y2=2.885
r245 16 17 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=2.885
+ $X2=2.2 $Y2=2.885
r246 14 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.36 $Y=1.76
+ $X2=2.495 $Y2=1.76
r247 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.36 $Y=1.76
+ $X2=2.2 $Y2=1.76
r248 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=2.96
+ $X2=2.2 $Y2=2.885
r249 11 13 522.167 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=2.125 $Y=2.96
+ $X2=2.125 $Y2=4.585
r250 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=1.685
+ $X2=2.2 $Y2=1.76
r251 8 10 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.125 $Y=1.685
+ $X2=2.125 $Y2=1.075
r252 6 38 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.015
r253 3 37 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=1.685
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%B 3 7 11 15 19 22 26 30 33 39 42 43 46
+ 51 55 58 64 69 74 78 79 81 83 84 85 86
c230 86 0 6.46001e-20 $X=3.67 $Y=2.592
c231 69 0 1.26882e-19 $X=0.485 $Y=2.59
c232 55 0 9.53445e-20 $X=2.305 $Y=2.59
r233 86 93 0.459737 $w=1.9e-07 $l=6.95999e-07 $layer=MET1_cond $X=3.67 $Y=2.592
+ $X2=2.975 $Y2=2.59
r234 85 95 0.124897 $w=2.19e-07 $l=2.05998e-07 $layer=MET1_cond $X=4.06 $Y=2.592
+ $X2=4.265 $Y2=2.59
r235 85 86 0.386904 $w=1.65e-07 $l=3.9e-07 $layer=MET1_cond $X=4.06 $Y=2.592
+ $X2=3.67 $Y2=2.592
r236 84 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.45 $Y=2.59
+ $X2=2.305 $Y2=2.59
r237 83 93 0.0970649 $w=1.9e-07 $l=1.45e-07 $layer=MET1_cond $X=2.83 $Y=2.59
+ $X2=2.975 $Y2=2.59
r238 83 84 0.365895 $w=1.7e-07 $l=3.8e-07 $layer=MET1_cond $X=2.83 $Y=2.59
+ $X2=2.45 $Y2=2.59
r239 79 88 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.63 $Y=2.59
+ $X2=0.485 $Y2=2.59
r240 79 81 0.0144432 $w=1.7e-07 $l=1.5e-08 $layer=MET1_cond $X=0.63 $Y=2.59
+ $X2=0.645 $Y2=2.59
r241 78 91 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.16 $Y=2.59
+ $X2=2.305 $Y2=2.59
r242 78 81 1.45877 $w=1.7e-07 $l=1.515e-06 $layer=MET1_cond $X=2.16 $Y=2.59
+ $X2=0.645 $Y2=2.59
r243 74 76 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.015 $Y=2.43
+ $X2=2.015 $Y2=2.59
r244 69 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.485 $Y=2.59
+ $X2=0.485 $Y2=2.59
r245 69 71 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.485 $Y=2.59
+ $X2=0.485 $Y2=2.76
r246 64 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.265 $Y=2.59
+ $X2=4.265 $Y2=2.59
r247 61 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=2.59
+ $X2=2.975 $Y2=2.59
r248 58 61 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.975 $Y=1.85
+ $X2=2.975 $Y2=2.59
r249 55 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.305 $Y=2.59
+ $X2=2.305 $Y2=2.59
r250 53 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.59
+ $X2=2.015 $Y2=2.59
r251 53 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.1 $Y=2.59
+ $X2=2.305 $Y2=2.59
r252 49 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=2.76
+ $X2=0.485 $Y2=2.76
r253 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.57 $Y=2.76
+ $X2=0.895 $Y2=2.76
r254 46 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=2.59 $X2=4.265 $Y2=2.59
r255 46 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.59
+ $X2=4.265 $Y2=2.755
r256 46 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=2.59
+ $X2=4.265 $Y2=2.425
r257 42 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.85 $X2=2.975 $Y2=1.85
r258 42 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.85
+ $X2=2.975 $Y2=2.015
r259 42 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.85
+ $X2=2.975 $Y2=1.685
r260 39 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=2.43 $X2=2.015 $Y2=2.43
r261 36 39 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.765 $Y=2.43
+ $X2=2.015 $Y2=2.43
r262 33 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=2.76 $X2=0.895 $Y2=2.76
r263 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.76
+ $X2=0.895 $Y2=2.925
r264 33 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=2.76
+ $X2=0.895 $Y2=2.595
r265 30 48 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=4.275 $Y=4.585
+ $X2=4.275 $Y2=2.755
r266 26 47 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=4.275 $Y=1.075
+ $X2=4.275 $Y2=2.425
r267 22 44 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=2.985 $Y=4.585
+ $X2=2.985 $Y2=2.015
r268 19 43 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.985 $Y=1.075
+ $X2=2.985 $Y2=1.685
r269 13 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.595
+ $X2=1.765 $Y2=2.43
r270 13 15 1020.4 $w=1.5e-07 $l=1.99e-06 $layer=POLY_cond $X=1.765 $Y=2.595
+ $X2=1.765 $Y2=4.585
r271 9 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.265
+ $X2=1.765 $Y2=2.43
r272 9 11 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=1.765 $Y=2.265
+ $X2=1.765 $Y2=1.075
r273 7 35 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=0.905 $Y=4.585
+ $X2=0.905 $Y2=2.925
r274 3 34 779.404 $w=1.5e-07 $l=1.52e-06 $layer=POLY_cond $X=0.905 $Y=1.075
+ $X2=0.905 $Y2=2.595
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%CI 3 7 11 15 19 23 26 30 32 36 42 45 51
+ 55 56 57 58 60 66
c184 56 0 3.15979e-20 $X=1.47 $Y=2.22
c185 11 0 1.47588e-19 $X=3.415 $Y=1.075
c186 7 0 1.26882e-19 $X=1.335 $Y=4.585
r187 58 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.56 $Y=2.22
+ $X2=3.415 $Y2=2.22
r188 57 66 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.6 $Y=2.22
+ $X2=4.745 $Y2=2.22
r189 57 58 1.0014 $w=1.7e-07 $l=1.04e-06 $layer=MET1_cond $X=4.6 $Y=2.22
+ $X2=3.56 $Y2=2.22
r190 56 60 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.47 $Y=2.22
+ $X2=1.325 $Y2=2.22
r191 55 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.27 $Y=2.22
+ $X2=3.415 $Y2=2.22
r192 55 56 1.73319 $w=1.7e-07 $l=1.8e-06 $layer=MET1_cond $X=3.27 $Y=2.22
+ $X2=1.47 $Y2=2.22
r193 45 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.745 $Y=2.22
+ $X2=4.745 $Y2=2.22
r194 45 48 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.745 $Y=2.22
+ $X2=4.745 $Y2=2.4
r195 42 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.415 $Y=2.22
+ $X2=3.415 $Y2=2.22
r196 40 51 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=2.505
+ $X2=3.415 $Y2=2.59
r197 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.415 $Y=2.505
+ $X2=3.415 $Y2=2.22
r198 36 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.325 $Y=2.22
+ $X2=1.325 $Y2=2.22
r199 32 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=2.4 $X2=4.745 $Y2=2.4
r200 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=2.4
+ $X2=4.745 $Y2=2.565
r201 32 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=2.4
+ $X2=4.745 $Y2=2.235
r202 30 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=2.59 $X2=3.415 $Y2=2.59
r203 26 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=2.22 $X2=1.325 $Y2=2.22
r204 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.22
+ $X2=1.325 $Y2=2.385
r205 26 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=2.22
+ $X2=1.325 $Y2=2.055
r206 23 34 1035.79 $w=1.5e-07 $l=2.02e-06 $layer=POLY_cond $X=4.685 $Y=4.585
+ $X2=4.685 $Y2=2.565
r207 19 33 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=4.685 $Y=1.075
+ $X2=4.685 $Y2=2.235
r208 13 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.755
+ $X2=3.415 $Y2=2.59
r209 13 15 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.415 $Y=2.755
+ $X2=3.415 $Y2=4.585
r210 9 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=2.425
+ $X2=3.415 $Y2=2.59
r211 9 11 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=3.415 $Y=2.425
+ $X2=3.415 $Y2=1.075
r212 7 28 1128.09 $w=1.5e-07 $l=2.2e-06 $layer=POLY_cond $X=1.335 $Y=4.585
+ $X2=1.335 $Y2=2.385
r213 3 27 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=2.055
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%CON 1 3 9 11 14 18 22 25 27 32 38 43 46
+ 50 54 58 63 68 70 71 72 73 80
c192 73 0 1.47588e-19 $X=4.115 $Y=1.48
c193 54 0 3.15979e-20 $X=1.665 $Y=1.765
c194 43 0 1.74961e-19 $X=1.665 $Y=3.025
c195 32 0 1.77566e-19 $X=1.55 $Y=0.825
c196 27 0 1.71092e-19 $X=6.41 $Y=2.74
c197 25 0 1.22485e-19 $X=3.845 $Y=1.85
r198 73 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.115 $Y=1.48
+ $X2=3.97 $Y2=1.48
r199 72 80 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.995 $Y=1.48
+ $X2=6.14 $Y2=1.48
r200 72 73 1.81022 $w=1.7e-07 $l=1.88e-06 $layer=MET1_cond $X=5.995 $Y=1.48
+ $X2=4.115 $Y2=1.48
r201 71 75 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.48
+ $X2=1.55 $Y2=1.48
r202 70 78 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.825 $Y=1.48
+ $X2=3.97 $Y2=1.48
r203 70 71 2.05094 $w=1.7e-07 $l=2.13e-06 $layer=MET1_cond $X=3.825 $Y=1.48
+ $X2=1.695 $Y2=1.48
r204 66 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.14 $Y=1.48
+ $X2=6.14 $Y2=1.48
r205 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.14 $Y=1.48
+ $X2=6.41 $Y2=1.48
r206 61 63 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.85
+ $X2=3.97 $Y2=1.85
r207 56 58 6.89435 $w=1.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=3.117
+ $X2=1.665 $Y2=3.117
r208 52 54 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.55 $Y=1.765
+ $X2=1.665 $Y2=1.765
r209 48 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.565
+ $X2=6.41 $Y2=1.48
r210 48 50 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.41 $Y=1.565
+ $X2=6.41 $Y2=2.74
r211 46 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.97 $Y=1.48
+ $X2=3.97 $Y2=1.48
r212 44 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=1.765
+ $X2=3.97 $Y2=1.85
r213 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.97 $Y=1.765
+ $X2=3.97 $Y2=1.48
r214 43 58 1.22693 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=1.665 $Y=3.025
+ $X2=1.665 $Y2=3.117
r215 42 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.85
+ $X2=1.665 $Y2=1.765
r216 42 43 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.665 $Y=1.85
+ $X2=1.665 $Y2=3.025
r217 38 40 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.55 $Y=3.795
+ $X2=1.55 $Y2=5.835
r218 36 56 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.55 $Y=3.21
+ $X2=1.55 $Y2=3.117
r219 36 38 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.55 $Y=3.21
+ $X2=1.55 $Y2=3.795
r220 35 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.48
+ $X2=1.55 $Y2=1.48
r221 32 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.55 $Y2=1.48
r222 30 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.68
+ $X2=1.55 $Y2=1.765
r223 30 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.55 $Y=1.68 $X2=1.55
+ $Y2=1.48
r224 27 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=2.74 $X2=6.41 $Y2=2.74
r225 27 29 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.74
+ $X2=6.442 $Y2=2.905
r226 27 28 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.442 $Y=2.74
+ $X2=6.442 $Y2=2.575
r227 25 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.85 $X2=3.845 $Y2=1.85
r228 22 29 861.447 $w=1.5e-07 $l=1.68e-06 $layer=POLY_cond $X=6.535 $Y=4.585
+ $X2=6.535 $Y2=2.905
r229 18 28 769.149 $w=1.5e-07 $l=1.5e-06 $layer=POLY_cond $X=6.535 $Y=1.075
+ $X2=6.535 $Y2=2.575
r230 12 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=2.015
+ $X2=3.845 $Y2=1.85
r231 12 14 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=3.845 $Y=2.015
+ $X2=3.845 $Y2=4.585
r232 9 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.685
+ $X2=3.845 $Y2=1.85
r233 9 11 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.845 $Y=1.685
+ $X2=3.845 $Y2=1.075
r234 3 40 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r235 3 38 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.795
r236 1 32 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%A_784_115# 1 3 11 15 18 20 21 22 23 26
+ 28 32 35 37 40 43
c125 40 0 1.48211e-20 $X=4.31 $Y=0.99
c126 37 0 9.63581e-20 $X=5.415 $Y=3.25
c127 20 0 6.46001e-20 $X=3.845 $Y=3.03
c128 18 0 3.07391e-19 $X=5.585 $Y=2.755
c129 15 0 1.71513e-19 $X=5.585 $Y=4.585
c130 11 0 1.71092e-19 $X=5.585 $Y=1.075
r131 43 45 7.30282 $w=2.84e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=2.755
+ $X2=5.585 $Y2=2.755
r132 38 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.06 $Y=0.99
+ $X2=4.31 $Y2=0.99
r133 36 43 3.73949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=2.92
+ $X2=5.415 $Y2=2.755
r134 36 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.415 $Y=2.92
+ $X2=5.415 $Y2=3.25
r135 34 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=1.075
+ $X2=4.31 $Y2=0.99
r136 34 35 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=4.31 $Y=1.075
+ $X2=4.31 $Y2=2.135
r137 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.33 $Y=3.335
+ $X2=5.415 $Y2=3.25
r138 32 33 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=5.33 $Y=3.335
+ $X2=4.145 $Y2=3.335
r139 28 30 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=4.06 $Y=3.795
+ $X2=4.06 $Y2=5.835
r140 26 33 5.48216 $w=2.66e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=3.42
+ $X2=4.145 $Y2=3.335
r141 26 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.06 $Y=3.42
+ $X2=4.06 $Y2=3.795
r142 23 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=0.905
+ $X2=4.06 $Y2=0.99
r143 23 25 5.74118 $w=1.7e-07 $l=8e-08 $layer=LI1_cond $X=4.06 $Y=0.905 $X2=4.06
+ $Y2=0.825
r144 21 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.225 $Y=2.22
+ $X2=4.31 $Y2=2.135
r145 21 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.225 $Y=2.22
+ $X2=3.93 $Y2=2.22
r146 20 33 15.5724 $w=2.66e-07 $l=4.29564e-07 $layer=LI1_cond $X=3.845 $Y=3.03
+ $X2=4.145 $Y2=3.335
r147 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=2.305
+ $X2=3.93 $Y2=2.22
r148 19 20 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.845 $Y=2.305
+ $X2=3.845 $Y2=3.03
r149 18 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.585
+ $Y=2.755 $X2=5.585 $Y2=2.755
r150 13 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.92
+ $X2=5.585 $Y2=2.755
r151 13 15 853.755 $w=1.5e-07 $l=1.665e-06 $layer=POLY_cond $X=5.585 $Y=2.92
+ $X2=5.585 $Y2=4.585
r152 9 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=2.59
+ $X2=5.585 $Y2=2.755
r153 9 11 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=5.585 $Y=2.59
+ $X2=5.585 $Y2=1.075
r154 3 30 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.92
+ $Y=3.085 $X2=4.06 $Y2=5.835
r155 3 28 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=3.92
+ $Y=3.085 $X2=4.06 $Y2=3.795
r156 1 25 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.575 $X2=4.06 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%A_27_617# 1 2 11 15 19
r13 19 21 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.12 $Y=3.795
+ $X2=1.12 $Y2=5.835
r14 17 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.12 $Y=3.545
+ $X2=1.12 $Y2=3.795
r15 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=3.46
+ $X2=1.12 $Y2=3.545
r16 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=3.46
+ $X2=0.345 $Y2=3.46
r17 11 13 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=0.26 $Y=3.795
+ $X2=0.26 $Y2=5.835
r18 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.545
+ $X2=0.345 $Y2=3.46
r19 9 11 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.26 $Y=3.545
+ $X2=0.26 $Y2=3.795
r20 2 21 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r21 2 19 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.795
r22 1 13 171.429 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r23 1 11 171.429 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%A_526_617# 1 2 11 15 19
r12 19 21 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=3.63 $Y=3.795
+ $X2=3.63 $Y2=5.835
r13 17 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.63 $Y=3.54
+ $X2=3.63 $Y2=3.795
r14 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=3.455
+ $X2=3.63 $Y2=3.54
r15 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=3.455
+ $X2=2.855 $Y2=3.455
r16 11 13 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.77 $Y=3.795
+ $X2=2.77 $Y2=5.835
r17 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=3.54
+ $X2=2.855 $Y2=3.455
r18 9 11 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.77 $Y=3.54
+ $X2=2.77 $Y2=3.795
r19 2 21 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=3.49
+ $Y=3.085 $X2=3.63 $Y2=5.835
r20 2 19 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=3.49
+ $Y=3.085 $X2=3.63 $Y2=3.795
r21 1 13 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=2.63
+ $Y=3.085 $X2=2.77 $Y2=5.835
r22 1 11 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=2.63
+ $Y=3.085 $X2=2.77 $Y2=3.795
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%S 1 3 11 17 22 25 29 32
c49 32 0 1.32911e-19 $X=5.8 $Y=3.335
c50 29 0 1.41304e-19 $X=5.925 $Y=3.25
c51 25 0 1.66087e-19 $X=5.925 $Y=2.22
r52 27 29 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=3.25
+ $X2=5.925 $Y2=3.25
r53 23 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=2.22
+ $X2=5.925 $Y2=2.22
r54 22 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=3.165
+ $X2=5.925 $Y2=3.25
r55 21 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=2.305
+ $X2=5.925 $Y2=2.22
r56 21 22 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.925 $Y=2.305
+ $X2=5.925 $Y2=3.165
r57 17 19 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=5.8 $Y=3.795
+ $X2=5.8 $Y2=5.835
r58 15 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.8 $Y=3.335 $X2=5.8
+ $Y2=3.335
r59 15 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=3.335 $X2=5.8
+ $Y2=3.25
r60 15 17 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.8 $Y=3.335 $X2=5.8
+ $Y2=3.795
r61 9 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.135 $X2=5.8
+ $Y2=2.22
r62 9 11 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=5.8 $Y=2.135 $X2=5.8
+ $Y2=0.825
r63 3 19 171.429 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=5.66
+ $Y=3.085 $X2=5.8 $Y2=5.835
r64 3 17 171.429 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=3 $X=5.66
+ $Y=3.085 $X2=5.8 $Y2=3.795
r65 1 11 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=5.66
+ $Y=0.575 $X2=5.8 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%CO 1 3 10 20
r15 15 17 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.75 $Y=3.455
+ $X2=6.75 $Y2=5.835
r16 13 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.75 $Y=2.96
+ $X2=6.75 $Y2=2.96
r17 13 15 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.75 $Y=2.96
+ $X2=6.75 $Y2=3.455
r18 10 13 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=6.75 $Y=0.825
+ $X2=6.75 $Y2=2.96
r19 3 17 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=6.61
+ $Y=3.085 $X2=6.75 $Y2=5.835
r20 3 15 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=6.61
+ $Y=3.085 $X2=6.75 $Y2=3.455
r21 1 10 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=6.61
+ $Y=0.575 $X2=6.75 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%A_27_115# 1 2 11 13 14 17
c21 14 0 1.24216e-19 $X=0.345 $Y=1.345
r22 15 17 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.12 $Y=1.26
+ $X2=1.12 $Y2=0.825
r23 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.345
+ $X2=1.12 $Y2=1.26
r24 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.345
+ $X2=0.345 $Y2=1.345
r25 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.26
+ $X2=0.345 $Y2=1.345
r26 9 11 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=1.26
+ $X2=0.26 $Y2=0.825
r27 2 17 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
r28 1 11 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__ADDF_1%A_526_115# 1 2 11 13 14 17
c33 13 0 1.07664e-19 $X=3.545 $Y=1.345
r34 15 17 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.63 $Y=1.26
+ $X2=3.63 $Y2=0.825
r35 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=1.345
+ $X2=3.63 $Y2=1.26
r36 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=1.345
+ $X2=2.855 $Y2=1.345
r37 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.26
+ $X2=2.855 $Y2=1.345
r38 9 11 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.77 $Y=1.26
+ $X2=2.77 $Y2=0.825
r39 2 17 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.49
+ $Y=0.575 $X2=3.63 $Y2=0.825
r40 1 11 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.63
+ $Y=0.575 $X2=2.77 $Y2=0.825
.ends

