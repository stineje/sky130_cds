* File: sky130_osu_sc_15T_ls__and2_4.pex.spice
* Created: Fri Nov 12 14:53:40 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_LS__AND2_4%GND 1 2 3 37 39 47 49 56 58 66 75 77
r73 75 77 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r74 64 66 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.74
r75 59 71 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r76 58 64 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.305
r77 54 71 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r78 54 56 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.74
r79 49 71 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r80 45 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.305
+ $X2=1.05 $Y2=0.74
r81 37 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r82 37 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r83 37 45 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.05 $Y2=0.305
r84 37 39 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=0.965 $Y2=0.152
r85 37 50 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.152
+ $X2=1.135 $Y2=0.152
r86 37 58 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r87 37 59 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r88 37 49 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r89 37 50 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.135 $Y2=0.152
r90 37 39 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.965 $Y2=0.152
r91 3 66 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.74
r92 2 56 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.74
r93 1 47 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.575 $X2=1.05 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_4%VDD 1 2 3 4 33 37 41 47 51 57 61 68 78
+ 82
r53 78 82 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=2.38 $Y2=5.397
r54 73 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r55 68 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.215
+ $X2=2.84 $Y2=4.575
r56 66 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.575
r57 64 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=5.36
+ $X2=2.38 $Y2=5.36
r58 62 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r59 62 64 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r60 61 66 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.245
r61 61 64 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r62 57 60 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.215
+ $X2=1.98 $Y2=4.575
r63 55 76 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r64 55 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.575
r65 52 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r66 52 54 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r67 51 76 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r68 51 54 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r69 47 50 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.12 $Y=3.555
+ $X2=1.12 $Y2=4.575
r70 45 75 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r71 45 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.575
r72 42 73 3.16604 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=0.172 $Y2=5.397
r73 42 44 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.345 $Y=5.397
+ $X2=1.02 $Y2=5.397
r74 41 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r75 41 44 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r76 37 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.895
+ $X2=0.26 $Y2=4.575
r77 35 73 4.3922 $w=1.7e-07 $l=1.90997e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.172 $Y2=5.397
r78 35 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.26 $Y=5.245
+ $X2=0.26 $Y2=4.575
r79 33 64 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r80 33 54 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r81 33 44 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r82 33 73 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r83 4 71 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.575
r84 4 68 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.215
r85 3 60 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.575
r86 3 57 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.215
r87 2 50 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.575
r88 2 47 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.555
r89 1 40 400 $w=1.7e-07 $l=1.81142e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.575
r90 1 37 400 $w=1.7e-07 $l=1.13077e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.895
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_4%A 3 7 12 15 23
r32 21 23 0.00293427 $w=2.13e-07 $l=5e-09 $layer=MET1_cond $X=0.27 $Y=3.07
+ $X2=0.275 $Y2=3.07
r33 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=3.07
+ $X2=0.27 $Y2=3.07
r34 15 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.27 $Y=2.505
+ $X2=0.27 $Y2=3.07
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.505 $X2=0.27 $Y2=2.505
r36 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.505
+ $X2=0.475 $Y2=2.505
r37 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=2.505
r38 5 7 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=0.475 $Y=2.67
+ $X2=0.475 $Y2=3.825
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=2.505
r40 1 3 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=0.475 $Y=2.34
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_4%B 3 7 10 14 22
c41 7 0 1.37149e-19 $X=0.905 $Y=3.825
r42 20 22 0.00292056 $w=2.14e-07 $l=5e-09 $layer=MET1_cond $X=0.95 $Y=2.7
+ $X2=0.955 $Y2=2.7
r43 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=2.7 $X2=0.95
+ $Y2=2.7
r44 14 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.95 $Y=2.165
+ $X2=0.95 $Y2=2.7
r45 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.165 $X2=0.95 $Y2=2.165
r46 10 12 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2.33
r47 10 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.922 $Y=2.165
+ $X2=0.922 $Y2=2
r48 7 12 766.585 $w=1.5e-07 $l=1.495e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.33
r49 3 11 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.835 $Y=0.945
+ $X2=0.835 $Y2=2
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_4%A_27_115# 1 3 11 13 15 17 18 22 24 26 27
+ 28 29 33 35 37 38 40 44 46 48 49 55 56 57 60 62 63 68 74 76 77 78
c135 33 0 1.33323e-19 $X=2.195 $Y=0.945
c136 22 0 1.33323e-19 $X=1.765 $Y=0.945
r137 77 78 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=3.305
+ $X2=0.65 $Y2=3.475
r138 72 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=0.61 $Y2=1.675
r139 72 74 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.695 $Y=1.675
+ $X2=1.43 $Y2=1.675
r140 68 70 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.69 $Y=3.555
+ $X2=0.69 $Y2=4.575
r141 68 78 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=3.555
+ $X2=0.69 $Y2=3.475
r142 64 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=1.675
r143 64 77 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=3.305
r144 62 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.61 $Y2=1.675
r145 62 63 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=1.675
+ $X2=0.345 $Y2=1.675
r146 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.345 $Y2=1.675
r147 58 60 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.26 $Y=1.59
+ $X2=0.26 $Y2=0.74
r148 53 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.675 $X2=1.43 $Y2=1.675
r149 51 53 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.675
+ $X2=1.43 $Y2=1.675
r150 50 51 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.37 $Y2=1.675
r151 46 48 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r152 42 44 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.625 $Y2=0.945
r153 41 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r154 40 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.7
r155 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r156 39 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.585
+ $X2=2.195 $Y2=1.585
r157 38 42 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.625 $Y2=1.51
r158 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.27 $Y2=1.585
r159 35 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=2.625
r160 35 37 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r161 31 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=1.585
r162 31 33 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=0.945
r163 30 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r164 29 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r165 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r166 27 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=2.195 $Y2=1.585
r167 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=1.84 $Y2=1.585
r168 24 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r169 24 26 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r170 20 28 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.84 $Y2=1.585
r171 20 53 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.43 $Y2=1.675
r172 20 22 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=0.945
r173 19 49 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.625
+ $X2=1.352 $Y2=2.625
r174 18 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r175 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.445 $Y2=2.625
r176 17 49 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.55
+ $X2=1.352 $Y2=2.625
r177 16 51 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=1.675
r178 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=2.55
r179 13 49 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.352 $Y2=2.625
r180 13 15 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r181 9 50 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=1.675
r182 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.945
r183 3 70 300 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=4.575
r184 3 68 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.825 $X2=0.69 $Y2=3.555
r185 1 60 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_OSU_SC_15T_LS__AND2_4%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c78 54 0 1.33323e-19 $X=2.41 $Y=1.335
c79 45 0 1.33323e-19 $X=1.55 $Y=1.335
c80 24 0 1.37149e-19 $X=1.55 $Y=2.33
r81 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.215
+ $X2=2.41 $Y2=2.33
r82 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r83 54 55 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.215
r84 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.33
+ $X2=1.55 $Y2=2.33
r85 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=2.41 $Y2=2.33
r86 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=1.695 $Y2=2.33
r87 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r88 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r89 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r90 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r91 46 48 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r92 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r93 45 48 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r94 41 43 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.215
+ $X2=2.41 $Y2=4.575
r95 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=2.33
r96 38 41 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=3.215
r97 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r98 32 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.41 $Y=0.74
+ $X2=2.41 $Y2=1.22
r99 27 29 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.215
+ $X2=1.55 $Y2=4.575
r100 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r101 24 27 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=3.215
r102 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r103 18 21 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.55 $Y=0.74
+ $X2=1.55 $Y2=1.22
r104 6 43 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.575
r105 6 41 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.215
r106 5 29 240 $w=1.7e-07 $l=1.81865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.575
r107 5 27 240 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.215
r108 2 32 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.74
r109 1 18 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.74
.ends

