* File: sky130_osu_sc_12T_ms__aoi21_l.spice
* Created: Fri Nov 12 15:21:12 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* 
.include "sky130_osu_sc_12T_ms__aoi21_l.pex.spice"
.subckt sky130_osu_sc_12T_ms__aoi21_l  GND VDD A0 A1 B0 Y
* 
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1002 A_110_114# N_A0_M1002_g N_GND_M1002_s N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75000.9 A=0.078 P=1.34 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_110_114# N_GND_M1002_b NSHORT L=0.15 W=0.52
+ AD=0.0964364 AS=0.0546 PD=1.01636 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75000.5 A=0.078 P=1.34 MULT=1
MM1003 N_GND_M1003_d N_B0_M1003_g N_Y_M1001_d N_GND_M1002_b NSHORT L=0.15 W=0.36
+ AD=0.0954 AS=0.0667636 PD=1.25 PS=0.703636 NRD=0 NRS=19.992 M=1 R=2.4 SA=75001
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1000 N_VDD_M1000_d N_A0_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_A_27_521#_M1004_d N_A1_M1004_g N_VDD_M1000_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_B0_M1005_g N_A_27_521#_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1000_b NWDIODE A=3.9552 P=7.96
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_ms__aoi21_l.pxi.spice"
*
.ends
*
*
