* File: sky130_osu_sc_15T_ms__or2_4.pex.spice
* Created: Fri Nov 12 14:46:09 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_15T_MS__OR2_4%GND 1 2 3 4 41 45 47 54 56 63 65 73 84 86
r72 84 86 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=2.38 $Y2=0.152
r73 71 73 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.84 $Y=0.305
+ $X2=2.84 $Y2=0.865
r74 66 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.152
+ $X2=1.98 $Y2=0.152
r75 65 71 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.755 $Y=0.152
+ $X2=2.84 $Y2=0.305
r76 61 80 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.152
r77 61 63 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.98 $Y=0.305
+ $X2=1.98 $Y2=0.865
r78 57 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.152
+ $X2=1.12 $Y2=0.152
r79 56 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.152
+ $X2=1.98 $Y2=0.152
r80 52 79 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.152
r81 52 54 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0.305
+ $X2=1.12 $Y2=0.865
r82 47 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0.152
+ $X2=1.12 $Y2=0.152
r83 43 45 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.26 $Y=0.305
+ $X2=0.26 $Y2=0.865
r84 41 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=0.19
+ $X2=2.38 $Y2=0.19
r85 41 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=0.19
+ $X2=0.34 $Y2=0.19
r86 41 43 4.39984 $w=1.7e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.26 $Y2=0.305
r87 41 48 3.15839 $w=3.05e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0.152
+ $X2=0.345 $Y2=0.152
r88 41 65 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.755 $Y2=0.152
r89 41 66 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.38 $Y=0.152
+ $X2=2.065 $Y2=0.152
r90 41 56 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.895 $Y2=0.152
r91 41 57 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.205 $Y2=0.152
r92 41 47 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.035 $Y2=0.152
r93 41 48 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.345 $Y2=0.152
r94 4 73 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.865
r95 3 63 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.865
r96 2 54 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.865
r97 1 45 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_4%VDD 1 2 3 29 31 40 44 50 54 61 68 72
r47 68 72 0.950071 $w=3.05e-07 $l=2.04e-06 $layer=MET1_cond $X=0.34 $Y=5.397
+ $X2=2.38 $Y2=5.397
r48 61 64 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.84 $Y=3.205
+ $X2=2.84 $Y2=4.565
r49 59 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.84 $Y=5.245
+ $X2=2.84 $Y2=4.565
r50 57 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.38 $Y=5.36
+ $X2=2.38 $Y2=5.36
r51 55 66 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=1.98 $Y2=5.397
r52 55 57 11.9023 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=5.397
+ $X2=2.38 $Y2=5.397
r53 54 59 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.84 $Y2=5.245
r54 54 57 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.755 $Y=5.397
+ $X2=2.38 $Y2=5.397
r55 50 53 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.98 $Y=3.205
+ $X2=1.98 $Y2=4.565
r56 48 66 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=5.397
r57 48 53 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.98 $Y=5.245
+ $X2=1.98 $Y2=4.565
r58 45 65 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.12 $Y2=5.397
r59 45 47 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=5.397
+ $X2=1.7 $Y2=5.397
r60 44 66 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.98 $Y2=5.397
r61 44 47 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.895 $Y=5.397
+ $X2=1.7 $Y2=5.397
r62 40 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=3.885
+ $X2=1.12 $Y2=4.565
r63 38 65 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=5.397
r64 38 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=5.245
+ $X2=1.12 $Y2=4.565
r65 33 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.34 $Y=5.36
+ $X2=0.34 $Y2=5.36
r66 33 37 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.34 $Y=5.397
+ $X2=1.02 $Y2=5.397
r67 31 65 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.12 $Y2=5.397
r68 31 37 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=5.397
+ $X2=1.02 $Y2=5.397
r69 29 57 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=5.245 $X2=2.38 $Y2=5.33
r70 29 47 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=5.245 $X2=1.7 $Y2=5.33
r71 29 37 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=5.245 $X2=1.02 $Y2=5.33
r72 29 33 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=5.245 $X2=0.34 $Y2=5.33
r73 3 64 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=4.565
r74 3 61 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=2.825 $X2=2.84 $Y2=3.205
r75 2 53 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=4.565
r76 2 50 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.825 $X2=1.98 $Y2=3.205
r77 1 43 400 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=4.565
r78 1 40 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.825 $X2=1.12 $Y2=3.885
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_4%B 3 7 12 15 21
r28 18 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.27 $Y=2.7 $X2=0.27
+ $Y2=2.7
r29 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.27 $Y=2.415
+ $X2=0.27 $Y2=2.7
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=2.415 $X2=0.27 $Y2=2.415
r31 10 12 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=2.415
+ $X2=0.475 $Y2=2.415
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.58
+ $X2=0.475 $Y2=2.415
r33 5 7 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=0.475 $Y=2.58
+ $X2=0.475 $Y2=3.825
r34 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.25
+ $X2=0.475 $Y2=2.415
r35 1 3 669.16 $w=1.5e-07 $l=1.305e-06 $layer=POLY_cond $X=0.475 $Y=2.25
+ $X2=0.475 $Y2=0.945
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_4%A 3 7 10 14 20
c44 7 0 1.37149e-19 $X=0.905 $Y=3.825
r45 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.95 $Y=3.07
+ $X2=0.95 $Y2=3.07
r46 14 17 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.95 $Y=2.125
+ $X2=0.95 $Y2=3.07
r47 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.125 $X2=0.95 $Y2=2.125
r48 10 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.125
+ $X2=0.95 $Y2=2.29
r49 10 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.125
+ $X2=0.95 $Y2=1.96
r50 7 12 787.096 $w=1.5e-07 $l=1.535e-06 $layer=POLY_cond $X=0.905 $Y=3.825
+ $X2=0.905 $Y2=2.29
r51 3 11 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=0.905 $Y=0.945
+ $X2=0.905 $Y2=1.96
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_4%A_27_565# 1 3 11 13 15 17 18 22 24 26 27
+ 28 29 33 35 37 38 40 44 46 48 49 55 56 57 60 64 65 67 70 74 76
c135 33 0 1.33323e-19 $X=2.195 $Y=0.945
c136 22 0 1.33323e-19 $X=1.765 $Y=0.945
r137 72 76 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.775 $Y=1.675
+ $X2=0.65 $Y2=1.675
r138 72 74 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.775 $Y=1.675
+ $X2=1.43 $Y2=1.675
r139 68 76 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.65 $Y2=1.675
r140 68 70 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.69 $Y=1.59
+ $X2=0.69 $Y2=0.865
r141 66 76 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.65 $Y2=1.675
r142 66 67 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=0.61 $Y=1.76
+ $X2=0.61 $Y2=3.285
r143 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.525 $Y=3.37
+ $X2=0.61 $Y2=3.285
r144 64 65 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.525 $Y=3.37
+ $X2=0.345 $Y2=3.37
r145 60 62 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.26 $Y=3.545
+ $X2=0.26 $Y2=4.565
r146 58 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.345 $Y2=3.37
r147 58 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=3.545
r148 53 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.675 $X2=1.43 $Y2=1.675
r149 51 53 12.412 $w=2.33e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.675
+ $X2=1.43 $Y2=1.675
r150 50 51 7.24034 $w=2.33e-07 $l=3.5e-08 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.37 $Y2=1.675
r151 46 48 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.625 $Y=2.7
+ $X2=2.625 $Y2=3.825
r152 42 44 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.625 $Y2=0.945
r153 41 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.625
+ $X2=2.195 $Y2=2.625
r154 40 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.625 $Y2=2.7
r155 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.625
+ $X2=2.27 $Y2=2.625
r156 39 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.585
+ $X2=2.195 $Y2=1.585
r157 38 42 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.625 $Y2=1.51
r158 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.585
+ $X2=2.27 $Y2=1.585
r159 35 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=2.625
r160 35 37 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.195 $Y=2.7
+ $X2=2.195 $Y2=3.825
r161 31 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=1.585
r162 31 33 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.195 $Y2=0.945
r163 30 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.625
+ $X2=1.765 $Y2=2.625
r164 29 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=2.195 $Y2=2.625
r165 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.625
+ $X2=1.84 $Y2=2.625
r166 27 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=2.195 $Y2=1.585
r167 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.585
+ $X2=1.84 $Y2=1.585
r168 24 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=2.625
r169 24 26 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.765 $Y=2.7
+ $X2=1.765 $Y2=3.825
r170 20 28 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.84 $Y2=1.585
r171 20 53 69.3004 $w=2.33e-07 $l=4.09268e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.43 $Y2=1.675
r172 20 22 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.765 $Y2=0.945
r173 19 49 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.445 $Y=2.625
+ $X2=1.352 $Y2=2.625
r174 18 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.765 $Y2=2.625
r175 18 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.69 $Y=2.625
+ $X2=1.445 $Y2=2.625
r176 17 49 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=1.37 $Y=2.55
+ $X2=1.352 $Y2=2.625
r177 16 51 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=1.675
r178 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.37 $Y=1.84
+ $X2=1.37 $Y2=2.55
r179 13 49 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.352 $Y2=2.625
r180 13 15 361.5 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.335 $Y=2.7
+ $X2=1.335 $Y2=3.825
r181 9 50 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=1.675
r182 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=0.945
r183 3 62 300 $w=1.7e-07 $l=1.80142e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=4.565
r184 3 60 300 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.825 $X2=0.26 $Y2=3.545
r185 1 70 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_OSU_SC_15T_MS__OR2_4%Y 1 2 5 6 18 24 32 38 45 46 48 50 52 54
+ 55
c77 54 0 1.33323e-19 $X=2.41 $Y=1.335
c78 45 0 1.33323e-19 $X=1.55 $Y=1.335
c79 24 0 1.37149e-19 $X=1.55 $Y=2.33
r80 55 63 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=2.215
+ $X2=2.41 $Y2=2.33
r81 54 61 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=1.22
r82 54 55 0.847336 $w=1.7e-07 $l=8.8e-07 $layer=MET1_cond $X=2.41 $Y=1.335
+ $X2=2.41 $Y2=2.215
r83 53 59 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=2.33
+ $X2=1.55 $Y2=2.33
r84 52 63 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=2.41 $Y2=2.33
r85 52 53 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=2.33
+ $X2=1.695 $Y2=2.33
r86 51 57 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.695 $Y=1.22
+ $X2=1.55 $Y2=1.22
r87 50 61 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=2.41 $Y2=1.22
r88 50 51 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.265 $Y=1.22
+ $X2=1.695 $Y2=1.22
r89 46 59 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=2.33
r90 46 48 0.245535 $w=1.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.55 $Y=2.215
+ $X2=1.55 $Y2=1.96
r91 45 57 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.22
r92 45 48 0.601801 $w=1.7e-07 $l=6.25e-07 $layer=MET1_cond $X=1.55 $Y=1.335
+ $X2=1.55 $Y2=1.96
r93 41 43 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.41 $Y=3.205
+ $X2=2.41 $Y2=4.565
r94 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=2.33
r95 38 41 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.41 $Y=2.33
+ $X2=2.41 $Y2=3.205
r96 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.41 $Y=1.22
+ $X2=2.41 $Y2=1.22
r97 32 35 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.41 $Y=0.865
+ $X2=2.41 $Y2=1.22
r98 27 29 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.55 $Y=3.205
+ $X2=1.55 $Y2=4.565
r99 24 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=2.33
r100 24 27 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.55 $Y=2.33
+ $X2=1.55 $Y2=3.205
r101 21 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.55 $Y=1.22
+ $X2=1.55 $Y2=1.22
r102 18 21 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.55 $Y=0.865
+ $X2=1.55 $Y2=1.22
r103 6 43 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=4.565
r104 6 41 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.825 $X2=2.41 $Y2=3.205
r105 5 29 240 $w=1.7e-07 $l=1.80865e-06 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=4.565
r106 5 27 240 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.825 $X2=1.55 $Y2=3.205
r107 2 32 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.865
r108 1 18 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.865
.ends

