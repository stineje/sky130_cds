magic
tech sky130A
magscale 1 2
timestamp 1646761263
<< checkpaint >>
rect -1529 2461 2577 2602
rect -1760 -1129 6260 2461
rect -1529 -1260 2577 -1129
<< nwell >>
rect 0 1089 255 1090
rect -269 529 1317 1089
<< nmoslvt >>
rect -180 115 -150 263
rect -94 115 -64 263
rect 96 115 126 263
rect 182 115 212 263
rect 254 115 284 263
rect 374 115 404 263
rect 446 115 476 263
rect 532 115 562 263
rect 740 115 770 263
rect 826 115 856 263
rect 1016 115 1046 263
rect 1088 115 1118 263
rect 1188 115 1218 263
<< pmos >>
rect -180 565 -150 965
rect -108 565 -78 965
rect 96 565 126 965
rect 182 565 212 965
rect 254 565 284 965
rect 374 565 404 965
rect 446 565 476 965
rect 532 565 562 965
rect 740 565 770 965
rect 826 565 856 965
rect 1016 565 1046 965
rect 1102 565 1132 965
rect 1188 565 1218 965
<< ndiff >>
rect -233 215 -180 263
rect -233 131 -225 215
rect -191 131 -180 215
rect -233 115 -180 131
rect -150 215 -94 263
rect -150 131 -139 215
rect -105 131 -94 215
rect -150 115 -94 131
rect -64 215 -11 263
rect -64 131 -53 215
rect -19 131 -11 215
rect -64 115 -11 131
rect 43 215 96 263
rect 43 131 51 215
rect 85 131 96 215
rect 43 115 96 131
rect 126 215 182 263
rect 126 131 137 215
rect 171 131 182 215
rect 126 115 182 131
rect 212 115 254 263
rect 284 215 374 263
rect 284 131 295 215
rect 363 131 374 215
rect 284 115 374 131
rect 404 115 446 263
rect 476 215 532 263
rect 476 131 487 215
rect 521 131 532 215
rect 476 115 532 131
rect 562 215 615 263
rect 562 131 573 215
rect 607 131 615 215
rect 562 115 615 131
rect 687 215 740 263
rect 687 131 695 215
rect 729 131 740 215
rect 687 115 740 131
rect 770 215 826 263
rect 770 131 781 215
rect 815 131 826 215
rect 770 115 826 131
rect 856 215 909 263
rect 856 131 867 215
rect 901 131 909 215
rect 856 115 909 131
rect 963 215 1016 263
rect 963 131 971 215
rect 1005 131 1016 215
rect 963 115 1016 131
rect 1046 115 1088 263
rect 1118 215 1188 263
rect 1118 131 1129 215
rect 1163 131 1188 215
rect 1118 115 1188 131
rect 1218 215 1271 263
rect 1218 131 1229 215
rect 1263 131 1271 215
rect 1218 115 1271 131
<< pdiff >>
rect -233 949 -180 965
rect -233 605 -225 949
rect -191 605 -180 949
rect -233 565 -180 605
rect -150 565 -108 965
rect -78 949 -25 965
rect -78 741 -67 949
rect -33 741 -25 949
rect -78 565 -25 741
rect 43 949 96 965
rect 43 673 51 949
rect 85 673 96 949
rect 43 565 96 673
rect 126 949 182 965
rect 126 673 137 949
rect 171 673 182 949
rect 126 565 182 673
rect 212 565 254 965
rect 284 949 374 965
rect 284 605 295 949
rect 363 605 374 949
rect 284 565 374 605
rect 404 565 446 965
rect 476 949 532 965
rect 476 605 487 949
rect 521 605 532 949
rect 476 565 532 605
rect 562 949 615 965
rect 562 605 573 949
rect 607 605 615 949
rect 562 565 615 605
rect 687 949 740 965
rect 687 605 695 949
rect 729 605 740 949
rect 687 565 740 605
rect 770 949 826 965
rect 770 605 781 949
rect 815 605 826 949
rect 770 565 826 605
rect 856 949 909 965
rect 856 605 867 949
rect 901 605 909 949
rect 856 565 909 605
rect 963 949 1016 965
rect 963 741 971 949
rect 1005 741 1016 949
rect 963 565 1016 741
rect 1046 949 1102 965
rect 1046 673 1057 949
rect 1091 673 1102 949
rect 1046 565 1102 673
rect 1132 949 1188 965
rect 1132 673 1143 949
rect 1177 673 1188 949
rect 1132 565 1188 673
rect 1218 949 1271 965
rect 1218 605 1229 949
rect 1263 605 1271 949
rect 1218 565 1271 605
<< ndiffc >>
rect -225 131 -191 215
rect -139 131 -105 215
rect -53 131 -19 215
rect 51 131 85 215
rect 137 131 171 215
rect 295 131 363 215
rect 487 131 521 215
rect 573 131 607 215
rect 695 131 729 215
rect 781 131 815 215
rect 867 131 901 215
rect 971 131 1005 215
rect 1129 131 1163 215
rect 1229 131 1263 215
<< pdiffc >>
rect -225 605 -191 949
rect -67 741 -33 949
rect 51 673 85 949
rect 137 673 171 949
rect 295 605 363 949
rect 487 605 521 949
rect 573 605 607 949
rect 695 605 729 949
rect 781 605 815 949
rect 867 605 901 949
rect 971 741 1005 949
rect 1057 673 1091 949
rect 1143 673 1177 949
rect 1229 605 1263 949
<< psubdiff >>
rect -233 27 -209 61
rect -175 27 -151 61
rect -97 27 -73 61
rect -39 27 -15 61
rect 88 27 112 61
rect 146 27 170 61
rect 224 27 248 61
rect 282 27 306 61
rect 360 27 384 61
rect 418 27 442 61
rect 496 27 520 61
rect 554 27 578 61
rect 632 27 656 61
rect 690 27 714 61
rect 768 27 792 61
rect 826 27 850 61
rect 963 27 987 61
rect 1021 27 1045 61
rect 1099 27 1123 61
rect 1157 27 1181 61
<< nsubdiff >>
rect -233 1019 -209 1053
rect -175 1019 -151 1053
rect -97 1019 -73 1053
rect -39 1019 -15 1053
rect 88 1019 112 1053
rect 146 1019 170 1053
rect 224 1019 248 1053
rect 282 1019 306 1053
rect 360 1019 384 1053
rect 418 1019 442 1053
rect 496 1019 520 1053
rect 554 1019 578 1053
rect 632 1019 656 1053
rect 690 1019 714 1053
rect 768 1019 792 1053
rect 826 1019 850 1053
rect 963 1019 987 1053
rect 1021 1019 1045 1053
rect 1099 1019 1123 1053
rect 1157 1019 1181 1053
<< psubdiffcont >>
rect -209 27 -175 61
rect -73 27 -39 61
rect 112 27 146 61
rect 248 27 282 61
rect 384 27 418 61
rect 520 27 554 61
rect 656 27 690 61
rect 792 27 826 61
rect 987 27 1021 61
rect 1123 27 1157 61
<< nsubdiffcont >>
rect -209 1019 -175 1053
rect -73 1019 -39 1053
rect 112 1019 146 1053
rect 248 1019 282 1053
rect 384 1019 418 1053
rect 520 1019 554 1053
rect 656 1019 690 1053
rect 792 1019 826 1053
rect 987 1019 1021 1053
rect 1123 1019 1157 1053
<< poly >>
rect -180 965 -150 991
rect -108 965 -78 991
rect 96 965 126 991
rect 182 965 212 991
rect 254 965 284 991
rect 374 965 404 991
rect 446 965 476 991
rect 532 965 562 991
rect 740 965 770 991
rect 826 965 856 991
rect 1016 965 1046 991
rect 1102 965 1132 991
rect 1188 965 1218 991
rect -180 399 -150 565
rect -108 532 -78 565
rect 96 543 126 565
rect -108 516 -35 532
rect -108 482 -79 516
rect -45 482 -35 516
rect -108 466 -35 482
rect 86 509 126 543
rect -204 383 -150 399
rect -204 349 -194 383
rect -160 349 -150 383
rect -204 333 -150 349
rect -180 263 -150 333
rect -94 263 -64 466
rect 86 351 116 509
rect 182 466 212 565
rect 254 534 284 565
rect 374 534 404 565
rect 254 518 308 534
rect 254 484 264 518
rect 298 484 308 518
rect 254 468 308 484
rect 350 518 404 534
rect 350 484 360 518
rect 394 484 404 518
rect 350 468 404 484
rect 158 450 212 466
rect 158 416 168 450
rect 202 416 212 450
rect 350 423 380 468
rect 158 400 212 416
rect 86 335 140 351
rect 86 301 96 335
rect 130 301 140 335
rect 86 285 140 301
rect 96 263 126 285
rect 182 263 212 400
rect 254 393 380 423
rect 446 425 476 565
rect 532 535 562 565
rect 740 549 770 565
rect 532 504 573 535
rect 446 409 500 425
rect 254 263 284 393
rect 446 375 456 409
rect 490 375 500 409
rect 446 359 500 375
rect 350 335 404 351
rect 350 301 360 335
rect 394 301 404 335
rect 350 285 404 301
rect 374 263 404 285
rect 446 263 476 359
rect 543 351 573 504
rect 730 519 770 549
rect 730 425 760 519
rect 826 425 856 565
rect 1016 534 1046 565
rect 963 518 1046 534
rect 963 484 973 518
rect 1007 484 1046 518
rect 963 468 1046 484
rect 705 409 760 425
rect 705 375 715 409
rect 749 375 760 409
rect 705 359 760 375
rect 802 409 856 425
rect 802 375 812 409
rect 846 375 856 409
rect 802 359 856 375
rect 543 335 601 351
rect 543 311 557 335
rect 532 301 557 311
rect 591 301 601 335
rect 532 281 601 301
rect 730 308 760 359
rect 532 263 562 281
rect 730 278 770 308
rect 740 263 770 278
rect 826 263 856 359
rect 1016 263 1046 468
rect 1102 466 1132 565
rect 1188 540 1218 565
rect 1188 510 1225 540
rect 1088 450 1153 466
rect 1088 416 1109 450
rect 1143 416 1153 450
rect 1088 400 1153 416
rect 1088 263 1118 400
rect 1195 368 1225 510
rect 1195 352 1249 368
rect 1195 332 1205 352
rect 1188 318 1205 332
rect 1239 318 1249 352
rect 1188 302 1249 318
rect 1188 263 1218 302
rect -180 89 -150 115
rect -94 89 -64 115
rect 96 89 126 115
rect 182 89 212 115
rect 254 89 284 115
rect 374 89 404 115
rect 446 89 476 115
rect 532 89 562 115
rect 740 89 770 115
rect 826 89 856 115
rect 1016 89 1046 115
rect 1088 89 1118 115
rect 1188 89 1218 115
<< polycont >>
rect -79 482 -45 516
rect -194 349 -160 383
rect 264 484 298 518
rect 360 484 394 518
rect 168 416 202 450
rect 96 301 130 335
rect 456 375 490 409
rect 360 301 394 335
rect 973 484 1007 518
rect 715 375 749 409
rect 812 375 846 409
rect 557 301 591 335
rect 1109 416 1143 450
rect 1205 318 1239 352
<< locali >>
rect -267 1059 1317 1080
rect -267 1019 -209 1059
rect -175 1019 -73 1059
rect -39 1019 112 1059
rect 146 1019 248 1059
rect 282 1019 384 1059
rect 418 1019 520 1059
rect 554 1019 656 1059
rect 690 1019 792 1059
rect 826 1019 987 1059
rect 1021 1019 1123 1059
rect 1157 1019 1317 1059
rect -225 949 -191 965
rect -67 949 -33 1019
rect -67 725 -33 741
rect 51 949 85 965
rect 28 673 51 739
rect 28 656 85 673
rect 137 949 171 1019
rect 137 657 171 673
rect 295 949 363 965
rect -225 483 -191 605
rect -147 383 -113 523
rect -79 516 -45 597
rect -79 466 -45 482
rect -210 349 -194 383
rect -160 349 -113 383
rect 28 409 62 656
rect 295 602 363 605
rect -225 215 -191 231
rect -225 61 -191 131
rect 28 244 62 375
rect 96 568 363 602
rect 487 949 521 1019
rect 487 589 521 605
rect 573 949 607 965
rect 96 335 130 568
rect 360 518 394 534
rect 248 484 264 518
rect 298 484 314 518
rect 168 400 202 416
rect 280 335 314 484
rect 360 483 394 484
rect 573 483 607 605
rect 695 949 729 965
rect 695 518 729 597
rect 781 949 815 1019
rect 781 589 815 605
rect 867 949 901 965
rect 971 949 1005 1019
rect 971 725 1005 741
rect 1057 949 1091 965
rect 1041 673 1057 691
rect 1041 657 1091 673
rect 1143 949 1177 1019
rect 1143 657 1177 673
rect 1229 949 1263 965
rect 901 605 914 614
rect 867 580 914 605
rect 695 484 846 518
rect 573 419 607 449
rect 440 375 456 409
rect 490 375 506 409
rect 573 385 661 419
rect 812 409 846 484
rect 557 335 591 351
rect 130 301 239 335
rect 280 301 360 335
rect 394 301 557 335
rect 96 285 130 301
rect 205 251 239 301
rect 557 285 591 301
rect 627 251 661 385
rect 699 375 715 409
rect 749 375 765 409
rect 812 335 846 375
rect -139 215 -105 227
rect -139 115 -105 131
rect -53 215 -19 231
rect 28 215 85 244
rect 28 210 51 215
rect -53 61 -19 131
rect 51 115 85 131
rect 137 215 171 231
rect 205 217 363 251
rect 137 61 171 131
rect 295 215 363 217
rect 295 115 363 131
rect 487 215 521 231
rect 487 61 521 131
rect 573 217 661 251
rect 695 301 846 335
rect 880 335 914 580
rect 973 518 1007 597
rect 973 468 1007 484
rect 1041 352 1075 657
rect 1109 450 1143 523
rect 1229 483 1263 605
rect 1109 400 1143 416
rect 1205 352 1239 368
rect 573 215 607 217
rect 573 115 607 131
rect 695 215 729 301
rect 880 267 914 301
rect 867 233 914 267
rect 971 318 1205 352
rect 695 115 729 131
rect 781 215 815 231
rect 781 61 815 131
rect 867 215 901 233
rect 867 115 901 131
rect 971 215 1005 318
rect 1205 302 1239 318
rect 971 115 1005 131
rect 1129 215 1163 231
rect 1129 61 1163 131
rect 1229 215 1263 227
rect 1229 115 1263 131
rect -267 21 -209 61
rect -175 21 -73 61
rect -39 21 112 61
rect 146 21 248 61
rect 282 21 384 61
rect 418 21 520 61
rect 554 21 656 61
rect 690 21 792 61
rect 826 21 987 61
rect 1021 21 1123 61
rect 1157 21 1317 61
rect -267 0 1317 21
<< viali >>
rect -209 1053 -175 1059
rect -209 1025 -175 1053
rect -73 1053 -39 1059
rect -73 1025 -39 1053
rect 112 1053 146 1059
rect 112 1025 146 1053
rect 248 1053 282 1059
rect 248 1025 282 1053
rect 384 1053 418 1059
rect 384 1025 418 1053
rect 520 1053 554 1059
rect 520 1025 554 1053
rect 656 1053 690 1059
rect 656 1025 690 1053
rect 792 1053 826 1059
rect 792 1025 826 1053
rect 987 1053 1021 1059
rect 987 1025 1021 1053
rect 1123 1053 1157 1059
rect 1123 1025 1157 1053
rect -79 597 -45 631
rect -225 449 -191 483
rect -147 523 -113 557
rect 28 375 62 409
rect -139 227 -105 261
rect 264 484 298 518
rect 168 450 202 484
rect 360 449 394 483
rect 695 605 729 631
rect 695 597 729 605
rect 573 449 607 483
rect 456 375 490 409
rect 557 301 591 335
rect 715 375 749 409
rect 973 597 1007 631
rect 1109 523 1143 557
rect 1229 449 1263 483
rect 880 301 914 335
rect 1229 227 1263 261
rect -209 27 -175 55
rect -209 21 -175 27
rect -73 27 -39 55
rect -73 21 -39 27
rect 112 27 146 55
rect 112 21 146 27
rect 248 27 282 55
rect 248 21 282 27
rect 384 27 418 55
rect 384 21 418 27
rect 520 27 554 55
rect 520 21 554 27
rect 656 27 690 55
rect 656 21 690 27
rect 792 27 826 55
rect 792 21 826 27
rect 987 27 1021 55
rect 987 21 1021 27
rect 1123 27 1157 55
rect 1123 21 1157 27
<< metal1 >>
rect -267 1059 1317 1080
rect -267 1025 -209 1059
rect -175 1025 -73 1059
rect -39 1025 112 1059
rect 146 1025 248 1059
rect 282 1025 384 1059
rect 418 1025 520 1059
rect 554 1025 656 1059
rect 690 1025 792 1059
rect 826 1025 987 1059
rect 1021 1025 1123 1059
rect 1157 1025 1317 1059
rect -267 1019 1317 1025
rect -91 631 -33 637
rect -112 597 -79 631
rect -45 597 -33 631
rect -91 591 -33 597
rect 682 631 740 637
rect 961 631 1019 637
rect 682 597 695 631
rect 729 597 973 631
rect 1007 597 1041 631
rect 682 591 740 597
rect 961 591 1019 597
rect -159 557 -101 563
rect 1097 557 1155 563
rect -181 523 -147 557
rect -113 523 -101 557
rect 264 524 314 557
rect -159 517 -101 523
rect 252 523 314 524
rect 1077 523 1109 557
rect 1143 523 1155 557
rect 252 518 310 523
rect -237 483 -179 489
rect 156 484 215 490
rect -142 483 168 484
rect -237 449 -225 483
rect -191 450 168 483
rect 202 450 215 484
rect 252 484 264 518
rect 298 484 310 518
rect 1097 517 1155 523
rect 252 478 310 484
rect 348 483 406 489
rect 561 483 619 489
rect -191 449 215 450
rect -237 443 -179 449
rect -139 267 -105 449
rect 156 444 215 449
rect 348 449 360 483
rect 394 449 573 483
rect 607 449 619 483
rect 348 443 406 449
rect 561 443 619 449
rect 1217 483 1275 489
rect 1217 449 1229 483
rect 1263 449 1275 483
rect 1217 443 1275 449
rect 15 409 74 415
rect 15 375 28 409
rect 62 402 74 409
rect 444 409 503 415
rect 444 402 456 409
rect 62 375 456 402
rect 490 406 503 409
rect 703 409 761 415
rect 703 406 715 409
rect 490 378 715 406
rect 490 375 503 378
rect 15 374 503 375
rect 15 369 74 374
rect 444 369 503 374
rect 703 375 715 378
rect 749 375 761 409
rect 703 369 761 375
rect 543 335 603 341
rect 521 301 557 335
rect 591 301 603 335
rect 543 295 603 301
rect 867 335 927 344
rect 867 301 880 335
rect 914 301 942 335
rect 867 300 942 301
rect 867 292 927 300
rect 1229 267 1263 443
rect -151 261 -93 267
rect -151 227 -139 261
rect -105 227 -93 261
rect -151 221 -93 227
rect 1217 261 1275 267
rect 1217 227 1229 261
rect 1263 227 1275 261
rect 1217 221 1275 227
rect -267 55 1317 61
rect -267 21 -209 55
rect -175 21 -73 55
rect -39 21 112 55
rect 146 21 248 55
rect 282 21 384 55
rect 418 21 520 55
rect 554 21 656 55
rect 690 21 792 55
rect 826 21 987 55
rect 1021 21 1123 55
rect 1157 21 1317 55
rect -267 0 1317 21
<< labels >>
rlabel viali -131 540 -131 540 1 SE
port 1 n
rlabel viali -62 615 -62 615 1 E
port 2 n
rlabel viali 574 318 574 318 1 CK
port 3 n
rlabel metal1 1245 391 1245 391 1 ECK
port 4 n
rlabel metal1 895 314 895 318 1 Q
port 5 n
rlabel viali 1126 541 1126 541 1 CKa
port 6 n
rlabel viali -192 1038 -192 1038 1 vdd
rlabel viali -55 1039 -55 1039 1 vdd
rlabel viali 129 1040 129 1040 1 vdd
rlabel viali 265 1040 265 1040 1 vdd
rlabel viali 401 1040 401 1040 1 vdd
rlabel viali 538 1042 538 1042 1 vdd
rlabel viali 673 1041 673 1041 1 vdd
rlabel viali 809 1040 809 1040 1 vdd
rlabel viali 1005 1041 1005 1041 1 vdd
rlabel viali 1141 1041 1141 1041 1 vdd
rlabel viali -192 44 -192 44 1 gnd
rlabel viali -56 44 -56 44 1 gnd
rlabel viali 129 44 129 44 1 gnd
rlabel viali 264 42 264 42 1 gnd
rlabel viali 401 39 401 39 1 gnd
rlabel viali 537 39 537 39 1 gnd
rlabel viali 673 40 673 40 1 gnd
rlabel viali 809 40 809 40 1 gnd
rlabel viali 1004 40 1004 40 1 gnd
rlabel viali 1140 40 1140 40 1 gnd
<< end >>
