* File: sky130_osu_sc_18T_ls__buf_8.pex.spice
* Created: Thu Oct 29 17:35:07 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_OSU_SC_18T_LS__BUF_8%GND 1 2 3 4 5 40 44 46 53 55 62 64 71 75
+ 77 85 90 92
r119 90 92 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=0.152
+ $X2=3.74 $Y2=0.152
r120 83 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.152
+ $X2=3.27 $Y2=0.152
r121 77 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.152
+ $X2=0.69 $Y2=0.152
r122 73 85 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=4.13 $Y=0.305
+ $X2=4.045 $Y2=0.152
r123 73 75 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.13 $Y=0.305
+ $X2=4.13 $Y2=0.825
r124 69 84 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.152
r125 69 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=0.305
+ $X2=3.27 $Y2=0.825
r126 64 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.152
+ $X2=3.27 $Y2=0.152
r127 60 62 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=0.305
+ $X2=2.41 $Y2=0.825
r128 56 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0.152
+ $X2=1.55 $Y2=0.152
r129 51 79 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.152
r130 51 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=0.305
+ $X2=1.55 $Y2=0.825
r131 47 78 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.152
+ $X2=0.69 $Y2=0.152
r132 46 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0.152
+ $X2=1.55 $Y2=0.152
r133 42 78 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.152
r134 42 44 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=0.305
+ $X2=0.69 $Y2=0.825
r135 40 85 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=4.045 $Y2=0.152
r136 40 83 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=3.74 $Y=0.152
+ $X2=3.355 $Y2=0.152
r137 40 77 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.34 $Y=0.152
+ $X2=0.605 $Y2=0.152
r138 40 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=0.17
+ $X2=3.74 $Y2=0.17
r139 40 90 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=0.17
+ $X2=0.34 $Y2=0.17
r140 40 60 3.51065 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.41 $Y2=0.305
r141 40 55 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.325 $Y2=0.152
r142 40 65 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.152
+ $X2=2.495 $Y2=0.152
r143 40 64 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=3.185 $Y2=0.152
r144 40 65 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=3.06 $Y=0.152
+ $X2=2.495 $Y2=0.152
r145 40 55 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=2.325 $Y2=0.152
r146 40 56 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.7 $Y=0.152
+ $X2=1.635 $Y2=0.152
r147 40 46 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=1.465 $Y2=0.152
r148 40 47 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=0.152
+ $X2=0.775 $Y2=0.152
r149 5 75 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.575 $X2=4.13 $Y2=0.825
r150 4 71 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.575 $X2=3.27 $Y2=0.825
r151 3 62 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.575 $X2=2.41 $Y2=0.825
r152 2 53 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.575 $X2=1.55 $Y2=0.825
r153 1 44 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.575 $X2=0.69 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_8%VDD 1 2 3 4 5 34 38 42 48 52 58 62 68 74
+ 78 85 87 92
r82 92 99 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.74 $Y=6.49
+ $X2=3.74 $Y2=6.49
r83 87 92 1.58345 $w=3.05e-07 $l=3.4e-06 $layer=MET1_cond $X=0.34 $Y=6.507
+ $X2=3.74 $Y2=6.507
r84 87 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.34 $Y=6.49
+ $X2=0.34 $Y2=6.49
r85 85 99 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.045 $Y=6.507
+ $X2=3.74 $Y2=6.507
r86 83 99 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=3.355 $Y=6.507
+ $X2=3.74 $Y2=6.507
r87 83 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=6.507
+ $X2=3.27 $Y2=6.507
r88 78 96 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.34 $Y2=6.507
r89 78 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=6.507
+ $X2=0.69 $Y2=6.507
r90 74 77 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.13 $Y=3.455
+ $X2=4.13 $Y2=5.835
r91 72 85 7.55824 $w=3.05e-07 $l=1.898e-07 $layer=LI1_cond $X=4.13 $Y=6.355
+ $X2=4.045 $Y2=6.507
r92 72 77 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.13 $Y=6.355
+ $X2=4.13 $Y2=5.835
r93 68 71 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.27 $Y=3.455
+ $X2=3.27 $Y2=5.835
r94 66 84 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.27 $Y=6.355
+ $X2=3.27 $Y2=6.507
r95 66 71 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.27 $Y=6.355
+ $X2=3.27 $Y2=5.835
r96 63 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=2.41 $Y2=6.507
r97 63 65 21.3485 $w=3.03e-07 $l=5.65e-07 $layer=LI1_cond $X=2.495 $Y=6.507
+ $X2=3.06 $Y2=6.507
r98 62 84 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.27 $Y2=6.507
r99 62 65 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=6.507
+ $X2=3.06 $Y2=6.507
r100 58 61 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.41 $Y=3.455
+ $X2=2.41 $Y2=5.835
r101 56 82 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=6.507
r102 56 61 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.41 $Y=6.355
+ $X2=2.41 $Y2=5.835
r103 53 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.55 $Y2=6.507
r104 53 55 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=1.635 $Y=6.507
+ $X2=1.7 $Y2=6.507
r105 52 82 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=2.41 $Y2=6.507
r106 52 55 23.6156 $w=3.03e-07 $l=6.25e-07 $layer=LI1_cond $X=2.325 $Y=6.507
+ $X2=1.7 $Y2=6.507
r107 48 51 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.55 $Y=3.455
+ $X2=1.55 $Y2=5.835
r108 46 80 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=6.507
r109 46 51 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.55 $Y=6.355
+ $X2=1.55 $Y2=5.835
r110 43 79 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=0.69 $Y2=6.507
r111 43 45 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=0.775 $Y=6.507
+ $X2=1.02 $Y2=6.507
r112 42 80 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.55 $Y2=6.507
r113 42 45 16.8143 $w=3.03e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=6.507
+ $X2=1.02 $Y2=6.507
r114 38 41 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.69 $Y=4.135
+ $X2=0.69 $Y2=5.835
r115 36 79 3.51065 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=6.507
r116 36 41 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.69 $Y=6.355
+ $X2=0.69 $Y2=5.835
r117 34 99 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=3.535 $Y=6.355 $X2=3.74 $Y2=6.44
r118 34 96 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.135 $Y=6.355 $X2=0.34 $Y2=6.44
r119 34 82 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.175 $Y=6.355 $X2=2.38 $Y2=6.44
r120 34 65 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=2.855 $Y=6.355 $X2=3.06 $Y2=6.44
r121 34 55 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=1.495 $Y=6.355 $X2=1.7 $Y2=6.44
r122 34 45 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0.815 $Y=6.355 $X2=1.02 $Y2=6.44
r123 5 77 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.99
+ $Y=3.085 $X2=4.13 $Y2=5.835
r124 5 74 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.99
+ $Y=3.085 $X2=4.13 $Y2=3.455
r125 4 71 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=5.835
r126 4 68 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.13
+ $Y=3.085 $X2=3.27 $Y2=3.455
r127 3 61 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=5.835
r128 3 58 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.27
+ $Y=3.085 $X2=2.41 $Y2=3.455
r129 2 51 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=5.835
r130 2 48 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.41
+ $Y=3.085 $X2=1.55 $Y2=3.455
r131 1 41 200 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=5.835
r132 1 38 200 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=3.085 $X2=0.69 $Y2=4.135
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_8%A 3 7 10 15 16
r40 16 18 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.645
r41 16 17 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.48
+ $X2=0.585 $Y2=2.315
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=2.48 $X2=0.635 $Y2=2.48
r43 12 15 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=2.48
r44 10 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.635 $Y=3.33
+ $X2=0.635 $Y2=3.33
r45 7 18 994.766 $w=1.5e-07 $l=1.94e-06 $layer=POLY_cond $X=0.475 $Y=4.585
+ $X2=0.475 $Y2=2.645
r46 3 17 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=0.475 $Y=1.075
+ $X2=0.475 $Y2=2.315
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_8%A_27_115# 1 2 9 11 13 15 18 20 22 23 24
+ 25 26 29 31 33 34 36 40 42 44 45 47 51 54 55 57 58 60 64 66 68 69 71 75 77 79
+ 80 82 86 88 90 95 96 97 98 99 100 101 102 103 104 107 111 115 117 120
c232 77 0 1.33323e-19 $X=3.485 $Y=3.01
c233 75 0 1.33323e-19 $X=3.485 $Y=1.075
c234 66 0 1.33323e-19 $X=3.055 $Y=3.01
c235 64 0 1.33323e-19 $X=3.055 $Y=1.075
c236 55 0 1.33323e-19 $X=2.625 $Y=3.01
c237 51 0 1.33323e-19 $X=2.625 $Y=1.075
c238 42 0 1.33323e-19 $X=2.195 $Y=3.01
c239 40 0 1.33323e-19 $X=2.195 $Y=1.075
c240 31 0 1.33323e-19 $X=1.765 $Y=3.01
c241 29 0 1.33323e-19 $X=1.765 $Y=1.075
c242 20 0 1.33323e-19 $X=1.335 $Y=3.01
c243 18 0 1.33323e-19 $X=1.335 $Y=1.075
r244 121 125 36.879 $w=2.81e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=1.18 $Y2=1.935
r245 121 123 10.2918 $w=2.81e-07 $l=6e-08 $layer=POLY_cond $X=0.965 $Y=1.935
+ $X2=0.905 $Y2=1.935
r246 120 121 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.935 $X2=0.965 $Y2=1.935
r247 116 117 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.935
+ $X2=0.26 $Y2=1.935
r248 115 120 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.965 $Y2=1.935
r249 115 116 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.88 $Y=1.935
+ $X2=0.345 $Y2=1.935
r250 111 113 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=0.26 $Y=3.455
+ $X2=0.26 $Y2=5.835
r251 109 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=1.935
r252 109 111 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.26 $Y=2.02
+ $X2=0.26 $Y2=3.455
r253 105 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=1.935
r254 105 107 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.26 $Y=1.85
+ $X2=0.26 $Y2=0.825
r255 93 94 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=2.935
+ $X2=1.335 $Y2=2.935
r256 91 93 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.905 $Y=2.935
+ $X2=1.18 $Y2=2.935
r257 88 90 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.915 $Y=3.01
+ $X2=3.915 $Y2=4.585
r258 84 86 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.915 $Y=1.77
+ $X2=3.915 $Y2=1.075
r259 83 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=2.935
+ $X2=3.485 $Y2=2.935
r260 82 88 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=2.935
+ $X2=3.915 $Y2=3.01
r261 82 83 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=2.935
+ $X2=3.56 $Y2=2.935
r262 81 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.845
+ $X2=3.485 $Y2=1.845
r263 80 84 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=1.845
+ $X2=3.915 $Y2=1.77
r264 80 81 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.845
+ $X2=3.56 $Y2=1.845
r265 77 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=3.01
+ $X2=3.485 $Y2=2.935
r266 77 79 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.485 $Y=3.01
+ $X2=3.485 $Y2=4.585
r267 73 103 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.845
r268 73 75 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.485 $Y2=1.075
r269 72 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=2.935
+ $X2=3.055 $Y2=2.935
r270 71 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=2.935
+ $X2=3.485 $Y2=2.935
r271 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=2.935
+ $X2=3.13 $Y2=2.935
r272 70 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.845
+ $X2=3.055 $Y2=1.845
r273 69 103 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.485 $Y2=1.845
r274 69 70 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.845
+ $X2=3.13 $Y2=1.845
r275 66 102 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=3.01
+ $X2=3.055 $Y2=2.935
r276 66 68 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=3.055 $Y=3.01
+ $X2=3.055 $Y2=4.585
r277 62 101 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.845
r278 62 64 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.055 $Y=1.77
+ $X2=3.055 $Y2=1.075
r279 61 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=2.935
+ $X2=2.625 $Y2=2.935
r280 60 102 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=3.055 $Y2=2.935
r281 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=2.935
+ $X2=2.7 $Y2=2.935
r282 59 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.845 $X2=2.625
+ $Y2=1.845
r283 58 101 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=3.055 $Y2=1.845
r284 58 59 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.845
+ $X2=2.7 $Y2=1.845
r285 55 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=2.935
r286 55 57 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.625 $Y=3.01
+ $X2=2.625 $Y2=4.585
r287 54 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=2.86
+ $X2=2.625 $Y2=2.935
r288 53 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.92
+ $X2=2.625 $Y2=1.845
r289 53 54 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.625 $Y=1.92 $X2=2.625
+ $Y2=2.86
r290 49 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.845
r291 49 51 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.625 $Y=1.77
+ $X2=2.625 $Y2=1.075
r292 48 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=2.935
+ $X2=2.195 $Y2=2.935
r293 47 100 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.625 $Y2=2.935
r294 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=2.935
+ $X2=2.27 $Y2=2.935
r295 46 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.195 $Y2=1.845
r296 45 99 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.625 $Y2=1.845
r297 45 46 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.845
+ $X2=2.27 $Y2=1.845
r298 42 98 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=2.935
r299 42 44 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=2.195 $Y=3.01
+ $X2=2.195 $Y2=4.585
r300 38 97 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.845
r301 38 40 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.77
+ $X2=2.195 $Y2=1.075
r302 37 96 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=2.935
+ $X2=1.765 $Y2=2.935
r303 36 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=2.195 $Y2=2.935
r304 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=2.935
+ $X2=1.84 $Y2=2.935
r305 35 95 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.765 $Y2=1.845
r306 34 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=2.195 $Y2=1.845
r307 34 35 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.845
+ $X2=1.84 $Y2=1.845
r308 31 96 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=2.935
r309 31 33 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.765 $Y=3.01
+ $X2=1.765 $Y2=4.585
r310 27 95 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.845
r311 27 29 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.765 $Y=1.77
+ $X2=1.765 $Y2=1.075
r312 26 94 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=2.935
+ $X2=1.335 $Y2=2.935
r313 25 96 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.765 $Y2=2.935
r314 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=2.935
+ $X2=1.41 $Y2=2.935
r315 23 95 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.765 $Y2=1.845
r316 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.69 $Y=1.845
+ $X2=1.41 $Y2=1.845
r317 20 94 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=2.935
r318 20 22 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=1.335 $Y=3.01
+ $X2=1.335 $Y2=4.585
r319 16 24 23.2782 $w=2.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.41 $Y2=1.845
r320 16 125 26.5872 $w=2.81e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.18 $Y2=1.935
r321 16 18 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.335 $Y=1.77
+ $X2=1.335 $Y2=1.075
r322 15 93 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=2.86
+ $X2=1.18 $Y2=2.935
r323 14 125 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=1.935
r324 14 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.18 $Y=2.1
+ $X2=1.18 $Y2=2.86
r325 11 91 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=2.935
r326 11 13 506.1 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=0.905 $Y=3.01
+ $X2=0.905 $Y2=4.585
r327 7 123 17.4353 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.935
r328 7 9 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=1.075
r329 2 113 150 $w=1.7e-07 $l=2.81181e-06 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=5.835
r330 2 111 150 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=3.085 $X2=0.26 $Y2=3.455
r331 1 107 91 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.575 $X2=0.26 $Y2=0.825
.ends

.subckt PM_SKY130_OSU_SC_18T_LS__BUF_8%Y 1 2 3 4 5 6 7 8 25 26 28 30 32 35 36 37
+ 38 39 41 42 43 44 45 46 47 53 59 65 71 73 85 97 109
c167 47 0 1.33323e-19 $X=3.7 $Y=2.845
c168 46 0 1.33323e-19 $X=3.7 $Y=1.595
c169 45 0 2.66647e-19 $X=2.985 $Y=2.96
c170 43 0 2.66647e-19 $X=2.985 $Y=1.48
c171 39 0 2.66647e-19 $X=2.125 $Y=2.96
c172 37 0 2.66647e-19 $X=2.125 $Y=1.48
c173 26 0 1.33323e-19 $X=1.12 $Y=2.845
c174 25 0 1.33323e-19 $X=1.12 $Y=1.595
r175 116 118 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=3.7 $Y=3.455
+ $X2=3.7 $Y2=5.835
r176 104 106 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=2.84 $Y=3.455
+ $X2=2.84 $Y2=5.835
r177 92 94 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.98 $Y=3.455
+ $X2=1.98 $Y2=5.835
r178 80 82 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=1.12 $Y=3.455
+ $X2=1.12 $Y2=5.835
r179 71 116 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.7 $Y=2.96
+ $X2=3.7 $Y2=3.455
r180 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=2.96 $X2=3.7
+ $Y2=2.96
r181 68 109 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.7 $Y=1.48
+ $X2=3.7 $Y2=0.825
r182 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=1.48 $X2=3.7
+ $Y2=1.48
r183 65 104 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=3.455
r184 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=2.96
+ $X2=2.84 $Y2=2.96
r185 62 97 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.84 $Y=1.48
+ $X2=2.84 $Y2=0.825
r186 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=1.48
+ $X2=2.84 $Y2=1.48
r187 59 92 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=3.455
r188 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=2.96
+ $X2=1.98 $Y2=2.96
r189 56 85 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=0.825
r190 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.98 $Y=1.48
+ $X2=1.98 $Y2=1.48
r191 53 80 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=3.455
r192 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.96
+ $X2=1.12 $Y2=2.96
r193 50 73 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=0.825
r194 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.48
+ $X2=1.12 $Y2=1.48
r195 47 70 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.7 $Y=2.845
+ $X2=3.7 $Y2=2.96
r196 46 67 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=3.7 $Y=1.595
+ $X2=3.7 $Y2=1.48
r197 46 47 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=3.7 $Y=1.595
+ $X2=3.7 $Y2=2.845
r198 45 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=2.96
+ $X2=2.84 $Y2=2.96
r199 44 70 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.555 $Y=2.96
+ $X2=3.7 $Y2=2.96
r200 44 45 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.555 $Y=2.96
+ $X2=2.985 $Y2=2.96
r201 43 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=1.48
+ $X2=2.84 $Y2=1.48
r202 42 67 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=3.555 $Y=1.48
+ $X2=3.7 $Y2=1.48
r203 42 43 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=3.555 $Y=1.48
+ $X2=2.985 $Y2=1.48
r204 41 64 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=2.845
+ $X2=2.84 $Y2=2.96
r205 40 61 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=1.48
r206 40 41 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=2.84 $Y=1.595
+ $X2=2.84 $Y2=2.845
r207 39 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=2.96
+ $X2=1.98 $Y2=2.96
r208 38 64 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.84 $Y2=2.96
r209 38 39 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=2.96
+ $X2=2.125 $Y2=2.96
r210 37 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.125 $Y=1.48
+ $X2=1.98 $Y2=1.48
r211 36 61 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.84 $Y2=1.48
r212 36 37 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=2.695 $Y=1.48
+ $X2=2.125 $Y2=1.48
r213 35 58 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=2.845
+ $X2=1.98 $Y2=2.96
r214 34 55 0.0257089 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=1.48
r215 34 35 1.2036 $w=1.7e-07 $l=1.25e-06 $layer=MET1_cond $X=1.98 $Y=1.595
+ $X2=1.98 $Y2=2.845
r216 33 52 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=2.96
+ $X2=1.12 $Y2=2.96
r217 32 58 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.98 $Y2=2.96
r218 32 33 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=2.96
+ $X2=1.265 $Y2=2.96
r219 31 49 0.0389498 $w=1.7e-07 $l=1.45e-07 $layer=MET1_cond $X=1.265 $Y=1.48
+ $X2=1.12 $Y2=1.48
r220 30 55 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.98 $Y2=1.48
r221 30 31 0.548843 $w=1.7e-07 $l=5.7e-07 $layer=MET1_cond $X=1.835 $Y=1.48
+ $X2=1.265 $Y2=1.48
r222 26 52 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.96
r223 26 28 0.553657 $w=1.7e-07 $l=5.75e-07 $layer=MET1_cond $X=1.12 $Y=2.845
+ $X2=1.12 $Y2=2.27
r224 25 49 0.0308913 $w=1.7e-07 $l=1.15e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=1.48
r225 25 28 0.649946 $w=1.7e-07 $l=6.75e-07 $layer=MET1_cond $X=1.12 $Y=1.595
+ $X2=1.12 $Y2=2.27
r226 8 118 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=5.835
r227 8 116 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=3.085 $X2=3.7 $Y2=3.455
r228 7 106 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=5.835
r229 7 104 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=2.7
+ $Y=3.085 $X2=2.84 $Y2=3.455
r230 6 94 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=5.835
r231 6 92 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=1.84
+ $Y=3.085 $X2=1.98 $Y2=3.455
r232 5 82 150 $w=1.7e-07 $l=2.81913e-06 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=5.835
r233 5 80 150 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=3.085 $X2=1.12 $Y2=3.455
r234 4 109 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.575 $X2=3.7 $Y2=0.825
r235 3 97 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.575 $X2=2.84 $Y2=0.825
r236 2 85 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.575 $X2=1.98 $Y2=0.825
r237 1 73 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.575 $X2=1.12 $Y2=0.825
.ends

